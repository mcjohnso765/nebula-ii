* NGSPICE file created from team_02.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_2 abstract view
.subckt sky130_fd_sc_hd__o2111ai_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_8 abstract view
.subckt sky130_fd_sc_hd__inv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_4 abstract view
.subckt sky130_fd_sc_hd__o211a_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__bufinv_16 abstract view
.subckt sky130_fd_sc_hd__bufinv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_2 abstract view
.subckt sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_1 abstract view
.subckt sky130_fd_sc_hd__nor4b_1 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_8 abstract view
.subckt sky130_fd_sc_hd__clkinv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_16 abstract view
.subckt sky130_fd_sc_hd__inv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41ai_2 abstract view
.subckt sky130_fd_sc_hd__o41ai_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_12 abstract view
.subckt sky130_fd_sc_hd__inv_12 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_4 abstract view
.subckt sky130_fd_sc_hd__a221oi_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_4 abstract view
.subckt sky130_fd_sc_hd__or4bb_4 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_2 abstract view
.subckt sky130_fd_sc_hd__or4bb_2 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinvlp_4 abstract view
.subckt sky130_fd_sc_hd__clkinvlp_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_16 abstract view
.subckt sky130_fd_sc_hd__clkinv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_2 abstract view
.subckt sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_2 abstract view
.subckt sky130_fd_sc_hd__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_4 abstract view
.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_4 abstract view
.subckt sky130_fd_sc_hd__o41a_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_2 abstract view
.subckt sky130_fd_sc_hd__a2111oi_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_1 abstract view
.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_2 abstract view
.subckt sky130_fd_sc_hd__a41o_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_2 abstract view
.subckt sky130_fd_sc_hd__o41a_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_4 abstract view
.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_4 abstract view
.subckt sky130_fd_sc_hd__and3b_4 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_2 abstract view
.subckt sky130_fd_sc_hd__dfstp_2 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_1 abstract view
.subckt sky130_fd_sc_hd__o32ai_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311ai_4 abstract view
.subckt sky130_fd_sc_hd__o311ai_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_4 abstract view
.subckt sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_4 abstract view
.subckt sky130_fd_sc_hd__a221o_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

.subckt team_02 ACK_I ADR_O[0] ADR_O[10] ADR_O[11] ADR_O[12] ADR_O[13] ADR_O[14] ADR_O[15]
+ ADR_O[16] ADR_O[17] ADR_O[18] ADR_O[19] ADR_O[1] ADR_O[20] ADR_O[21] ADR_O[22] ADR_O[23]
+ ADR_O[24] ADR_O[25] ADR_O[26] ADR_O[27] ADR_O[28] ADR_O[29] ADR_O[2] ADR_O[30] ADR_O[31]
+ ADR_O[3] ADR_O[4] ADR_O[5] ADR_O[6] ADR_O[7] ADR_O[8] ADR_O[9] CYC_O DAT_I[0] DAT_I[10]
+ DAT_I[11] DAT_I[12] DAT_I[13] DAT_I[14] DAT_I[15] DAT_I[16] DAT_I[17] DAT_I[18]
+ DAT_I[19] DAT_I[1] DAT_I[20] DAT_I[21] DAT_I[22] DAT_I[23] DAT_I[24] DAT_I[25] DAT_I[26]
+ DAT_I[27] DAT_I[28] DAT_I[29] DAT_I[2] DAT_I[30] DAT_I[31] DAT_I[3] DAT_I[4] DAT_I[5]
+ DAT_I[6] DAT_I[7] DAT_I[8] DAT_I[9] DAT_O[0] DAT_O[10] DAT_O[11] DAT_O[12] DAT_O[13]
+ DAT_O[14] DAT_O[15] DAT_O[16] DAT_O[17] DAT_O[18] DAT_O[19] DAT_O[1] DAT_O[20] DAT_O[21]
+ DAT_O[22] DAT_O[23] DAT_O[24] DAT_O[25] DAT_O[26] DAT_O[27] DAT_O[28] DAT_O[29]
+ DAT_O[2] DAT_O[30] DAT_O[31] DAT_O[3] DAT_O[4] DAT_O[5] DAT_O[6] DAT_O[7] DAT_O[8]
+ DAT_O[9] SEL_O[0] SEL_O[1] SEL_O[2] SEL_O[3] STB_O WE_O clk en gpio_in[0] gpio_in[10]
+ gpio_in[11] gpio_in[12] gpio_in[13] gpio_in[14] gpio_in[15] gpio_in[16] gpio_in[17]
+ gpio_in[18] gpio_in[19] gpio_in[1] gpio_in[20] gpio_in[21] gpio_in[22] gpio_in[23]
+ gpio_in[24] gpio_in[25] gpio_in[26] gpio_in[27] gpio_in[28] gpio_in[29] gpio_in[2]
+ gpio_in[30] gpio_in[31] gpio_in[3] gpio_in[4] gpio_in[5] gpio_in[6] gpio_in[7] gpio_in[8]
+ gpio_in[9] gpio_out[0] gpio_out[10] gpio_out[11] gpio_out[12] gpio_out[13] gpio_out[14]
+ gpio_out[15] gpio_out[16] gpio_out[17] gpio_out[18] gpio_out[19] gpio_out[1] gpio_out[20]
+ gpio_out[21] gpio_out[22] gpio_out[23] gpio_out[24] gpio_out[25] gpio_out[26] gpio_out[27]
+ gpio_out[28] gpio_out[29] gpio_out[2] gpio_out[30] gpio_out[31] gpio_out[3] gpio_out[4]
+ gpio_out[5] gpio_out[6] gpio_out[7] gpio_out[8] gpio_out[9] nrst vccd1 vssd1
XPHY_EDGE_ROW_176_Left_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09671_ _04653_ _04706_ _04707_ net889 vssd1 vssd1 vccd1 vccd1 _00120_ sky130_fd_sc_hd__o211a_1
X_06883_ top.DUT.register\[14\]\[18\] net585 net464 top.DUT.register\[13\]\[18\] _02021_
+ vssd1 vssd1 vccd1 vccd1 _02022_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_124_2300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08622_ _03744_ vssd1 vssd1 vccd1 vccd1 _03745_ sky130_fd_sc_hd__inv_2
X_08553_ net434 _03678_ _03672_ net427 vssd1 vssd1 vccd1 vccd1 _03679_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA_fanout162_A _04906_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_194_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_194_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07298__B1 net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11094__A1 _01405_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07504_ top.DUT.register\[22\]\[14\] net649 net752 top.DUT.register\[26\]\[14\] _02642_
+ vssd1 vssd1 vccd1 vccd1 _02643_ sky130_fd_sc_hd__a221o_1
X_08484_ _03566_ _03612_ _02568_ vssd1 vssd1 vccd1 vccd1 _03613_ sky130_fd_sc_hd__o21a_1
XANTENNA__07837__A2 net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06229__A top.ramload\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_159_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_186_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07435_ top.DUT.register\[14\]\[15\] net584 net504 top.DUT.register\[27\]\[15\] vssd1
+ vssd1 vccd1 vccd1 _02574_ sky130_fd_sc_hd__a22o_1
XFILLER_0_147_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_185_Left_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1071_A net1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout427_A _03259_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_1974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07366_ top.DUT.register\[7\]\[8\] net662 net640 top.DUT.register\[8\]\[8\] vssd1
+ vssd1 vccd1 vccd1 _02505_ sky130_fd_sc_hd__a22o_1
X_09105_ _04172_ _04179_ vssd1 vssd1 vccd1 vccd1 _04180_ sky130_fd_sc_hd__nand2b_1
X_06317_ _01447_ _01469_ _01468_ _01448_ vssd1 vssd1 vccd1 vccd1 _00003_ sky130_fd_sc_hd__a2bb2o_1
X_07297_ top.DUT.register\[3\]\[12\] net551 net451 top.DUT.register\[29\]\[12\] _02435_
+ vssd1 vssd1 vccd1 vccd1 _02436_ sky130_fd_sc_hd__a221o_1
XANTENNA__09974__S net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09036_ _04108_ _04109_ _04110_ _03412_ vssd1 vssd1 vccd1 vccd1 _04111_ sky130_fd_sc_hd__or4b_1
XTAP_TAPCELL_ROW_135_2473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06248_ top.ramload\[9\] net855 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedData\[9\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_170_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout796_A net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11149__A2 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold340 top.DUT.register\[11\]\[9\] vssd1 vssd1 vccd1 vccd1 net1456 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10913__S net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_157 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06179_ _01413_ _01419_ vssd1 vssd1 vccd1 vccd1 _01421_ sky130_fd_sc_hd__nor2_1
XANTENNA__08450__Y _03580_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold351 top.DUT.register\[6\]\[4\] vssd1 vssd1 vccd1 vccd1 net1467 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13721__RESET_B net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold362 top.DUT.register\[2\]\[4\] vssd1 vssd1 vccd1 vccd1 net1478 sky130_fd_sc_hd__dlygate4sd3_1
Xhold373 top.ramaddr\[25\] vssd1 vssd1 vccd1 vccd1 net1489 sky130_fd_sc_hd__dlygate4sd3_1
Xhold384 top.DUT.register\[26\]\[6\] vssd1 vssd1 vccd1 vccd1 net1500 sky130_fd_sc_hd__dlygate4sd3_1
Xhold395 top.DUT.register\[14\]\[11\] vssd1 vssd1 vccd1 vccd1 net1511 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout963_A net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06576__A2 net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout820 _01579_ vssd1 vssd1 vccd1 vccd1 net820 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout584_X net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07773__B2 top.DUT.register\[19\]\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout831 net832 vssd1 vssd1 vccd1 vccd1 net831 sky130_fd_sc_hd__clkbuf_2
Xfanout842 _05041_ vssd1 vssd1 vccd1 vccd1 net842 sky130_fd_sc_hd__buf_2
X_09938_ net828 _04652_ vssd1 vssd1 vccd1 vccd1 _04943_ sky130_fd_sc_hd__nor2_1
Xfanout853 net854 vssd1 vssd1 vccd1 vccd1 net853 sky130_fd_sc_hd__clkbuf_2
Xfanout864 net865 vssd1 vssd1 vccd1 vccd1 net864 sky130_fd_sc_hd__clkbuf_2
Xfanout875 net876 vssd1 vssd1 vccd1 vccd1 net875 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_181_3161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout886 top.ru.state\[5\] vssd1 vssd1 vccd1 vccd1 net886 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout751_X net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout897 net899 vssd1 vssd1 vccd1 vccd1 net897 sky130_fd_sc_hd__clkbuf_4
X_09869_ top.pc\[25\] _04560_ vssd1 vssd1 vccd1 vccd1 _04880_ sky130_fd_sc_hd__nand2_1
Xhold1040 top.DUT.register\[7\]\[9\] vssd1 vssd1 vccd1 vccd1 net2156 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1051 top.lcd.cnt_20ms\[8\] vssd1 vssd1 vccd1 vccd1 net2167 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11900_ _05782_ vssd1 vssd1 vccd1 vccd1 _05783_ sky130_fd_sc_hd__inv_2
Xhold1062 top.DUT.register\[3\]\[25\] vssd1 vssd1 vccd1 vccd1 net2178 sky130_fd_sc_hd__dlygate4sd3_1
X_12880_ clknet_leaf_28_clk _00472_ net1010 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[11\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1073 top.DUT.register\[4\]\[30\] vssd1 vssd1 vccd1 vccd1 net2189 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1084 top.DUT.register\[25\]\[0\] vssd1 vssd1 vccd1 vccd1 net2200 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1095 top.DUT.register\[19\]\[11\] vssd1 vssd1 vccd1 vccd1 net2211 sky130_fd_sc_hd__dlygate4sd3_1
X_11831_ _05678_ _05689_ vssd1 vssd1 vccd1 vccd1 _05714_ sky130_fd_sc_hd__and2b_1
XANTENNA__09278__A1 net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_185_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_64_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_64_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11762_ _05572_ _05634_ vssd1 vssd1 vccd1 vccd1 _05645_ sky130_fd_sc_hd__nand2_1
XANTENNA__07828__A2 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06139__A top.lcd.nextState\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13501_ clknet_leaf_13_clk _01093_ net941 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[31\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_10713_ net1925 net217 net335 vssd1 vssd1 vccd1 vccd1 _00874_ sky130_fd_sc_hd__mux2_1
X_11693_ _05493_ _05543_ vssd1 vssd1 vccd1 vccd1 _05576_ sky130_fd_sc_hd__and2_1
XANTENNA__06500__A2 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_181_823 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13432_ clknet_leaf_127_clk _01024_ net921 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[29\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_10644_ net190 net1799 net343 vssd1 vssd1 vccd1 vccd1 _00808_ sky130_fd_sc_hd__mux2_1
XANTENNA__06426__X _01565_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_192_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13363_ clknet_leaf_123_clk _00955_ net927 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[27\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_10575_ net1432 net213 net353 vssd1 vssd1 vccd1 vccd1 _00741_ sky130_fd_sc_hd__mux2_1
XANTENNA__10095__S net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_692 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09169__B _02808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_210_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12314_ top.pad.button_control.r_counter\[5\] top.pad.button_control.r_counter\[4\]
+ _06116_ vssd1 vssd1 vccd1 vccd1 _06120_ sky130_fd_sc_hd__and3_1
XANTENNA__09737__X _04763_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07461__B1 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13294_ clknet_leaf_41_clk _00886_ net1047 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[24\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_121_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_210_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08431__A2_N net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12245_ top.lcd.cnt_20ms\[12\] top.lcd.cnt_20ms\[11\] _06074_ top.lcd.cnt_20ms\[13\]
+ vssd1 vssd1 vccd1 vccd1 _06078_ sky130_fd_sc_hd__a31o_1
XANTENNA__10823__S net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12176_ _05083_ _05968_ net1311 net847 vssd1 vssd1 vccd1 vccd1 _01284_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__06567__A2 net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_166_2934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11127_ net55 net867 vssd1 vssd1 vccd1 vccd1 _05069_ sky130_fd_sc_hd__and2_1
XFILLER_0_155_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11058_ net1187 net866 net837 top.ramstore\[9\] vssd1 vssd1 vccd1 vccd1 _01169_ sky130_fd_sc_hd__a22o_1
XFILLER_0_3_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11312__A2 _05136_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_204_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10009_ net155 net1615 net625 vssd1 vssd1 vccd1 vccd1 _00214_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_199_3433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_106_2041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09124__S _04045_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_488 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07819__A2 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_15_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07220_ _02331_ _02356_ vssd1 vssd1 vccd1 vccd1 _02359_ sky130_fd_sc_hd__or2_2
XFILLER_0_6_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07151_ top.DUT.register\[21\]\[11\] net655 net738 top.DUT.register\[12\]\[11\] _02287_
+ vssd1 vssd1 vccd1 vccd1 _02290_ sky130_fd_sc_hd__a221o_1
XFILLER_0_42_512 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09079__B top.a1.instruction\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07082_ _02198_ _02219_ vssd1 vssd1 vccd1 vccd1 _02221_ sky130_fd_sc_hd__nand2_1
XANTENNA__07452__B1 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10733__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_442 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09744__A2 _04172_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_2392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout138 net139 vssd1 vssd1 vccd1 vccd1 net138 sky130_fd_sc_hd__buf_2
Xfanout149 _04938_ vssd1 vssd1 vccd1 vccd1 net149 sky130_fd_sc_hd__buf_1
XANTENNA__06231__B net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07984_ top.DUT.register\[5\]\[31\] net653 net749 top.DUT.register\[17\]\[31\] vssd1
+ vssd1 vccd1 vccd1 _03123_ sky130_fd_sc_hd__a22o_1
X_09723_ _04172_ _02340_ _02355_ vssd1 vssd1 vccd1 vccd1 _04751_ sky130_fd_sc_hd__or3b_1
X_06935_ top.DUT.register\[1\]\[21\] net756 net712 top.DUT.register\[11\]\[21\] vssd1
+ vssd1 vccd1 vccd1 _02074_ sky130_fd_sc_hd__a22o_1
XANTENNA__11303__A2 _05123_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout377_A net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09654_ _04674_ _04689_ _04681_ vssd1 vssd1 vccd1 vccd1 _04695_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_97_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09542__B _04590_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06866_ _01983_ _02004_ vssd1 vssd1 vccd1 vccd1 _02005_ sky130_fd_sc_hd__nor2_1
X_08605_ _02266_ _03727_ vssd1 vssd1 vccd1 vccd1 _03728_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_210_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06797_ top.DUT.register\[9\]\[17\] net470 net552 top.DUT.register\[3\]\[17\] _01935_
+ vssd1 vssd1 vccd1 vccd1 _01936_ sky130_fd_sc_hd__a221o_1
X_09585_ _04627_ _04631_ vssd1 vssd1 vccd1 vccd1 _04632_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_179_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout544_A net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06730__A2 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09969__S net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08536_ _03647_ _03656_ _03662_ vssd1 vssd1 vccd1 vccd1 _03663_ sky130_fd_sc_hd__or3b_4
XPHY_EDGE_ROW_193_Left_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_46_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_166_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10908__S net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout332_X net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout711_A _01638_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08467_ _03060_ _03573_ vssd1 vssd1 vccd1 vccd1 _03596_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_137_2502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1074_X net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07418_ top.DUT.register\[23\]\[9\] net671 net746 top.DUT.register\[17\]\[9\] _02549_
+ vssd1 vssd1 vccd1 vccd1 _02557_ sky130_fd_sc_hd__a221o_1
XFILLER_0_80_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08398_ net296 _03529_ _03528_ vssd1 vssd1 vccd1 vccd1 _03530_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_52_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_93_clk_A clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07349_ top.DUT.register\[15\]\[8\] net680 net676 top.DUT.register\[31\]\[8\] vssd1
+ vssd1 vccd1 vccd1 _02488_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_150_2702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10360_ net1550 net142 net379 vssd1 vssd1 vccd1 vccd1 _00536_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout799_X net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06797__A2 net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09019_ _01875_ _02753_ _03042_ _03518_ vssd1 vssd1 vccd1 vccd1 _04094_ sky130_fd_sc_hd__or4_1
X_10291_ net1700 net156 net388 vssd1 vssd1 vccd1 vccd1 _00469_ sky130_fd_sc_hd__mux2_1
XANTENNA__10643__S net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12030_ _05899_ _05912_ vssd1 vssd1 vccd1 vccd1 _05913_ sky130_fd_sc_hd__nor2_1
Xhold170 top.ramaddr\[13\] vssd1 vssd1 vccd1 vccd1 net1286 sky130_fd_sc_hd__dlygate4sd3_1
Xhold181 top.ramstore\[3\] vssd1 vssd1 vccd1 vccd1 net1297 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06422__A top.a1.instruction\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold192 top.a1.row2\[9\] vssd1 vssd1 vccd1 vccd1 net1308 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout966_X net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout650 _01612_ vssd1 vssd1 vccd1 vccd1 net650 sky130_fd_sc_hd__clkbuf_4
XANTENNA_clkbuf_leaf_31_clk_A clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_148_2664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout661 net662 vssd1 vssd1 vccd1 vccd1 net661 sky130_fd_sc_hd__buf_4
XANTENNA__07805__X _02944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout672 _01597_ vssd1 vssd1 vccd1 vccd1 net672 sky130_fd_sc_hd__clkbuf_4
Xfanout683 _01511_ vssd1 vssd1 vccd1 vccd1 net683 sky130_fd_sc_hd__buf_2
XFILLER_0_189_208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout694 net696 vssd1 vssd1 vccd1 vccd1 net694 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_70_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12932_ clknet_leaf_36_clk _00524_ net1042 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[13\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_161_2864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12863_ clknet_leaf_15_clk _00455_ net961 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[11\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_46_clk_A clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06721__A2 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11814_ net131 _05666_ vssd1 vssd1 vccd1 vccd1 _05697_ sky130_fd_sc_hd__and2b_1
XANTENNA__11058__B2 top.ramstore\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12794_ clknet_leaf_5_clk _00386_ net936 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[9\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_194_3352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07540__X _02679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_194_3363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_32_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11745_ _05626_ _05627_ vssd1 vssd1 vccd1 vccd1 _05628_ sky130_fd_sc_hd__or2_1
XANTENNA__10818__S net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_480 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11676_ _05527_ _05528_ _05549_ vssd1 vssd1 vccd1 vccd1 _05559_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_12_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13415_ clknet_leaf_6_clk _01007_ net938 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[28\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_180_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10627_ net142 net1675 net348 vssd1 vssd1 vccd1 vccd1 _00792_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_104_clk_A clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_181_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07434__B1 net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13346_ clknet_leaf_8_clk _00938_ net947 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[26\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_10558_ net1377 net158 net355 vssd1 vssd1 vccd1 vccd1 _00725_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06788__A2 net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10553__S net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13277_ clknet_leaf_119_clk _00869_ net954 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[24\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_10489_ net2304 net165 net364 vssd1 vssd1 vccd1 vccd1 _00659_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12228_ _01383_ _06054_ _06067_ net978 vssd1 vssd1 vccd1 vccd1 _01317_ sky130_fd_sc_hd__o211a_1
XANTENNA__09726__A2 net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_119_clk_A clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12159_ _06035_ _06041_ vssd1 vssd1 vccd1 vccd1 _06042_ sky130_fd_sc_hd__nand2_1
XFILLER_0_208_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_68 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06960__A2 net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06720_ top.DUT.register\[10\]\[25\] net770 net742 top.DUT.register\[2\]\[25\] vssd1
+ vssd1 vccd1 vccd1 _01859_ sky130_fd_sc_hd__a22o_1
XFILLER_0_189_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09930__X _04936_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06651_ _01789_ vssd1 vssd1 vccd1 vccd1 _01790_ sky130_fd_sc_hd__inv_2
XANTENNA__06712__A2 net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06582_ _01711_ _01720_ vssd1 vssd1 vccd1 vccd1 _01721_ sky130_fd_sc_hd__nor2_2
X_09370_ _04428_ _04429_ vssd1 vssd1 vccd1 vccd1 _04430_ sky130_fd_sc_hd__or2_1
XFILLER_0_74_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07450__X _02589_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08321_ _02852_ _03050_ vssd1 vssd1 vccd1 vccd1 _03456_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_24_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10728__S net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08953__A2_N _04050_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08252_ net298 _03370_ _03367_ vssd1 vssd1 vccd1 vccd1 _03389_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07673__B1 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_2232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07203_ _01509_ net793 vssd1 vssd1 vccd1 vccd1 _02342_ sky130_fd_sc_hd__nor2_1
XFILLER_0_15_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08183_ net302 _03320_ vssd1 vssd1 vccd1 vccd1 _03321_ sky130_fd_sc_hd__or2_1
XFILLER_0_172_664 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06226__B net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07134_ top.DUT.register\[12\]\[11\] net531 net515 top.DUT.register\[7\]\[11\] _02272_
+ vssd1 vssd1 vccd1 vccd1 _02273_ sky130_fd_sc_hd__a221o_1
XFILLER_0_42_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07425__B1 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_591 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_2421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08968__A2_N net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10971__B net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_2432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07065_ top.DUT.register\[24\]\[22\] net644 net739 top.DUT.register\[12\]\[22\] _02203_
+ vssd1 vssd1 vccd1 vccd1 _02204_ sky130_fd_sc_hd__a221o_1
XANTENNA__10463__S net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout494_A net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout661_A net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07967_ top.DUT.register\[16\]\[31\] net545 net513 top.DUT.register\[24\]\[31\] _03105_
+ vssd1 vssd1 vccd1 vccd1 _03106_ sky130_fd_sc_hd__a221o_1
XFILLER_0_199_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout759_A _01617_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09706_ net2284 net256 net633 vssd1 vssd1 vccd1 vccd1 _00125_ sky130_fd_sc_hd__mux2_1
X_06918_ top.DUT.register\[10\]\[21\] net521 net505 top.DUT.register\[27\]\[21\] vssd1
+ vssd1 vccd1 vccd1 _02057_ sky130_fd_sc_hd__a22o_1
XANTENNA__08169__A _01983_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07898_ top.DUT.register\[22\]\[1\] net576 net556 top.DUT.register\[28\]\[1\] vssd1
+ vssd1 vccd1 vccd1 _03037_ sky130_fd_sc_hd__a22o_1
X_09637_ _04677_ _04678_ vssd1 vssd1 vccd1 vccd1 _04679_ sky130_fd_sc_hd__nor2_1
XANTENNA__11307__B _05130_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06849_ top.DUT.register\[20\]\[19\] net665 net650 top.DUT.register\[22\]\[19\] _01987_
+ vssd1 vssd1 vccd1 vccd1 _01988_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout547_X net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout926_A net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06703__A2 net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_143_2594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09568_ _04614_ _04615_ vssd1 vssd1 vccd1 vccd1 _04616_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_167_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08519_ _02475_ net431 net499 _02474_ vssd1 vssd1 vccd1 vccd1 _03646_ sky130_fd_sc_hd__a22o_1
XANTENNA__10638__S net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_194_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout714_X net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09499_ top.pc\[25\] _04543_ vssd1 vssd1 vccd1 vccd1 _04551_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_176_3082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08616__B net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_176_3093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11323__A top.a1.dataIn\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11530_ _05370_ _05371_ _05396_ _05398_ _05366_ vssd1 vssd1 vccd1 vccd1 _05413_ sky130_fd_sc_hd__a221o_1
XFILLER_0_65_467 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07927__A_N _02329_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08463__A1_N net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_163_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_128 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_137_Right_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11461_ _05287_ net278 _05306_ vssd1 vssd1 vccd1 vccd1 _05344_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_80_448 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13200_ clknet_leaf_29_clk _00792_ net1017 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[21\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07416__B1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10412_ net1477 net189 net369 vssd1 vssd1 vccd1 vccd1 _00584_ sky130_fd_sc_hd__mux2_1
X_11392_ _05273_ _05274_ _05243_ vssd1 vssd1 vccd1 vccd1 _05275_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_59_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13131_ clknet_leaf_50_clk _00723_ net1059 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[19\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10373__S net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10343_ net1745 net196 net379 vssd1 vssd1 vccd1 vccd1 _00519_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09708__A2 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07248__A _02329_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13062_ clknet_leaf_33_clk _00654_ net1044 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[17\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_10274_ net2024 net220 net385 vssd1 vssd1 vccd1 vccd1 _00452_ sky130_fd_sc_hd__mux2_1
XANTENNA__06152__A top.a1.dataIn\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12013_ _05865_ net126 _05866_ vssd1 vssd1 vccd1 vccd1 _05896_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08931__A3 _03187_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06942__A2 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout480 _04964_ vssd1 vssd1 vccd1 vccd1 net480 sky130_fd_sc_hd__buf_6
XFILLER_0_136_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout491 _04721_ vssd1 vssd1 vccd1 vccd1 net491 sky130_fd_sc_hd__buf_2
XANTENNA__08079__A _02242_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12915_ clknet_leaf_120_clk _00507_ net932 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[13\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_17_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12846_ clknet_leaf_43_clk _00438_ net1064 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[10\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09910__B net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_185_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07711__A net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_173_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12777_ clknet_leaf_21_clk _00369_ net1033 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[8\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_145_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10548__S net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_620 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07430__B _02567_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11728_ _05606_ _05607_ vssd1 vssd1 vccd1 vccd1 _05611_ sky130_fd_sc_hd__or2_1
XANTENNA__07655__B1 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_104_Right_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11659_ _05529_ _05535_ _05537_ _05541_ _05494_ vssd1 vssd1 vccd1 vccd1 _05542_ sky130_fd_sc_hd__o2111ai_2
XTAP_TAPCELL_ROW_211_3606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_211_3617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_211_3628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07958__A1 _01722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold906 top.DUT.register\[3\]\[20\] vssd1 vssd1 vccd1 vccd1 net2022 sky130_fd_sc_hd__dlygate4sd3_1
Xhold917 top.DUT.register\[21\]\[16\] vssd1 vssd1 vccd1 vccd1 net2033 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10283__S net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13329_ clknet_leaf_115_clk _00921_ net966 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[26\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_114_2151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold928 top.DUT.register\[24\]\[1\] vssd1 vssd1 vccd1 vccd1 net2044 sky130_fd_sc_hd__dlygate4sd3_1
Xhold939 top.DUT.register\[25\]\[12\] vssd1 vssd1 vccd1 vccd1 net2055 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_712 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_2162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_3_1_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_3_1_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_20_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08870_ _01745_ _01785_ _03095_ vssd1 vssd1 vccd1 vccd1 _03981_ sky130_fd_sc_hd__nor3_1
XANTENNA__13431__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07186__A2 net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_209_3579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_208_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07821_ top.DUT.register\[25\]\[0\] net778 net702 top.DUT.register\[3\]\[0\] vssd1
+ vssd1 vccd1 vccd1 _02960_ sky130_fd_sc_hd__a22o_1
XANTENNA__10190__A1 _04712_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06933__A2 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_208_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07752_ top.DUT.register\[7\]\[3\] net517 _02890_ vssd1 vssd1 vccd1 vccd1 _02891_
+ sky130_fd_sc_hd__a21o_1
X_06703_ top.DUT.register\[9\]\[25\] net470 net559 top.DUT.register\[2\]\[25\] _01841_
+ vssd1 vssd1 vccd1 vccd1 _01842_ sky130_fd_sc_hd__a221o_1
XFILLER_0_79_537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11127__B net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07683_ top.DUT.register\[30\]\[4\] net760 net748 top.DUT.register\[17\]\[4\] vssd1
+ vssd1 vccd1 vccd1 _02822_ sky130_fd_sc_hd__a22o_1
XANTENNA__09883__A1 net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_177_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09422_ top.pc\[20\] _04461_ vssd1 vssd1 vccd1 vccd1 _04479_ sky130_fd_sc_hd__nor2_1
X_06634_ top.DUT.register\[14\]\[27\] net733 _01767_ _01769_ _01772_ vssd1 vssd1 vccd1
+ vccd1 _01773_ sky130_fd_sc_hd__a2111o_1
XANTENNA__12219__B1 net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07894__B1 net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08717__A _03342_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09353_ top.pc\[16\] _04403_ vssd1 vssd1 vccd1 vccd1 _04414_ sky130_fd_sc_hd__nor2_1
XANTENNA__10458__S net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06565_ top.DUT.register\[6\]\[28\] net569 net453 top.DUT.register\[29\]\[28\] _01703_
+ vssd1 vssd1 vccd1 vccd1 _01704_ sky130_fd_sc_hd__a221o_1
XFILLER_0_19_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout242_A _04745_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08304_ net297 _03438_ vssd1 vssd1 vccd1 vccd1 _03439_ sky130_fd_sc_hd__nand2_1
XFILLER_0_191_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07646__B1 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06496_ net788 _01596_ _01618_ vssd1 vssd1 vccd1 vccd1 _01635_ sky130_fd_sc_hd__and3_4
X_09284_ _04347_ _04348_ vssd1 vssd1 vccd1 vccd1 _04349_ sky130_fd_sc_hd__and2b_1
XFILLER_0_90_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06237__A top.ramload\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07110__A2 net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08235_ net295 _03371_ _03370_ vssd1 vssd1 vccd1 vccd1 _03372_ sky130_fd_sc_hd__o21a_1
XFILLER_0_144_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_160_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout507_A _01565_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08166_ _02198_ net329 vssd1 vssd1 vccd1 vccd1 _03304_ sky130_fd_sc_hd__nand2_1
XFILLER_0_160_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07117_ top.DUT.register\[21\]\[16\] net656 net723 top.DUT.register\[29\]\[16\] _02254_
+ vssd1 vssd1 vccd1 vccd1 _02256_ sky130_fd_sc_hd__a221o_1
X_08097_ _03232_ _03235_ net291 vssd1 vssd1 vccd1 vccd1 _03236_ sky130_fd_sc_hd__mux2_1
XANTENNA__10046__X _04954_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09982__S net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07048_ top.DUT.register\[24\]\[22\] net512 net440 top.DUT.register\[5\]\[22\] _02186_
+ vssd1 vssd1 vccd1 vccd1 _02187_ sky130_fd_sc_hd__a221o_1
XANTENNA__09835__X _04850_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload90 clknet_leaf_58_clk vssd1 vssd1 vccd1 vccd1 clkload90/Y sky130_fd_sc_hd__inv_8
XFILLER_0_30_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout876_A net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout497_X net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10921__S net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08374__A1 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07177__A2 net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09283__A top.pc\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_2623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08999_ _03505_ _03543_ _04073_ vssd1 vssd1 vccd1 vccd1 _04074_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout664_X net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06924__A2 net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_178_3111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10961_ top.a1.dataInTemp\[0\] net785 vssd1 vssd1 vccd1 vccd1 _05004_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_206_Right_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_178_3122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09874__A1 _03929_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12700_ clknet_leaf_130_clk _00292_ net909 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[6\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_13680_ clknet_leaf_91_clk _01256_ net996 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07885__B1 net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10892_ top.DUT.register\[30\]\[4\] net255 net481 vssd1 vssd1 vccd1 vccd1 _01053_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12631_ clknet_leaf_129_clk _00223_ net911 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[4\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_195_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_167_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10368__S net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_191_3311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10595__C net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_183_759 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12562_ clknet_leaf_31_clk _00154_ net1021 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[2\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_404 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13304__CLK clknet_leaf_128_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07101__A2 net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11513_ _05391_ _05393_ _05395_ _05383_ vssd1 vssd1 vccd1 vccd1 _05396_ sky130_fd_sc_hd__o31a_2
XTAP_TAPCELL_ROW_22_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12493_ clknet_leaf_87_clk _00085_ net1006 vssd1 vssd1 vccd1 vccd1 top.pc\[5\] sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_156_2785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11444_ top.a1.dataIn\[17\] _05287_ net278 vssd1 vssd1 vccd1 vccd1 _05327_ sky130_fd_sc_hd__and3_1
XFILLER_0_33_150 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11375_ top.a1.dataIn\[21\] top.a1.dataIn\[19\] _05220_ vssd1 vssd1 vccd1 vccd1 _05258_
+ sky130_fd_sc_hd__or3_1
XFILLER_0_21_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_189_3284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13114_ clknet_leaf_4_clk _00706_ net939 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[19\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_10326_ net151 net2303 net383 vssd1 vssd1 vccd1 vccd1 _00503_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13045_ clknet_leaf_34_clk _00637_ net1043 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[17\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_4_2__f_clk clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_2__leaf_clk sky130_fd_sc_hd__clkbuf_16
XANTENNA__08970__A1_N _01829_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10257_ net161 net1300 net391 vssd1 vssd1 vccd1 vccd1 _00436_ sky130_fd_sc_hd__mux2_1
XANTENNA__10831__S net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10188_ net689 _04967_ vssd1 vssd1 vccd1 vccd1 _04968_ sky130_fd_sc_hd__or2_1
XANTENNA__06376__B1 net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06915__A2 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08117__A1 net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_205_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_85_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_159_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07876__B1 net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07340__A2 net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12829_ clknet_leaf_13_clk _00421_ net953 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[10\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10278__S net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06350_ top.pad.button_control.r_counter\[14\] top.pad.button_control.r_counter\[13\]
+ top.pad.button_control.r_counter\[12\] top.pad.button_control.r_counter\[11\] vssd1
+ vssd1 vccd1 vccd1 _01490_ sky130_fd_sc_hd__or4_1
XFILLER_0_173_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06281_ top.lcd.cnt_500hz\[7\] top.lcd.cnt_500hz\[6\] top.lcd.cnt_500hz\[11\] top.lcd.cnt_500hz\[4\]
+ vssd1 vssd1 vccd1 vccd1 _01444_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_71_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08020_ _01589_ _03157_ _03152_ vssd1 vssd1 vccd1 vccd1 _03159_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_112_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold703 top.DUT.register\[27\]\[12\] vssd1 vssd1 vccd1 vccd1 net1819 sky130_fd_sc_hd__dlygate4sd3_1
Xhold714 top.DUT.register\[29\]\[11\] vssd1 vssd1 vccd1 vccd1 net1830 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold725 top.DUT.register\[18\]\[3\] vssd1 vssd1 vccd1 vccd1 net1841 sky130_fd_sc_hd__dlygate4sd3_1
Xhold736 top.a1.row2\[27\] vssd1 vssd1 vccd1 vccd1 net1852 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_96_1887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold747 top.DUT.register\[21\]\[17\] vssd1 vssd1 vccd1 vccd1 net1863 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06377__A_N top.a1.instruction\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold758 top.ramaddr\[9\] vssd1 vssd1 vccd1 vccd1 net1874 sky130_fd_sc_hd__dlygate4sd3_1
X_09971_ net1524 net166 net630 vssd1 vssd1 vccd1 vccd1 _00179_ sky130_fd_sc_hd__mux2_1
Xhold769 top.DUT.register\[25\]\[20\] vssd1 vssd1 vccd1 vccd1 net1885 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07800__B1 net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08922_ net1335 net831 net800 _04030_ vssd1 vssd1 vccd1 vccd1 _00048_ sky130_fd_sc_hd__a22o_1
XANTENNA__10741__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07159__A2 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08853_ _01790_ _03094_ vssd1 vssd1 vccd1 vccd1 _03965_ sky130_fd_sc_hd__and2_1
XANTENNA__08211__S net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout192_A _04850_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07804_ _02936_ _02938_ _02940_ _02942_ vssd1 vssd1 vccd1 vccd1 _02943_ sky130_fd_sc_hd__or4_4
X_08784_ _03856_ _03898_ net289 vssd1 vssd1 vccd1 vccd1 _03899_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_127_2353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07735_ top.DUT.register\[5\]\[3\] net653 net713 top.DUT.register\[11\]\[3\] _02873_
+ vssd1 vssd1 vccd1 vccd1 _02874_ sky130_fd_sc_hd__a221o_1
XANTENNA__08659__A2 _03185_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout457_A net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_211_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_2542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07867__B1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07666_ top.a1.instruction\[24\] _01507_ net793 top.a1.instruction\[16\] _02804_
+ vssd1 vssd1 vccd1 vccd1 _02805_ sky130_fd_sc_hd__a221o_2
XTAP_TAPCELL_ROW_140_2553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07331__A2 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09405_ _04461_ _04462_ vssd1 vssd1 vccd1 vccd1 _04463_ sky130_fd_sc_hd__or2_1
X_06617_ top.DUT.register\[10\]\[27\] net521 net505 top.DUT.register\[27\]\[27\] vssd1
+ vssd1 vccd1 vccd1 _01756_ sky130_fd_sc_hd__a22o_1
XFILLER_0_192_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09608__A1 net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07597_ top.DUT.register\[22\]\[6\] net647 net718 top.DUT.register\[19\]\[6\] vssd1
+ vssd1 vccd1 vccd1 _02736_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout624_A net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07619__B1 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09336_ _04396_ _04397_ vssd1 vssd1 vccd1 vccd1 _04398_ sky130_fd_sc_hd__or2_1
X_06548_ top.DUT.register\[4\]\[29\] net669 net716 top.DUT.register\[27\]\[29\] vssd1
+ vssd1 vccd1 vccd1 _01687_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_173_3041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10916__S net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09267_ _04331_ _04332_ vssd1 vssd1 vccd1 vccd1 _04333_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_145_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08831__A2 net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06479_ top.a1.instruction\[22\] top.a1.instruction\[23\] vssd1 vssd1 vccd1 vccd1
+ _01618_ sky130_fd_sc_hd__nor2_2
X_08218_ _03220_ _03242_ net291 vssd1 vssd1 vccd1 vccd1 _03355_ sky130_fd_sc_hd__mux2_1
XFILLER_0_172_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_576 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09198_ top.pc\[6\] top.pc\[7\] _04236_ vssd1 vssd1 vccd1 vccd1 _04268_ sky130_fd_sc_hd__and3_1
XANTENNA__11179__B1 net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout993_A net1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08149_ _03285_ _03286_ vssd1 vssd1 vccd1 vccd1 _03287_ sky130_fd_sc_hd__nand2_1
XFILLER_0_160_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07398__A2 net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12628__RESET_B net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11160_ _01409_ _05088_ vssd1 vssd1 vccd1 vccd1 _05089_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout781_X net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_698 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10111_ net1451 net141 net613 vssd1 vssd1 vccd1 vccd1 _00312_ sky130_fd_sc_hd__mux2_1
XANTENNA__10651__S net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11091_ net67 net864 vssd1 vssd1 vccd1 vccd1 _05051_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_8_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10042_ net1373 net158 net621 vssd1 vssd1 vccd1 vccd1 _00245_ sky130_fd_sc_hd__mux2_1
XANTENNA__09544__B1 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold30 top.a1.row1\[12\] vssd1 vssd1 vccd1 vccd1 net1146 sky130_fd_sc_hd__dlygate4sd3_1
Xhold41 net123 vssd1 vssd1 vccd1 vccd1 net1157 sky130_fd_sc_hd__dlygate4sd3_1
Xhold52 top.a1.row1\[113\] vssd1 vssd1 vccd1 vccd1 net1168 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold63 net112 vssd1 vssd1 vccd1 vccd1 net1179 sky130_fd_sc_hd__dlygate4sd3_1
Xhold74 top.lcd.cnt_20ms\[5\] vssd1 vssd1 vccd1 vccd1 net1190 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_188_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold85 top.a1.row1\[19\] vssd1 vssd1 vccd1 vccd1 net1201 sky130_fd_sc_hd__dlygate4sd3_1
X_13801_ clknet_leaf_71_clk _01370_ net1086 vssd1 vssd1 vccd1 vccd1 top.pad.keyCode\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07570__A2 net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07813__X _02952_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold96 top.a1.row1\[18\] vssd1 vssd1 vccd1 vccd1 net1212 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_input18_A DAT_I[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11993_ _05803_ _05875_ vssd1 vssd1 vccd1 vccd1 _05876_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09847__A1 net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08628__Y _03750_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_10__f_clk clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_10__leaf_clk
+ sky130_fd_sc_hd__clkbuf_16
X_13732_ clknet_leaf_96_clk _01303_ vssd1 vssd1 vccd1 vccd1 top.a1.dataInTemp\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_67_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09460__B _04514_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10944_ net1446 net174 net591 vssd1 vssd1 vccd1 vccd1 _01105_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_67_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07322__A2 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10098__S net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_158_2814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13663_ clknet_leaf_92_clk _01239_ net995 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[113\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06530__B1 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10875_ net184 net1783 net597 vssd1 vssd1 vccd1 vccd1 _01036_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12614_ clknet_leaf_41_clk _00206_ net1046 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[3\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13594_ clknet_leaf_63_clk net1153 net1090 vssd1 vssd1 vccd1 vccd1 net86 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_171_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12545_ clknet_leaf_16_clk _00137_ net961 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[1\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_136_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_170_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10826__S net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_612 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12476_ clknet_leaf_63_clk _00071_ net1090 vssd1 vssd1 vccd1 vccd1 top.ramstore\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08092__A _02678_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06605__A _01721_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_5 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11427_ _05266_ _05273_ _05274_ _05285_ vssd1 vssd1 vccd1 vccd1 _05310_ sky130_fd_sc_hd__or4bb_1
XANTENNA__07389__A2 net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_2110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09916__A _04151_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11358_ top.a1.dataIn\[25\] _05232_ _05231_ _05207_ vssd1 vssd1 vccd1 vccd1 _05241_
+ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__06597__B1 net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10561__S net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10309_ net208 net1488 net382 vssd1 vssd1 vccd1 vccd1 _00486_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_169_2976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11289_ net879 _05120_ _05128_ top.lcd.nextState\[3\] vssd1 vssd1 vccd1 vccd1 _05179_
+ sky130_fd_sc_hd__and4b_1
XANTENNA__08338__A1 net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_169_2987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13028_ clknet_leaf_36_clk _00620_ net1049 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[16\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_206_3538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1050 net1052 vssd1 vssd1 vccd1 vccd1 net1050 sky130_fd_sc_hd__clkbuf_2
Xfanout1061 net1070 vssd1 vssd1 vccd1 vccd1 net1061 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_177_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1072 net1073 vssd1 vssd1 vccd1 vccd1 net1072 sky130_fd_sc_hd__clkbuf_4
Xfanout1083 net1087 vssd1 vssd1 vccd1 vccd1 net1083 sky130_fd_sc_hd__clkbuf_4
Xfanout1094 net1095 vssd1 vssd1 vccd1 vccd1 net1094 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_179_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_109_2083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07520_ _02390_ _02478_ _02614_ _02658_ vssd1 vssd1 vccd1 vccd1 _02659_ sky130_fd_sc_hd__or4b_1
XANTENNA__07849__B1 net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_687 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08510__A1 net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_2272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08510__B2 _03334_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07451_ _02580_ _02589_ vssd1 vssd1 vccd1 vccd1 _02590_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_122_2283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06521__B1 net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06402_ top.a1.instruction\[16\] net685 _01522_ _01531_ vssd1 vssd1 vccd1 vccd1 _01541_
+ sky130_fd_sc_hd__and4_4
XFILLER_0_91_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07382_ _02513_ _02520_ vssd1 vssd1 vccd1 vccd1 _02521_ sky130_fd_sc_hd__nor2_2
XFILLER_0_123_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09121_ _02904_ _02934_ _02943_ _04195_ vssd1 vssd1 vccd1 vccd1 _04196_ sky130_fd_sc_hd__o31a_1
XFILLER_0_134_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06333_ net893 _01479_ vssd1 vssd1 vccd1 vccd1 _01480_ sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_123_clk clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_123_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__10736__S net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_1916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06264_ top.ramload\[25\] net853 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedData\[25\]
+ sky130_fd_sc_hd__and2_1
X_09052_ _03645_ _03673_ _03696_ _03711_ vssd1 vssd1 vccd1 vccd1 _04127_ sky130_fd_sc_hd__or4_1
XFILLER_0_72_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08003_ net807 _03141_ net437 vssd1 vssd1 vccd1 vccd1 _03142_ sky130_fd_sc_hd__o21a_2
XFILLER_0_130_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold500 top.DUT.register\[2\]\[6\] vssd1 vssd1 vccd1 vccd1 net1616 sky130_fd_sc_hd__dlygate4sd3_1
X_06195_ top.ru.state\[6\] net887 top.Wen vssd1 vssd1 vccd1 vccd1 _00012_ sky130_fd_sc_hd__a21o_1
XFILLER_0_142_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold511 top.DUT.register\[18\]\[22\] vssd1 vssd1 vccd1 vccd1 net1627 sky130_fd_sc_hd__dlygate4sd3_1
Xhold522 top.DUT.register\[21\]\[21\] vssd1 vssd1 vccd1 vccd1 net1638 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout205_A net206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_440 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06234__B net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold533 top.DUT.register\[11\]\[5\] vssd1 vssd1 vccd1 vccd1 net1649 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_164 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold544 top.DUT.register\[16\]\[22\] vssd1 vssd1 vccd1 vccd1 net1660 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06588__B1 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold555 top.DUT.register\[22\]\[24\] vssd1 vssd1 vccd1 vccd1 net1671 sky130_fd_sc_hd__dlygate4sd3_1
Xhold566 top.DUT.register\[27\]\[1\] vssd1 vssd1 vccd1 vccd1 net1682 sky130_fd_sc_hd__dlygate4sd3_1
Xhold577 top.DUT.register\[27\]\[14\] vssd1 vssd1 vccd1 vccd1 net1693 sky130_fd_sc_hd__dlygate4sd3_1
Xhold588 top.DUT.register\[22\]\[10\] vssd1 vssd1 vccd1 vccd1 net1704 sky130_fd_sc_hd__dlygate4sd3_1
X_09954_ net2254 net231 net627 vssd1 vssd1 vccd1 vccd1 _00162_ sky130_fd_sc_hd__mux2_1
XANTENNA__10471__S net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold599 top.DUT.register\[23\]\[28\] vssd1 vssd1 vccd1 vccd1 net1715 sky130_fd_sc_hd__dlygate4sd3_1
X_08905_ _01659_ _04013_ vssd1 vssd1 vccd1 vccd1 _04014_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_5_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09885_ net489 _04886_ _04894_ vssd1 vssd1 vccd1 vccd1 _04895_ sky130_fd_sc_hd__and3_2
XANTENNA_fanout574_A _01519_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08836_ net424 _03948_ _03946_ vssd1 vssd1 vccd1 vccd1 _03949_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07552__A2 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08767_ net284 _03739_ vssd1 vssd1 vccd1 vccd1 _03883_ sky130_fd_sc_hd__nor2_1
XANTENNA__06760__B1 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout362_X net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout741_A _01624_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout839_A net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07718_ top.a1.instruction\[24\] _01577_ _02856_ vssd1 vssd1 vccd1 vccd1 _02857_
+ sky130_fd_sc_hd__o21a_4
XFILLER_0_200_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_196_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08177__A _01722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08698_ net317 _03441_ _03442_ _03536_ vssd1 vssd1 vccd1 vccd1 _03817_ sky130_fd_sc_hd__o31a_1
XFILLER_0_184_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07081__A _02198_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11100__A3 net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_165_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_24_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07649_ top.DUT.register\[11\]\[5\] net710 net702 top.DUT.register\[3\]\[5\] _02780_
+ vssd1 vssd1 vccd1 vccd1 _02788_ sky130_fd_sc_hd__a221o_1
XANTENNA__06512__B1 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_177_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout627_X net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10660_ net141 net1784 net344 vssd1 vssd1 vccd1 vccd1 _00824_ sky130_fd_sc_hd__mux2_1
XANTENNA__08464__X _03594_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08905__A _01659_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_62_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09319_ top.pc\[14\] _04370_ vssd1 vssd1 vccd1 vccd1 _04382_ sky130_fd_sc_hd__or2_1
XFILLER_0_91_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10646__S net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10591_ net1522 net157 net352 vssd1 vssd1 vccd1 vccd1 _00757_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_114_clk clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_114_clk
+ sky130_fd_sc_hd__clkbuf_8
X_12330_ top.pad.button_control.r_counter\[10\] top.pad.button_control.r_counter\[9\]
+ _06126_ top.pad.button_control.r_counter\[11\] vssd1 vssd1 vccd1 vccd1 _06130_ sky130_fd_sc_hd__a31o_1
XANTENNA__12809__RESET_B net1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_153_2744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12261_ _01434_ net686 _06087_ vssd1 vssd1 vccd1 vccd1 _01336_ sky130_fd_sc_hd__and3_1
XFILLER_0_121_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11212_ _05112_ net1219 net471 vssd1 vssd1 vccd1 vccd1 _01256_ sky130_fd_sc_hd__mux2_1
XANTENNA__08568__B2 net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_186_3232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_186_3243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12192_ net1120 top.a1.dataIn\[0\] _06049_ vssd1 vssd1 vccd1 vccd1 _01299_ sky130_fd_sc_hd__mux2_1
XANTENNA__06579__B1 net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput42 net42 vssd1 vssd1 vccd1 vccd1 ADR_O[11] sky130_fd_sc_hd__buf_2
XFILLER_0_120_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10381__S net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput53 net53 vssd1 vssd1 vccd1 vccd1 ADR_O[21] sky130_fd_sc_hd__buf_2
X_11143_ net64 net868 vssd1 vssd1 vccd1 vccd1 _05077_ sky130_fd_sc_hd__and2_1
XANTENNA__09455__B _04499_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput64 net64 vssd1 vssd1 vccd1 vccd1 ADR_O[31] sky130_fd_sc_hd__buf_2
XFILLER_0_101_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput75 net75 vssd1 vssd1 vccd1 vccd1 DAT_O[11] sky130_fd_sc_hd__buf_2
XFILLER_0_101_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput86 net86 vssd1 vssd1 vccd1 vccd1 DAT_O[21] sky130_fd_sc_hd__clkbuf_4
XANTENNA__07791__A2 net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput97 net97 vssd1 vssd1 vccd1 vccd1 DAT_O[31] sky130_fd_sc_hd__clkbuf_4
X_11074_ net90 net871 net835 net1162 vssd1 vssd1 vccd1 vccd1 _01185_ sky130_fd_sc_hd__a22o_1
XANTENNA__06160__A top.a1.dataIn\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_208_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10025_ net1858 net222 net619 vssd1 vssd1 vccd1 vccd1 _00228_ sky130_fd_sc_hd__mux2_1
XFILLER_0_208_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output124_A net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06751__B1 net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_201_3457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_201_3468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11976_ _05847_ _05849_ _05755_ _05835_ vssd1 vssd1 vccd1 vccd1 _05859_ sky130_fd_sc_hd__a211oi_1
XPHY_EDGE_ROW_88_Left_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13715_ clknet_leaf_96_clk _01286_ net984 vssd1 vssd1 vccd1 vccd1 top.a1.row2\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_10927_ net246 top.DUT.register\[31\]\[7\] _04972_ vssd1 vssd1 vccd1 vccd1 _01088_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_197_3394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13646_ clknet_leaf_94_clk _00007_ net983 vssd1 vssd1 vccd1 vccd1 top.ru.state\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_10858_ net266 net1767 net594 vssd1 vssd1 vccd1 vccd1 _01019_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_156_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13577_ clknet_leaf_46_clk net1223 net1066 vssd1 vssd1 vccd1 vccd1 net99 sky130_fd_sc_hd__dfrtp_1
XANTENNA__10556__S net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_105_clk clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_105_clk
+ sky130_fd_sc_hd__clkbuf_8
X_10789_ net1424 net152 net485 vssd1 vssd1 vccd1 vccd1 _00950_ sky130_fd_sc_hd__mux2_1
X_12528_ clknet_leaf_85_clk _00120_ net1006 vssd1 vssd1 vccd1 vccd1 top.pc\[1\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_54_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12459_ clknet_leaf_46_clk _00054_ net1066 vssd1 vssd1 vccd1 vccd1 top.ramstore\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_169_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07718__X _02857_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_1835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_1846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10291__S net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout309 net310 vssd1 vssd1 vccd1 vccd1 net309 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__07782__A2 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06951_ _02069_ _02089_ vssd1 vssd1 vccd1 vccd1 _02090_ sky130_fd_sc_hd__and2_2
XANTENNA__06990__B1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06501__C _01607_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09670_ net899 net139 top.pc\[1\] vssd1 vssd1 vccd1 vccd1 _04707_ sky130_fd_sc_hd__a21o_1
XFILLER_0_118_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06882_ top.DUT.register\[28\]\[18\] net556 net528 top.DUT.register\[26\]\[18\] vssd1
+ vssd1 vccd1 vccd1 _02021_ sky130_fd_sc_hd__a22o_1
XANTENNA__07534__A2 net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_2301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09381__A _01930_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_2312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08731__B2 _03848_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08621_ net423 _03730_ _03743_ vssd1 vssd1 vccd1 vccd1 _03744_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_179_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06742__B1 net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08552_ net296 _03676_ _03677_ net319 vssd1 vssd1 vccd1 vccd1 _03678_ sky130_fd_sc_hd__a211o_1
XANTENNA__07613__B _02749_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08629__A2_N _03185_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_350 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07503_ top.DUT.register\[12\]\[14\] net739 net736 top.DUT.register\[16\]\[14\] vssd1
+ vssd1 vccd1 vccd1 _02642_ sky130_fd_sc_hd__a22o_1
XFILLER_0_175_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11135__B net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08483_ _02523_ _02569_ vssd1 vssd1 vccd1 vccd1 _03612_ sky130_fd_sc_hd__or2_1
XFILLER_0_187_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout155_A _04929_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06229__B net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07434_ top.DUT.register\[20\]\[15\] net563 net512 top.DUT.register\[24\]\[15\] _02572_
+ vssd1 vssd1 vccd1 vccd1 _02573_ sky130_fd_sc_hd__a221o_1
XFILLER_0_190_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_102_1975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_170_3000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07365_ top.DUT.register\[1\]\[8\] net755 net747 top.DUT.register\[17\]\[8\] vssd1
+ vssd1 vccd1 vccd1 _02504_ sky130_fd_sc_hd__a22o_1
XANTENNA__10466__S net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1064_A net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06516__Y _01655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09104_ _02357_ _04149_ _04178_ vssd1 vssd1 vccd1 vccd1 _04179_ sky130_fd_sc_hd__a21oi_1
X_06316_ _01447_ _01469_ vssd1 vssd1 vccd1 vccd1 _01470_ sky130_fd_sc_hd__nor2_1
XFILLER_0_33_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_640 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07296_ top.DUT.register\[6\]\[12\] net567 net559 top.DUT.register\[2\]\[12\] vssd1
+ vssd1 vccd1 vccd1 _02435_ sky130_fd_sc_hd__a22o_1
X_09035_ _02220_ _02751_ _02945_ _03041_ vssd1 vssd1 vccd1 vccd1 _04110_ sky130_fd_sc_hd__or4_1
XFILLER_0_5_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06247_ net1117 net852 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedData\[8\] sky130_fd_sc_hd__and2_1
XFILLER_0_130_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_2474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12346__A2 net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09747__B1 net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold330 top.DUT.register\[31\]\[24\] vssd1 vssd1 vccd1 vccd1 net1446 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10357__A1 net156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold341 top.DUT.register\[1\]\[12\] vssd1 vssd1 vccd1 vccd1 net1457 sky130_fd_sc_hd__dlygate4sd3_1
X_06178_ _01419_ vssd1 vssd1 vccd1 vccd1 _01420_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout691_A net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold352 top.DUT.register\[8\]\[8\] vssd1 vssd1 vccd1 vccd1 net1468 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold363 top.DUT.register\[23\]\[18\] vssd1 vssd1 vccd1 vccd1 net1479 sky130_fd_sc_hd__dlygate4sd3_1
Xhold374 top.DUT.register\[9\]\[27\] vssd1 vssd1 vccd1 vccd1 net1490 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_159_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold385 top.DUT.register\[11\]\[13\] vssd1 vssd1 vccd1 vccd1 net1501 sky130_fd_sc_hd__dlygate4sd3_1
Xhold396 top.DUT.register\[6\]\[19\] vssd1 vssd1 vccd1 vccd1 net1512 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09990__S net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout810 net812 vssd1 vssd1 vccd1 vccd1 net810 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07773__A2 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout821 net822 vssd1 vssd1 vccd1 vccd1 net821 sky130_fd_sc_hd__buf_2
Xfanout832 _01499_ vssd1 vssd1 vccd1 vccd1 net832 sky130_fd_sc_hd__buf_2
X_09937_ _04940_ _04941_ vssd1 vssd1 vccd1 vccd1 _04942_ sky130_fd_sc_hd__xnor2_1
Xfanout843 net844 vssd1 vssd1 vccd1 vccd1 net843 sky130_fd_sc_hd__buf_2
XANTENNA_fanout577_X net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout854 net855 vssd1 vssd1 vccd1 vccd1 net854 sky130_fd_sc_hd__buf_2
XANTENNA_fanout956_A net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06981__B1 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout865 net866 vssd1 vssd1 vccd1 vccd1 net865 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout876 net877 vssd1 vssd1 vccd1 vccd1 net876 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_181_3162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout887 top.busy_o vssd1 vssd1 vccd1 vccd1 net887 sky130_fd_sc_hd__buf_2
X_09868_ top.pc\[24\] _04543_ _04871_ vssd1 vssd1 vccd1 vccd1 _04879_ sky130_fd_sc_hd__a21o_1
Xfanout898 net899 vssd1 vssd1 vccd1 vccd1 net898 sky130_fd_sc_hd__clkbuf_2
Xhold1030 top.ramaddr\[18\] vssd1 vssd1 vccd1 vccd1 net2146 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07525__A2 net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13079__RESET_B net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1041 top.DUT.register\[6\]\[0\] vssd1 vssd1 vccd1 vccd1 net2157 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07363__X _02502_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1052 top.DUT.register\[26\]\[26\] vssd1 vssd1 vccd1 vccd1 net2168 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08722__B2 net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08819_ net883 top.pc\[25\] net694 _03932_ vssd1 vssd1 vccd1 vccd1 _03933_ sky130_fd_sc_hd__a22o_1
Xhold1063 top.DUT.register\[7\]\[14\] vssd1 vssd1 vccd1 vccd1 net2179 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1074 top.DUT.register\[29\]\[24\] vssd1 vssd1 vccd1 vccd1 net2190 sky130_fd_sc_hd__dlygate4sd3_1
X_09799_ top.pc\[18\] _04453_ vssd1 vssd1 vccd1 vccd1 _04817_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout744_X net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1085 top.DUT.register\[20\]\[11\] vssd1 vssd1 vccd1 vccd1 net2201 sky130_fd_sc_hd__dlygate4sd3_1
X_11830_ _05687_ _05712_ vssd1 vssd1 vccd1 vccd1 _05713_ sky130_fd_sc_hd__xor2_2
Xhold1096 top.DUT.register\[27\]\[17\] vssd1 vssd1 vccd1 vccd1 net2212 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_169_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11761_ _05623_ _05629_ _05640_ _05641_ vssd1 vssd1 vccd1 vccd1 _05644_ sky130_fd_sc_hd__a211o_1
X_13500_ clknet_leaf_2_clk _01092_ net914 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[31\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10712_ net1844 net224 net337 vssd1 vssd1 vccd1 vccd1 _00873_ sky130_fd_sc_hd__mux2_1
X_11692_ _05574_ vssd1 vssd1 vccd1 vccd1 _05575_ sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_4_3__f_clk_X clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13431_ clknet_leaf_2_clk _01023_ net918 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[29\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10643_ net197 net2101 net343 vssd1 vssd1 vccd1 vccd1 _00807_ sky130_fd_sc_hd__mux2_1
XANTENNA__10376__S net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_181_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12643__RESET_B net1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13362_ clknet_leaf_23_clk _00954_ net1022 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[27\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06155__A top.a1.dataIn\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10574_ net2201 net219 net350 vssd1 vssd1 vccd1 vccd1 _00740_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_5_clk_A clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12313_ _06118_ _06119_ vssd1 vssd1 vccd1 vccd1 _01356_ sky130_fd_sc_hd__nor2_1
XFILLER_0_23_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_210_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13293_ clknet_leaf_50_clk _00885_ net1058 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[24\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_121_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_161_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12244_ net1227 _06075_ _06077_ vssd1 vssd1 vccd1 vccd1 _01323_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_210_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_75_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12175_ net1238 net846 net796 _05978_ vssd1 vssd1 vccd1 vccd1 _01283_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_166_2935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11126_ net906 net1296 net861 _05068_ vssd1 vssd1 vccd1 vccd1 _01214_ sky130_fd_sc_hd__a31o_1
X_11057_ net103 net868 _05045_ net1292 vssd1 vssd1 vccd1 vccd1 _01168_ sky130_fd_sc_hd__a22o_1
XFILLER_0_64_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10008_ net158 net2084 net624 vssd1 vssd1 vccd1 vccd1 _00213_ sky130_fd_sc_hd__mux2_1
XANTENNA__07714__A top.a1.instruction\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_199_3434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06724__B1 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_2031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_106_2042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11236__A top.lcd.nextState\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_204_777 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_148_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11959_ _05794_ _05822_ vssd1 vssd1 vccd1 vccd1 _05842_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10284__A0 top.DUT.register\[11\]\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13629_ clknet_leaf_72_clk _01216_ net1085 vssd1 vssd1 vccd1 vccd1 net56 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10286__S net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07150_ top.DUT.register\[20\]\[11\] net663 net750 top.DUT.register\[26\]\[11\] _02288_
+ vssd1 vssd1 vccd1 vccd1 _02289_ sky130_fd_sc_hd__a221o_1
XFILLER_0_27_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07081_ _02198_ _02219_ vssd1 vssd1 vccd1 vccd1 _02220_ sky130_fd_sc_hd__nor2_2
XFILLER_0_42_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09729__B1 net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_454 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_2393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07755__A2 net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08952__B2 net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_14__f_clk_X clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07983_ net333 vssd1 vssd1 vccd1 vccd1 _03122_ sky130_fd_sc_hd__inv_2
Xfanout139 _04207_ vssd1 vssd1 vccd1 vccd1 net139 sky130_fd_sc_hd__clkbuf_2
XANTENNA__06963__B1 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09722_ _02341_ _04149_ _04177_ vssd1 vssd1 vccd1 vccd1 _04750_ sky130_fd_sc_hd__and3_1
X_06934_ top.DUT.register\[24\]\[21\] net646 net735 top.DUT.register\[16\]\[21\] _02072_
+ vssd1 vssd1 vccd1 vccd1 _02073_ sky130_fd_sc_hd__a221o_1
XFILLER_0_198_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07507__A2 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09653_ _04675_ _04680_ vssd1 vssd1 vccd1 vccd1 _04694_ sky130_fd_sc_hd__nor2_1
X_06865_ _02003_ vssd1 vssd1 vccd1 vccd1 _02004_ sky130_fd_sc_hd__inv_2
XANTENNA__10511__A1 net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08604_ _03701_ _03726_ _02611_ vssd1 vssd1 vccd1 vccd1 _03727_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_179_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09584_ _04629_ _04630_ vssd1 vssd1 vccd1 vccd1 _04631_ sky130_fd_sc_hd__nor2_1
X_06796_ top.DUT.register\[6\]\[17\] net568 net536 top.DUT.register\[19\]\[17\] vssd1
+ vssd1 vccd1 vccd1 _01935_ sky130_fd_sc_hd__a22o_1
XFILLER_0_210_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_118_Right_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_179_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08535_ net423 _03642_ _03661_ net496 vssd1 vssd1 vccd1 vccd1 _03662_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_46_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout537_A net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08466_ net1874 net833 net803 _03595_ vssd1 vssd1 vccd1 vccd1 _00027_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_34_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07140__B1 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_137_2503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07417_ top.DUT.register\[5\]\[9\] net651 net639 top.DUT.register\[8\]\[9\] _02554_
+ vssd1 vssd1 vccd1 vccd1 _02556_ sky130_fd_sc_hd__a221o_1
XANTENNA__11152__Y _05082_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_190_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_162_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06494__A2 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08397_ net304 _03426_ vssd1 vssd1 vccd1 vccd1 _03529_ sky130_fd_sc_hd__or2_2
XFILLER_0_161_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout704_A _01642_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout325_X net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09985__S net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07348_ _02480_ _02482_ _02484_ _02486_ vssd1 vssd1 vccd1 vccd1 _02487_ sky130_fd_sc_hd__or4_1
XANTENNA__10578__A1 net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_150_2703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10924__S net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07279_ top.DUT.register\[30\]\[13\] net760 net641 top.DUT.register\[8\]\[13\] vssd1
+ vssd1 vccd1 vccd1 _02418_ sky130_fd_sc_hd__a22o_1
XFILLER_0_60_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09018_ _03889_ _03982_ _04006_ _04092_ vssd1 vssd1 vccd1 vccd1 _04093_ sky130_fd_sc_hd__or4_1
XFILLER_0_130_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10290_ net1899 net161 net387 vssd1 vssd1 vccd1 vccd1 _00468_ sky130_fd_sc_hd__mux2_1
XANTENNA__09196__A1 _01505_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_478 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold160 top.ramstore\[0\] vssd1 vssd1 vccd1 vccd1 net1276 sky130_fd_sc_hd__dlygate4sd3_1
Xhold171 top.DUT.register\[26\]\[4\] vssd1 vssd1 vccd1 vccd1 net1287 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06422__B top.a1.instruction\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold182 top.ramaddr\[23\] vssd1 vssd1 vccd1 vccd1 net1298 sky130_fd_sc_hd__dlygate4sd3_1
Xhold193 top.DUT.register\[15\]\[0\] vssd1 vssd1 vccd1 vccd1 net1309 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07746__A2 net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout861_X net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout640 _01619_ vssd1 vssd1 vccd1 vccd1 net640 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06954__B1 net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout651 _01610_ vssd1 vssd1 vccd1 vccd1 net651 sky130_fd_sc_hd__clkbuf_8
Xfanout662 _01606_ vssd1 vssd1 vccd1 vccd1 net662 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_148_2665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout673 net674 vssd1 vssd1 vccd1 vccd1 net673 sky130_fd_sc_hd__clkbuf_8
Xfanout684 _01510_ vssd1 vssd1 vccd1 vccd1 net684 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_70_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07093__X _02232_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout695 net696 vssd1 vssd1 vccd1 vccd1 net695 sky130_fd_sc_hd__clkbuf_2
X_12931_ clknet_leaf_57_clk _00523_ net1076 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[13\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06706__B1 net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_161_2854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_161_2865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12862_ clknet_leaf_20_clk _00454_ net1028 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[11\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_34_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_201_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11813_ _05625_ _05665_ vssd1 vssd1 vccd1 vccd1 _05696_ sky130_fd_sc_hd__or2_1
XANTENNA__11058__A2 net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12793_ clknet_leaf_15_clk _00385_ net961 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[9\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_205_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_194_3353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11744_ _01399_ _05620_ _05585_ vssd1 vssd1 vccd1 vccd1 _05627_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_55_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07131__B1 net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11675_ _05528_ _05549_ vssd1 vssd1 vccd1 vccd1 _05558_ sky130_fd_sc_hd__nand2_1
XFILLER_0_71_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_12_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13414_ clknet_leaf_40_clk _01006_ net1053 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[28\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_181_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_107 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10626_ net148 net2002 net348 vssd1 vssd1 vccd1 vccd1 _00791_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_77_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_180_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13345_ clknet_leaf_16_clk _00937_ net965 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[26\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_10557_ net2159 net159 net355 vssd1 vssd1 vccd1 vccd1 _00724_ sky130_fd_sc_hd__mux2_1
XANTENNA__10834__S net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_180_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07985__A2 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13276_ clknet_leaf_0_clk _00868_ net922 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[24\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_10488_ net2210 net168 net361 vssd1 vssd1 vccd1 vccd1 _00658_ sky130_fd_sc_hd__mux2_1
X_12227_ _01383_ _06066_ vssd1 vssd1 vccd1 vccd1 _06067_ sky130_fd_sc_hd__nand2_1
XFILLER_0_166_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12158_ _06038_ _06039_ _01403_ _06036_ vssd1 vssd1 vccd1 vccd1 _06041_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__06945__B1 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11109_ net45 net869 vssd1 vssd1 vccd1 vccd1 _05060_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_16_Left_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12089_ _05941_ _05971_ vssd1 vssd1 vccd1 vccd1 _05972_ sky130_fd_sc_hd__xor2_2
XANTENNA__11237__Y _05130_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11297__A2 _05136_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_182_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06650_ _01786_ _01788_ vssd1 vssd1 vccd1 vccd1 _01789_ sky130_fd_sc_hd__or2_1
XFILLER_0_189_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07370__B1 net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06581_ _01713_ _01715_ _01717_ _01719_ vssd1 vssd1 vccd1 vccd1 _01720_ sky130_fd_sc_hd__or4_1
XFILLER_0_188_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08320_ net498 _03446_ _03454_ net434 vssd1 vssd1 vccd1 vccd1 _03455_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_19_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_50_clk_X clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07122__B1 net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06347__X _01489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08275__A net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_145_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08251_ net321 net436 _03387_ _03386_ vssd1 vssd1 vccd1 vccd1 _03388_ sky130_fd_sc_hd__a31o_1
XFILLER_0_74_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_25_Left_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_119_2233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07202_ net795 _02331_ _02335_ _02339_ vssd1 vssd1 vccd1 vccd1 _02341_ sky130_fd_sc_hd__or4_1
XFILLER_0_61_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08182_ _03316_ _03319_ net288 vssd1 vssd1 vccd1 vccd1 _03320_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_41_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07133_ top.DUT.register\[14\]\[11\] net583 net547 top.DUT.register\[18\]\[11\] vssd1
+ vssd1 vccd1 vccd1 _02272_ sky130_fd_sc_hd__a22o_1
XFILLER_0_144_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10744__S net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09818__B _04487_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_2422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_2433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07976__A2 net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07064_ top.DUT.register\[30\]\[22\] net759 net750 top.DUT.register\[26\]\[22\] vssd1
+ vssd1 vccd1 vccd1 _02203_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_12_Right_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06242__B net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12182__B1 net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07728__A2 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_34_Left_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09553__B _04590_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07966_ top.DUT.register\[19\]\[31\] net538 net526 top.DUT.register\[11\]\[31\] vssd1
+ vssd1 vccd1 vccd1 _03105_ sky130_fd_sc_hd__a22o_1
X_09705_ _03460_ net405 net490 _04736_ vssd1 vssd1 vccd1 vccd1 _04737_ sky130_fd_sc_hd__o211a_4
X_06917_ top.DUT.register\[16\]\[21\] net544 net445 top.DUT.register\[1\]\[21\] _02055_
+ vssd1 vssd1 vccd1 vccd1 _02056_ sky130_fd_sc_hd__a221o_1
XFILLER_0_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07897_ top.DUT.register\[6\]\[1\] net569 net545 top.DUT.register\[16\]\[1\] _03035_
+ vssd1 vssd1 vccd1 vccd1 _03036_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout654_A _01610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_94_clk clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_94_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_179_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09636_ top.pad.keyCode\[1\] top.pad.keyCode\[2\] top.pad.keyCode\[3\] top.pad.keyCode\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04678_ sky130_fd_sc_hd__or4b_2
X_06848_ top.DUT.register\[23\]\[19\] net673 net740 top.DUT.register\[12\]\[19\] vssd1
+ vssd1 vccd1 vccd1 _01987_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_21_Right_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_143_2584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_2595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09567_ top.pc\[29\] _04605_ vssd1 vssd1 vccd1 vccd1 _04615_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout442_X net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06779_ _01897_ _01917_ vssd1 vssd1 vccd1 vccd1 _01918_ sky130_fd_sc_hd__nor2_1
XANTENNA__10919__S net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_251 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08518_ net317 _03644_ _03643_ vssd1 vssd1 vccd1 vccd1 _03645_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_93_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08185__A _01572_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_43_Left_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09498_ _04536_ _04542_ _04550_ _04051_ top.pc\[24\] vssd1 vssd1 vccd1 vccd1 _00104_
+ sky130_fd_sc_hd__o32a_1
XANTENNA__07113__B1 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_176_3083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_148_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08449_ _03332_ _03578_ net297 vssd1 vssd1 vccd1 vccd1 _03579_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_175_492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_479 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout707_X net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11460_ _05302_ _05337_ vssd1 vssd1 vccd1 vccd1 _05343_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_163_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08913__A _01659_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_5_0_clk_X clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10411_ net1460 net198 net372 vssd1 vssd1 vccd1 vccd1 _00583_ sky130_fd_sc_hd__mux2_1
X_11391_ _05242_ _05268_ vssd1 vssd1 vccd1 vccd1 _05274_ sky130_fd_sc_hd__xnor2_2
XANTENNA__10654__S net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_30_Right_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_59_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13130_ clknet_leaf_116_clk _00722_ net958 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[19\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07967__A2 net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10342_ net1614 net208 net379 vssd1 vssd1 vccd1 vccd1 _00518_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06433__A _01571_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13061_ clknet_leaf_35_clk _00653_ net1041 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[17\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_10273_ net2253 net227 net385 vssd1 vssd1 vccd1 vccd1 _00451_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_52_Left_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07248__B _02385_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08916__A1 net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12012_ _05874_ _05887_ vssd1 vssd1 vccd1 vccd1 _05895_ sky130_fd_sc_hd__xnor2_1
XANTENNA__08916__B2 _03259_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06927__B1 net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout470 _01524_ vssd1 vssd1 vccd1 vccd1 net470 sky130_fd_sc_hd__clkbuf_8
Xfanout481 _04964_ vssd1 vssd1 vccd1 vccd1 net481 sky130_fd_sc_hd__buf_4
XANTENNA__11279__A2 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout492 _03339_ vssd1 vssd1 vccd1 vccd1 net492 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_45_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_85_clk clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_85_clk
+ sky130_fd_sc_hd__clkbuf_8
X_12914_ clknet_leaf_23_clk _00506_ net1021 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[13\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_17_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12845_ clknet_leaf_42_clk _00437_ net1064 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[10\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_186_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_61_Left_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10829__S net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07270__Y _02409_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07711__B _02849_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12776_ clknet_leaf_7_clk _00368_ net946 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[8\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08095__A _02773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07104__B1 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11727_ _05606_ _05607_ vssd1 vssd1 vccd1 vccd1 _05610_ sky130_fd_sc_hd__nor2_1
XANTENNA__11233__B top.lcd.nextState\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11658_ _05495_ _05540_ vssd1 vssd1 vccd1 vccd1 _05541_ sky130_fd_sc_hd__nor2_1
XANTENNA__09919__A net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_211_3607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_211_3618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10609_ net208 net1976 net348 vssd1 vssd1 vccd1 vccd1 _00774_ sky130_fd_sc_hd__mux2_1
XFILLER_0_141_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_211_3629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10564__S net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11589_ _05436_ _05471_ vssd1 vssd1 vccd1 vccd1 _05472_ sky130_fd_sc_hd__or2_1
XFILLER_0_141_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold907 top.DUT.register\[13\]\[7\] vssd1 vssd1 vccd1 vccd1 net2023 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold918 top.DUT.register\[4\]\[23\] vssd1 vssd1 vccd1 vccd1 net2034 sky130_fd_sc_hd__dlygate4sd3_1
X_13328_ clknet_leaf_29_clk _00920_ net1018 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[25\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold929 top.DUT.register\[10\]\[7\] vssd1 vssd1 vccd1 vccd1 net2045 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_70_Left_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_114_2152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10962__A1 net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_114_2163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13259_ clknet_leaf_45_clk _00851_ net1065 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[23\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06630__A2 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_209_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_208_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06918__B1 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10714__A1 net206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07820_ top.DUT.register\[23\]\[0\] net671 net711 top.DUT.register\[11\]\[0\] _02958_
+ vssd1 vssd1 vccd1 vccd1 _02959_ sky130_fd_sc_hd__a221o_1
XANTENNA__08383__A2 net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09580__A1 _01679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_208_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07591__B1 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09941__X _04946_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12600__CLK clknet_leaf_128_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07751_ top.DUT.register\[15\]\[3\] net681 net677 top.DUT.register\[31\]\[3\] vssd1
+ vssd1 vccd1 vccd1 _02890_ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_92_clk_A clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_76_clk clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_76_clk
+ sky130_fd_sc_hd__clkbuf_8
X_06702_ top.DUT.register\[23\]\[25\] net571 net564 top.DUT.register\[20\]\[25\] vssd1
+ vssd1 vccd1 vccd1 _01841_ sky130_fd_sc_hd__a22o_1
XANTENNA__09332__A1 net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07682_ top.DUT.register\[16\]\[4\] net735 _02818_ _02820_ vssd1 vssd1 vccd1 vccd1
+ _02821_ sky130_fd_sc_hd__a211o_1
XANTENNA__07343__B1 net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09421_ top.pc\[20\] _04461_ vssd1 vssd1 vccd1 vccd1 _04478_ sky130_fd_sc_hd__and2_1
X_06633_ top.DUT.register\[12\]\[27\] net740 net735 top.DUT.register\[16\]\[27\] _01771_
+ vssd1 vssd1 vccd1 vccd1 _01772_ sky130_fd_sc_hd__a221o_1
XANTENNA__07902__A net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_177_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06697__A2 net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_177_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10739__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09352_ _04398_ _04399_ _04396_ vssd1 vssd1 vccd1 vccd1 _04413_ sky130_fd_sc_hd__o21bai_1
X_06564_ top.DUT.register\[18\]\[28\] net549 net514 top.DUT.register\[24\]\[28\] vssd1
+ vssd1 vccd1 vccd1 _01703_ sky130_fd_sc_hd__a22o_1
XFILLER_0_176_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06518__A _01571_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_210 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08303_ _03203_ _03212_ net314 vssd1 vssd1 vccd1 vccd1 _03438_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09283_ top.pc\[12\] _04336_ vssd1 vssd1 vccd1 vccd1 _04348_ sky130_fd_sc_hd__or2_1
XFILLER_0_142_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06495_ top.DUT.register\[4\]\[30\] net669 net732 top.DUT.register\[14\]\[30\] _01631_
+ vssd1 vssd1 vccd1 vccd1 _01634_ sky130_fd_sc_hd__a221o_1
XANTENNA__06237__B net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout235_A _04757_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_191_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08234_ net303 net333 vssd1 vssd1 vccd1 vccd1 _03371_ sky130_fd_sc_hd__nand2_2
XANTENNA_clkbuf_leaf_30_clk_A clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13106__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08165_ _02069_ net301 vssd1 vssd1 vccd1 vccd1 _03303_ sky130_fd_sc_hd__nand2_1
XANTENNA__10474__S net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_803 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07116_ top.DUT.register\[4\]\[16\] net668 net703 top.DUT.register\[3\]\[16\] _02251_
+ vssd1 vssd1 vccd1 vccd1 _02255_ sky130_fd_sc_hd__a221o_1
X_08096_ _03233_ _03234_ vssd1 vssd1 vccd1 vccd1 _03235_ sky130_fd_sc_hd__and2_1
XFILLER_0_42_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkload80 clknet_leaf_42_clk vssd1 vssd1 vccd1 vccd1 clkload80/Y sky130_fd_sc_hd__bufinv_16
XANTENNA_clkbuf_leaf_45_clk_A clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06621__A2 net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07047_ top.DUT.register\[13\]\[22\] net463 net504 top.DUT.register\[27\]\[22\] vssd1
+ vssd1 vccd1 vccd1 _02186_ sky130_fd_sc_hd__a22o_1
Xclkload91 clknet_leaf_78_clk vssd1 vssd1 vccd1 vccd1 clkload91/Y sky130_fd_sc_hd__inv_8
XANTENNA_fanout392_X net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout771_A _01614_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout869_A _01427_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08998_ net284 _03420_ _03477_ vssd1 vssd1 vccd1 vccd1 _04073_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07582__B1 net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_2624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07949_ _02267_ _03073_ _03086_ _03087_ vssd1 vssd1 vccd1 vccd1 _03088_ sky130_fd_sc_hd__o211a_1
XFILLER_0_203_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout657_X net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_170_Right_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_103_clk_A clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10960_ top.edg2.flip2 _05002_ top.edg2.flip1 vssd1 vssd1 vccd1 vccd1 _05003_ sky130_fd_sc_hd__nor3b_1
XTAP_TAPCELL_ROW_3_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_178_3112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11130__A1 net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_178_3123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09874__A2 net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06688__A2 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09619_ top.a1.state\[0\] top.a1.state\[2\] top.a1.state\[1\] vssd1 vssd1 vccd1 vccd1
+ _04664_ sky130_fd_sc_hd__nor3b_2
XANTENNA__10649__S net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10891_ net1358 net262 net480 vssd1 vssd1 vccd1 vccd1 _01052_ sky130_fd_sc_hd__mux2_1
XFILLER_0_167_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12630_ clknet_leaf_4_clk _00222_ net937 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[4\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_183_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_191_3312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_183_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_418 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_118_clk_A clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12561_ clknet_leaf_116_clk _00153_ net957 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[2\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_66_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_416 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11512_ _05351_ _05394_ vssd1 vssd1 vccd1 vccd1 _05395_ sky130_fd_sc_hd__nand2_1
XFILLER_0_93_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_760 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_451 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12492_ clknet_leaf_86_clk _00084_ net1006 vssd1 vssd1 vccd1 vccd1 top.pc\[4\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_108_367 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_156_2786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_191_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11443_ _05287_ net278 top.a1.dataIn\[17\] vssd1 vssd1 vccd1 vccd1 _05326_ sky130_fd_sc_hd__a21oi_1
XANTENNA__06860__A2 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10384__S net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_202_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11374_ _05249_ _05250_ _05224_ vssd1 vssd1 vccd1 vccd1 _05257_ sky130_fd_sc_hd__a21boi_1
XANTENNA__06163__A top.pc\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_189_3274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13204__RESET_B net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13113_ clknet_leaf_16_clk _00705_ net960 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[19\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_104_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10325_ net155 net1496 net383 vssd1 vssd1 vccd1 vccd1 _00502_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_189_3285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06612__A2 net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13044_ clknet_leaf_54_clk _00636_ net1075 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[17\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_10256_ net166 net1514 net391 vssd1 vssd1 vccd1 vccd1 _00435_ sky130_fd_sc_hd__mux2_1
XANTENNA__06450__X _01589_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12623__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08952__A2_N _04050_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10187_ top.a1.instruction\[7\] top.a1.instruction\[8\] _04154_ net786 vssd1 vssd1
+ vccd1 vccd1 _04967_ sky130_fd_sc_hd__or4b_1
XANTENNA__07573__B1 net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_58_clk clknet_4_12__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_58_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_72_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07325__B1 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_204_3499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06679__A2 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10559__S net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_768 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12828_ clknet_leaf_130_clk _00420_ net909 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[10\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_174_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12759_ clknet_leaf_128_clk _00351_ net912 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[8\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06280_ top.lcd.cnt_500hz\[5\] top.lcd.cnt_500hz\[8\] _01438_ vssd1 vssd1 vccd1 vccd1
+ _01443_ sky130_fd_sc_hd__or3b_1
XFILLER_0_142_602 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06851__A2 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10294__S net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold704 top.DUT.register\[28\]\[16\] vssd1 vssd1 vccd1 vccd1 net1820 sky130_fd_sc_hd__dlygate4sd3_1
Xhold715 top.DUT.register\[19\]\[6\] vssd1 vssd1 vccd1 vccd1 net1831 sky130_fd_sc_hd__dlygate4sd3_1
Xhold726 top.DUT.register\[5\]\[7\] vssd1 vssd1 vccd1 vccd1 net1842 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold737 top.DUT.register\[10\]\[25\] vssd1 vssd1 vccd1 vccd1 net1853 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_96_1888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06504__C _01607_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06603__A2 _01741_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09970_ net2193 net169 net627 vssd1 vssd1 vccd1 vccd1 _00178_ sky130_fd_sc_hd__mux2_1
Xhold748 top.DUT.register\[28\]\[25\] vssd1 vssd1 vccd1 vccd1 net1864 sky130_fd_sc_hd__dlygate4sd3_1
Xhold759 top.DUT.register\[29\]\[21\] vssd1 vssd1 vccd1 vccd1 net1875 sky130_fd_sc_hd__dlygate4sd3_1
X_08921_ net695 _04028_ _04029_ top.pc\[30\] net884 vssd1 vssd1 vccd1 vccd1 _04030_
+ sky130_fd_sc_hd__a32o_1
XANTENNA__06360__X _01499_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06801__A _01930_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08356__A2 net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08852_ net435 _03960_ _03963_ _03264_ vssd1 vssd1 vccd1 vccd1 _03964_ sky130_fd_sc_hd__o2bb2a_1
X_07803_ top.DUT.register\[25\]\[2\] net455 net511 top.DUT.register\[24\]\[2\] _02941_
+ vssd1 vssd1 vccd1 vccd1 _02942_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_108_Left_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08783_ _03200_ _03207_ vssd1 vssd1 vccd1 vccd1 _03898_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_127_2354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_49_clk clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_49_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_137_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07734_ top.DUT.register\[8\]\[3\] net641 net757 top.DUT.register\[1\]\[3\] vssd1
+ vssd1 vccd1 vccd1 _02873_ sky130_fd_sc_hd__a22o_1
XANTENNA__07316__B1 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11112__A1 net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08728__A net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10469__S net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07665_ top.a1.instruction\[11\] _01474_ vssd1 vssd1 vccd1 vccd1 _02804_ sky130_fd_sc_hd__and2_1
XFILLER_0_149_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout352_A net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_140_2543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09404_ top.pc\[18\] _04428_ top.pc\[19\] vssd1 vssd1 vccd1 vccd1 _04462_ sky130_fd_sc_hd__a21oi_1
X_06616_ top.DUT.register\[15\]\[27\] net682 net678 top.DUT.register\[31\]\[27\] vssd1
+ vssd1 vccd1 vccd1 _01755_ sky130_fd_sc_hd__a22o_1
XFILLER_0_153_72 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07596_ top.DUT.register\[14\]\[6\] net730 net702 top.DUT.register\[3\]\[6\] vssd1
+ vssd1 vccd1 vccd1 _02735_ sky130_fd_sc_hd__a22o_1
XFILLER_0_94_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_149_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_192_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09335_ top.pc\[15\] _04386_ vssd1 vssd1 vccd1 vccd1 _04397_ sky130_fd_sc_hd__nor2_1
X_06547_ top.DUT.register\[8\]\[29\] net641 net752 top.DUT.register\[26\]\[29\] _01680_
+ vssd1 vssd1 vccd1 vccd1 _01686_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_173_3042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout617_A _04954_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08292__A1 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_192_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09266_ _04313_ _04314_ _04316_ vssd1 vssd1 vccd1 vccd1 _04332_ sky130_fd_sc_hd__a21o_1
XANTENNA__07095__A2 net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06478_ net788 _01607_ _01611_ vssd1 vssd1 vccd1 vccd1 _01617_ sky130_fd_sc_hd__and3_4
XFILLER_0_35_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_173_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08217_ net2018 net830 net800 _03354_ vssd1 vssd1 vccd1 vccd1 _00019_ sky130_fd_sc_hd__a22o_1
XANTENNA__06842__A2 net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09197_ net899 top.pc\[6\] _04253_ _04267_ net892 vssd1 vssd1 vccd1 vccd1 _00086_
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_172_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout405_X net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09993__S net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08148_ _02849_ net330 vssd1 vssd1 vccd1 vccd1 _03286_ sky130_fd_sc_hd__nand2_1
XANTENNA__09846__X _04859_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12646__CLK clknet_leaf_40_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout986_A net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09792__A1 _04438_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08079_ _02242_ net299 vssd1 vssd1 vccd1 vccd1 _03218_ sky130_fd_sc_hd__nand2_1
XANTENNA__09792__B2 top.a1.dataIn\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10932__S net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10110_ net1811 net148 net613 vssd1 vssd1 vccd1 vccd1 _00311_ sky130_fd_sc_hd__mux2_1
XANTENNA__07807__A _02925_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11090_ net906 net1915 net861 _05050_ vssd1 vssd1 vccd1 vccd1 _01196_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_8_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout774_X net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10041_ net1333 net159 net621 vssd1 vssd1 vccd1 vccd1 _00244_ sky130_fd_sc_hd__mux2_1
XANTENNA_hold185_X net1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold20 top.ramstore\[30\] vssd1 vssd1 vccd1 vccd1 net1136 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07555__B1 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold31 top.ramstore\[29\] vssd1 vssd1 vccd1 vccd1 net1147 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09581__X _04628_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold42 top.a1.row1\[115\] vssd1 vssd1 vccd1 vccd1 net1158 sky130_fd_sc_hd__dlygate4sd3_1
Xhold53 top.a1.row1\[106\] vssd1 vssd1 vccd1 vccd1 net1169 sky130_fd_sc_hd__dlygate4sd3_1
Xhold64 net75 vssd1 vssd1 vccd1 vccd1 net1180 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_203_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold75 net113 vssd1 vssd1 vccd1 vccd1 net1191 sky130_fd_sc_hd__dlygate4sd3_1
Xhold86 top.ramstore\[12\] vssd1 vssd1 vccd1 vccd1 net1202 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_203_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13800_ clknet_leaf_70_clk _01369_ net1086 vssd1 vssd1 vccd1 vccd1 top.pad.keyCode\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold97 top.a1.row1\[0\] vssd1 vssd1 vccd1 vccd1 net1213 sky130_fd_sc_hd__dlygate4sd3_1
X_11992_ _05828_ _05840_ _05851_ _05827_ vssd1 vssd1 vccd1 vccd1 _05875_ sky130_fd_sc_hd__o31a_1
XFILLER_0_97_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07307__B1 net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13731_ clknet_leaf_96_clk _01302_ vssd1 vssd1 vccd1 vccd1 top.a1.dataInTemp\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_10943_ net1355 net178 net591 vssd1 vssd1 vccd1 vccd1 _01104_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_67_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10379__S net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_543 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_3_0_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_3_0_0_clk sky130_fd_sc_hd__clkbuf_8
X_13662_ clknet_leaf_90_clk _01238_ net1001 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[112\]
+ sky130_fd_sc_hd__dfrtp_1
X_10874_ net203 net1965 net596 vssd1 vssd1 vccd1 vccd1 _01035_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_158_2815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06158__A top.a1.dataIn\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_390 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12613_ clknet_leaf_33_clk _00205_ net1042 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[3\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_13593_ clknet_leaf_63_clk net1167 net1067 vssd1 vssd1 vccd1 vccd1 net85 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_360 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12544_ clknet_leaf_113_clk _00136_ net991 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[1\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06445__X _01584_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07086__A2 net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08373__A _03169_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_624 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12475_ clknet_leaf_47_clk _00070_ net1067 vssd1 vssd1 vccd1 vccd1 top.ramstore\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06833__A2 net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11426_ _05267_ _05275_ _05285_ vssd1 vssd1 vccd1 vccd1 _05309_ sky130_fd_sc_hd__and3_1
XANTENNA__09756__X _04779_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_6 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09783__A1 _04420_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_2111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11357_ top.a1.dataIn\[28\] _05239_ vssd1 vssd1 vccd1 vccd1 _05240_ sky130_fd_sc_hd__xor2_1
XANTENNA__09783__B2 top.a1.dataIn\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10842__S net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07794__B1 net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10308_ net213 net1728 net384 vssd1 vssd1 vccd1 vccd1 _00485_ sky130_fd_sc_hd__mux2_1
X_11288_ net881 _05129_ _05149_ vssd1 vssd1 vccd1 vccd1 _05178_ sky130_fd_sc_hd__o21bai_2
XTAP_TAPCELL_ROW_169_2977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13027_ clknet_leaf_61_clk _00619_ net1089 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[16\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_169_2988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10239_ net233 net2288 net389 vssd1 vssd1 vccd1 vccd1 _00418_ sky130_fd_sc_hd__mux2_1
XANTENNA__07546__B1 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_206_3539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1040 net1043 vssd1 vssd1 vccd1 vccd1 net1040 sky130_fd_sc_hd__clkbuf_4
Xfanout1051 net1052 vssd1 vssd1 vccd1 vccd1 net1051 sky130_fd_sc_hd__clkbuf_4
Xfanout1062 net1070 vssd1 vssd1 vccd1 vccd1 net1062 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07010__A2 net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1073 net1074 vssd1 vssd1 vccd1 vccd1 net1073 sky130_fd_sc_hd__clkbuf_4
Xfanout1084 net1085 vssd1 vssd1 vccd1 vccd1 net1084 sky130_fd_sc_hd__clkbuf_4
Xfanout1095 net1096 vssd1 vssd1 vccd1 vccd1 net1095 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_109_2084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10289__S net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_187_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_202_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_190_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_202_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07450_ _02582_ _02584_ _02586_ _02588_ vssd1 vssd1 vccd1 vccd1 _02589_ sky130_fd_sc_hd__or4_4
XTAP_TAPCELL_ROW_122_2273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_202_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_201_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06401_ _01511_ _01521_ _01527_ vssd1 vssd1 vccd1 vccd1 _01540_ sky130_fd_sc_hd__and3_4
XFILLER_0_45_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07381_ _02515_ _02517_ _02519_ vssd1 vssd1 vccd1 vccd1 _02520_ sky130_fd_sc_hd__or3_1
XFILLER_0_17_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09120_ _02904_ _02944_ vssd1 vssd1 vccd1 vccd1 _04195_ sky130_fd_sc_hd__nand2_1
X_06332_ _01391_ _01392_ vssd1 vssd1 vccd1 vccd1 _01479_ sky130_fd_sc_hd__nor2_2
XANTENNA__07077__A2 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_1917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09051_ _03390_ _03429_ _04063_ _04082_ vssd1 vssd1 vccd1 vccd1 _04126_ sky130_fd_sc_hd__or4_1
XANTENNA__06285__B1 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06263_ top.ramload\[24\] net853 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedData\[24\]
+ sky130_fd_sc_hd__and2_1
XANTENNA__09098__B _04172_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_6_Right_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08002_ _03133_ _03140_ vssd1 vssd1 vccd1 vccd1 _03141_ sky130_fd_sc_hd__nor2_4
XFILLER_0_53_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08026__A1 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold501 top.DUT.register\[18\]\[29\] vssd1 vssd1 vccd1 vccd1 net1617 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06194_ top.ru.state\[4\] net887 net1128 vssd1 vssd1 vccd1 vccd1 _00011_ sky130_fd_sc_hd__a21o_1
XFILLER_0_130_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold512 top.DUT.register\[8\]\[20\] vssd1 vssd1 vccd1 vccd1 net1628 sky130_fd_sc_hd__dlygate4sd3_1
Xhold523 top.DUT.register\[9\]\[11\] vssd1 vssd1 vccd1 vccd1 net1639 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_452 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold534 top.a1.hexop\[4\] vssd1 vssd1 vccd1 vccd1 net1650 sky130_fd_sc_hd__dlygate4sd3_1
Xhold545 top.DUT.register\[15\]\[9\] vssd1 vssd1 vccd1 vccd1 net1661 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10752__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold556 top.pad.button_control.r_counter\[10\] vssd1 vssd1 vccd1 vccd1 net1672 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold567 top.DUT.register\[2\]\[10\] vssd1 vssd1 vccd1 vccd1 net1683 sky130_fd_sc_hd__dlygate4sd3_1
Xhold578 top.DUT.register\[30\]\[9\] vssd1 vssd1 vccd1 vccd1 net1694 sky130_fd_sc_hd__dlygate4sd3_1
X_09953_ net1546 net238 net628 vssd1 vssd1 vccd1 vccd1 _00161_ sky130_fd_sc_hd__mux2_1
Xhold589 top.DUT.register\[28\]\[15\] vssd1 vssd1 vccd1 vccd1 net1705 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08904_ _01702_ _03992_ _01699_ vssd1 vssd1 vccd1 vccd1 _04013_ sky130_fd_sc_hd__a21oi_2
XTAP_TAPCELL_ROW_5_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06250__B net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09884_ _04151_ _04891_ _04893_ vssd1 vssd1 vccd1 vccd1 _04894_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07537__B1 net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07001__A2 net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08835_ _03093_ _03947_ vssd1 vssd1 vccd1 vccd1 _03948_ sky130_fd_sc_hd__nor2_1
XFILLER_0_99_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout567_A _01525_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08766_ _02136_ net492 vssd1 vssd1 vccd1 vccd1 _03882_ sky130_fd_sc_hd__nor2_1
XFILLER_0_79_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08458__A net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07717_ _02359_ _02805_ _02855_ vssd1 vssd1 vccd1 vccd1 _02856_ sky130_fd_sc_hd__a21o_1
XFILLER_0_79_143 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10199__S net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08697_ _03814_ _03815_ vssd1 vssd1 vccd1 vccd1 _03816_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout734_A net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout355_X net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1097_X net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09988__S net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07648_ top.DUT.register\[4\]\[5\] net667 net758 top.DUT.register\[30\]\[5\] _02783_
+ vssd1 vssd1 vccd1 vccd1 _02787_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_24_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06409__C _01546_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07579_ top.DUT.register\[20\]\[6\] net563 net559 top.DUT.register\[2\]\[6\] vssd1
+ vssd1 vccd1 vccd1 _02718_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout522_X net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10927__S _04972_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout901_A net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08905__B _04013_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_180_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09318_ top.pc\[14\] _04370_ vssd1 vssd1 vccd1 vccd1 _04381_ sky130_fd_sc_hd__and2_1
XANTENNA__07068__A2 net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10590_ net1847 net159 net352 vssd1 vssd1 vccd1 vccd1 _00756_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_62_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09249_ _02547_ top.pc\[10\] vssd1 vssd1 vccd1 vccd1 _04316_ sky130_fd_sc_hd__and2b_1
XANTENNA__06815__A2 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_153_2734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_153_2745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12260_ top.lcd.cnt_500hz\[1\] top.lcd.cnt_500hz\[0\] vssd1 vssd1 vccd1 vccd1 _06087_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_90_396 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11211_ net845 _05028_ _05038_ vssd1 vssd1 vccd1 vccd1 _05112_ sky130_fd_sc_hd__and3_1
XANTENNA__09765__A1 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08568__A2 net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10662__S net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12191_ net1001 _04656_ net850 vssd1 vssd1 vccd1 vccd1 _06049_ sky130_fd_sc_hd__and3_2
XTAP_TAPCELL_ROW_186_3233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11142_ net906 net1335 net862 _05076_ vssd1 vssd1 vccd1 vccd1 _01222_ sky130_fd_sc_hd__a31o_1
Xoutput43 net43 vssd1 vssd1 vccd1 vccd1 ADR_O[12] sky130_fd_sc_hd__buf_2
XANTENNA__07240__A2 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput54 net54 vssd1 vssd1 vccd1 vccd1 ADR_O[22] sky130_fd_sc_hd__buf_2
Xoutput65 net65 vssd1 vssd1 vccd1 vccd1 ADR_O[3] sky130_fd_sc_hd__buf_2
Xoutput76 net76 vssd1 vssd1 vccd1 vccd1 DAT_O[12] sky130_fd_sc_hd__clkbuf_4
Xoutput87 net87 vssd1 vssd1 vccd1 vccd1 DAT_O[22] sky130_fd_sc_hd__clkbuf_4
X_11073_ net89 net872 net836 net1130 vssd1 vssd1 vccd1 vccd1 _01184_ sky130_fd_sc_hd__a22o_1
Xoutput98 net98 vssd1 vssd1 vccd1 vccd1 DAT_O[3] sky130_fd_sc_hd__clkbuf_4
XANTENNA__07528__B1 net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08725__C1 _03740_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input30_A DAT_I[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10024_ net1846 net230 net619 vssd1 vssd1 vccd1 vccd1 _00227_ sky130_fd_sc_hd__mux2_1
XFILLER_0_208_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_187_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_201_3458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11975_ _05847_ _05849_ _05836_ vssd1 vssd1 vccd1 vccd1 _05858_ sky130_fd_sc_hd__a21boi_1
XANTENNA__09898__S net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13637__RESET_B net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13714_ clknet_leaf_96_clk _01285_ net984 vssd1 vssd1 vccd1 vccd1 top.a1.row2\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_10926_ net1746 net244 net593 vssd1 vssd1 vccd1 vccd1 _01087_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_197_3395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13645_ clknet_leaf_95_clk net1129 net983 vssd1 vssd1 vccd1 vccd1 top.ru.state\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10837__S net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10857_ net269 net2056 net596 vssd1 vssd1 vccd1 vccd1 _01018_ sky130_fd_sc_hd__mux2_1
XFILLER_0_171_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13576_ clknet_leaf_66_clk net1185 net1094 vssd1 vssd1 vccd1 vccd1 net98 sky130_fd_sc_hd__dfrtp_1
X_10788_ net1701 net156 net485 vssd1 vssd1 vccd1 vccd1 _00949_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_59_Right_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11241__B _01382_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06806__A2 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12527_ clknet_leaf_70_clk _00119_ vssd1 vssd1 vccd1 vccd1 top.a1.halfData\[5\] sky130_fd_sc_hd__dfxtp_2
X_12458_ clknet_leaf_65_clk _00053_ net1094 vssd1 vssd1 vccd1 vccd1 top.ramstore\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_152_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09756__A1 _04370_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11409_ _05288_ _05289_ _05290_ vssd1 vssd1 vccd1 vccd1 _05292_ sky130_fd_sc_hd__a21o_1
XANTENNA__10572__S net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12389_ clknet_leaf_94_clk top.ru.next_FetchedInstr\[1\] net981 vssd1 vssd1 vccd1
+ vccd1 top.a1.instruction\[1\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_93_1836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_1847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07767__B1 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07231__A2 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12519__RESET_B net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_185_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09508__A1 top.a1.instruction\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06950_ net808 net413 net438 vssd1 vssd1 vccd1 vccd1 _02089_ sky130_fd_sc_hd__o21a_1
XANTENNA__09084__D _04155_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_68_Right_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06881_ top.DUT.register\[23\]\[18\] net574 _02017_ _02019_ vssd1 vssd1 vccd1 vccd1
+ _02020_ sky130_fd_sc_hd__a211o_1
XFILLER_0_206_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08620_ _03742_ _03729_ _03741_ vssd1 vssd1 vccd1 vccd1 _03743_ sky130_fd_sc_hd__or3b_1
XANTENNA__11256__X _05149_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_2302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09381__B _01939_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_2313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_178_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_115 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08551_ net315 _03476_ vssd1 vssd1 vccd1 vccd1 _03677_ sky130_fd_sc_hd__and2_1
XFILLER_0_179_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07502_ top.DUT.register\[5\]\[14\] net652 net636 top.DUT.register\[6\]\[14\] _02639_
+ vssd1 vssd1 vccd1 vccd1 _02641_ sky130_fd_sc_hd__a221o_1
XANTENNA__07298__A2 net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08482_ net426 _03599_ _03610_ net428 _03609_ vssd1 vssd1 vccd1 vccd1 _03611_ sky130_fd_sc_hd__a221o_1
XFILLER_0_187_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_362 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11094__A3 net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07433_ top.DUT.register\[3\]\[15\] net552 net522 top.DUT.register\[10\]\[15\] vssd1
+ vssd1 vccd1 vccd1 _02572_ sky130_fd_sc_hd__a22o_1
XFILLER_0_134_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10747__S net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_77_Right_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout148_A _04938_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_170_3001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07364_ top.DUT.register\[4\]\[8\] net668 net731 top.DUT.register\[14\]\[8\] vssd1
+ vssd1 vccd1 vccd1 _02503_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_102_1976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09103_ _02341_ _04177_ _04149_ vssd1 vssd1 vccd1 vccd1 _04178_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_94_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06315_ _01331_ _01460_ vssd1 vssd1 vccd1 vccd1 _01469_ sky130_fd_sc_hd__and2_1
XFILLER_0_72_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07295_ _02432_ _02433_ vssd1 vssd1 vccd1 vccd1 _02434_ sky130_fd_sc_hd__nor2_2
XFILLER_0_150_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout315_A net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_374 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06245__B net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_652 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09034_ _01657_ _03179_ _03517_ vssd1 vssd1 vccd1 vccd1 _04109_ sky130_fd_sc_hd__or3_1
X_06246_ top.ramload\[7\] net852 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedData\[7\]
+ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_135_2464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_2475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09747__A1 _03663_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10482__S net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold320 top.DUT.register\[18\]\[19\] vssd1 vssd1 vccd1 vccd1 net1436 sky130_fd_sc_hd__dlygate4sd3_1
Xhold331 top.DUT.register\[25\]\[2\] vssd1 vssd1 vccd1 vccd1 net1447 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06177_ net904 _01409_ _01417_ vssd1 vssd1 vccd1 vccd1 _01419_ sky130_fd_sc_hd__or3_2
XFILLER_0_130_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold342 top.DUT.register\[20\]\[17\] vssd1 vssd1 vccd1 vccd1 net1458 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07758__B1 net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold353 top.DUT.register\[25\]\[23\] vssd1 vssd1 vccd1 vccd1 net1469 sky130_fd_sc_hd__dlygate4sd3_1
Xhold364 top.DUT.register\[2\]\[17\] vssd1 vssd1 vccd1 vccd1 net1480 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06261__A top.ramload\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold375 top.DUT.register\[24\]\[5\] vssd1 vssd1 vccd1 vccd1 net1491 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout800 net802 vssd1 vssd1 vccd1 vccd1 net800 sky130_fd_sc_hd__buf_2
Xhold386 top.DUT.register\[30\]\[14\] vssd1 vssd1 vccd1 vccd1 net1502 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_86_Right_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout811 net812 vssd1 vssd1 vccd1 vccd1 net811 sky130_fd_sc_hd__clkbuf_4
Xhold397 top.DUT.register\[26\]\[31\] vssd1 vssd1 vccd1 vccd1 net1513 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06430__B1 net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout822 _01578_ vssd1 vssd1 vccd1 vccd1 net822 sky130_fd_sc_hd__clkbuf_4
X_09936_ top.pc\[31\] _04644_ vssd1 vssd1 vccd1 vccd1 _04941_ sky130_fd_sc_hd__xnor2_1
Xfanout833 _01499_ vssd1 vssd1 vccd1 vccd1 net833 sky130_fd_sc_hd__buf_2
Xfanout844 _04666_ vssd1 vssd1 vccd1 vccd1 net844 sky130_fd_sc_hd__clkbuf_2
Xfanout855 _01433_ vssd1 vssd1 vccd1 vccd1 net855 sky130_fd_sc_hd__clkbuf_2
Xfanout866 _01427_ vssd1 vssd1 vccd1 vccd1 net866 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_181_3163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout877 _00012_ vssd1 vssd1 vccd1 vccd1 net877 sky130_fd_sc_hd__buf_4
X_09867_ net827 _04558_ _04877_ vssd1 vssd1 vccd1 vccd1 _04878_ sky130_fd_sc_hd__o21ba_1
XANTENNA_fanout472_X net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1020 top.ramload\[28\] vssd1 vssd1 vccd1 vccd1 net2136 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout888 top.a1.halfData\[0\] vssd1 vssd1 vccd1 vccd1 net888 sky130_fd_sc_hd__buf_2
Xhold1031 top.DUT.register\[5\]\[19\] vssd1 vssd1 vccd1 vccd1 net2147 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_175_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout899 net903 vssd1 vssd1 vccd1 vccd1 net899 sky130_fd_sc_hd__buf_4
XANTENNA__08722__A2 _03534_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_175_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1042 top.DUT.register\[26\]\[7\] vssd1 vssd1 vccd1 vccd1 net2158 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1053 top.DUT.register\[6\]\[2\] vssd1 vssd1 vccd1 vccd1 net2169 sky130_fd_sc_hd__dlygate4sd3_1
X_08818_ _03930_ _03931_ vssd1 vssd1 vccd1 vccd1 _03932_ sky130_fd_sc_hd__or2_1
XFILLER_0_197_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1064 top.DUT.register\[7\]\[20\] vssd1 vssd1 vccd1 vccd1 net2180 sky130_fd_sc_hd__dlygate4sd3_1
X_09798_ net829 _04446_ _04815_ vssd1 vssd1 vccd1 vccd1 _04816_ sky130_fd_sc_hd__o21ba_1
Xhold1075 top.DUT.register\[10\]\[18\] vssd1 vssd1 vccd1 vccd1 net2191 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1086 top.DUT.register\[21\]\[11\] vssd1 vssd1 vccd1 vccd1 net2202 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1097 top.pad.keyCode\[1\] vssd1 vssd1 vccd1 vccd1 net2213 sky130_fd_sc_hd__dlygate4sd3_1
X_08749_ _02221_ net431 net428 _03855_ _03862_ vssd1 vssd1 vccd1 vccd1 _03866_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout737_X net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_64_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11760_ _05638_ _05642_ vssd1 vssd1 vccd1 vccd1 _05643_ sky130_fd_sc_hd__and2b_1
XANTENNA__06497__B1 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_95_Right_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10711_ net1459 net190 net335 vssd1 vssd1 vccd1 vccd1 _00872_ sky130_fd_sc_hd__mux2_1
XANTENNA__10657__S net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout904_X net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11691_ _05546_ _05551_ vssd1 vssd1 vccd1 vccd1 _05574_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_48_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_193_652 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13430_ clknet_leaf_4_clk _01022_ net938 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[29\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_10642_ net209 net1540 net344 vssd1 vssd1 vccd1 vccd1 _00806_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_544 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_173 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08789__A2 net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13361_ clknet_leaf_112_clk _00953_ net990 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[27\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_10573_ top.DUT.register\[20\]\[10\] net228 net350 vssd1 vssd1 vccd1 vccd1 _00739_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07997__B1 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12312_ net2067 _06116_ net790 vssd1 vssd1 vccd1 vccd1 _06119_ sky130_fd_sc_hd__o21ai_1
X_13292_ clknet_4_15__leaf_clk _00884_ net1096 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[24\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_90_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07461__A2 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_251 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12243_ top.lcd.cnt_20ms\[12\] _06075_ net978 vssd1 vssd1 vccd1 vccd1 _06077_ sky130_fd_sc_hd__o21ai_1
XANTENNA__10392__S net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07749__B1 net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12174_ net1445 net848 net797 _05992_ vssd1 vssd1 vccd1 vccd1 _01282_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_75_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06171__A top.a1.halfData\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11125_ net54 net867 vssd1 vssd1 vccd1 vccd1 _05068_ sky130_fd_sc_hd__and2_1
XANTENNA__06421__B1 net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_166_2936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09482__A top.pc\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11056_ net102 net866 net837 net1207 vssd1 vssd1 vccd1 vccd1 _01167_ sky130_fd_sc_hd__a22o_1
XFILLER_0_204_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10007_ net159 net2183 net625 vssd1 vssd1 vccd1 vccd1 _00212_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_199_3424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_199_3435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_204_789 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09123__C1 _01505_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11958_ _05831_ net127 _05839_ _05828_ _05804_ vssd1 vssd1 vccd1 vccd1 _05841_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_80_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10909_ net1315 net194 net481 vssd1 vssd1 vccd1 vccd1 _01070_ sky130_fd_sc_hd__mux2_1
XANTENNA__10567__S net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_184_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11889_ _05725_ _05734_ _05752_ vssd1 vssd1 vccd1 vccd1 _05772_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_67_680 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13628_ clknet_leaf_75_clk _01215_ net1081 vssd1 vssd1 vccd1 vccd1 net55 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_184_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_183_195 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13559_ clknet_leaf_105_clk _01146_ net968 vssd1 vssd1 vccd1 vccd1 top.ramload\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_202_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07988__B1 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07080_ net823 _02218_ _01586_ vssd1 vssd1 vccd1 vccd1 _02219_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_89_68 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07452__A2 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09729__A1 _03569_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_2194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09944__X _04948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_479 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_130_2394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07982_ _03111_ _03120_ vssd1 vssd1 vccd1 vccd1 _03121_ sky130_fd_sc_hd__or2_4
XFILLER_0_10_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06933_ top.DUT.register\[21\]\[21\] net657 net721 top.DUT.register\[19\]\[21\] _02071_
+ vssd1 vssd1 vccd1 vccd1 _02072_ sky130_fd_sc_hd__a221o_1
X_09721_ net2082 net247 net631 vssd1 vssd1 vccd1 vccd1 _00128_ sky130_fd_sc_hd__mux2_1
X_06864_ net808 net414 net438 vssd1 vssd1 vccd1 vccd1 _02003_ sky130_fd_sc_hd__o21a_1
X_09652_ top.edg2.button_i _04688_ _04692_ vssd1 vssd1 vccd1 vccd1 _04693_ sky130_fd_sc_hd__or3_1
X_08603_ _02613_ _02654_ vssd1 vssd1 vccd1 vccd1 _03726_ sky130_fd_sc_hd__or2_1
XFILLER_0_96_208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09583_ _01572_ _04628_ vssd1 vssd1 vccd1 vccd1 _04630_ sky130_fd_sc_hd__nor2_1
X_06795_ top.DUT.register\[20\]\[17\] net563 net444 top.DUT.register\[1\]\[17\] _01933_
+ vssd1 vssd1 vccd1 vccd1 _01934_ sky130_fd_sc_hd__a221o_1
XFILLER_0_179_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout265_A _04729_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08534_ _03659_ _03660_ vssd1 vssd1 vccd1 vccd1 _03661_ sky130_fd_sc_hd__or2_1
XFILLER_0_210_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08736__A net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13141__RESET_B net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_490 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08465_ net886 top.pc\[9\] net697 _03594_ vssd1 vssd1 vccd1 vccd1 _03595_ sky130_fd_sc_hd__a22o_1
XFILLER_0_37_319 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10477__S net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout432_A net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07416_ top.DUT.register\[24\]\[9\] net643 net722 top.DUT.register\[29\]\[9\] vssd1
+ vssd1 vccd1 vccd1 _02555_ sky130_fd_sc_hd__a22o_1
XFILLER_0_18_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_137_2504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08396_ net315 _03527_ vssd1 vssd1 vccd1 vccd1 _03528_ sky130_fd_sc_hd__or2_1
XANTENNA__07691__A2 _02808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07347_ top.DUT.register\[29\]\[8\] net452 net508 top.DUT.register\[4\]\[8\] _02485_
+ vssd1 vssd1 vccd1 vccd1 _02486_ sky130_fd_sc_hd__a221o_1
XFILLER_0_45_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07979__B1 net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout318_X net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07639__X _02778_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07443__A2 net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07278_ top.DUT.register\[23\]\[13\] net674 net713 top.DUT.register\[11\]\[13\] vssd1
+ vssd1 vccd1 vccd1 _02417_ sky130_fd_sc_hd__a22o_1
XFILLER_0_131_711 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09017_ _03865_ _03966_ _04091_ _03708_ vssd1 vssd1 vccd1 vccd1 _04092_ sky130_fd_sc_hd__or4b_1
XANTENNA_fanout899_A net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06229_ top.ramload\[23\] net858 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedInstr\[23\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_60_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07358__Y _02497_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08928__C1 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold150 _01353_ vssd1 vssd1 vccd1 vccd1 net1266 sky130_fd_sc_hd__dlygate4sd3_1
Xhold161 top.DUT.register\[15\]\[30\] vssd1 vssd1 vccd1 vccd1 net1277 sky130_fd_sc_hd__dlygate4sd3_1
Xhold172 top.a1.row2\[24\] vssd1 vssd1 vccd1 vccd1 net1288 sky130_fd_sc_hd__dlygate4sd3_1
Xhold183 top.a1.row2\[8\] vssd1 vssd1 vccd1 vccd1 net1299 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold194 top.DUT.register\[15\]\[18\] vssd1 vssd1 vccd1 vccd1 net1310 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10940__S net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout630 _04948_ vssd1 vssd1 vccd1 vccd1 net630 sky130_fd_sc_hd__buf_4
Xfanout641 _01619_ vssd1 vssd1 vccd1 vccd1 net641 sky130_fd_sc_hd__clkbuf_8
Xfanout652 _01610_ vssd1 vssd1 vccd1 vccd1 net652 sky130_fd_sc_hd__clkbuf_4
X_09919_ net828 _04613_ vssd1 vssd1 vccd1 vccd1 _04926_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_148_2666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout663 _01605_ vssd1 vssd1 vccd1 vccd1 net663 sky130_fd_sc_hd__buf_6
XANTENNA_fanout854_X net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout674 _01597_ vssd1 vssd1 vccd1 vccd1 net674 sky130_fd_sc_hd__buf_4
Xfanout685 _01510_ vssd1 vssd1 vccd1 vccd1 net685 sky130_fd_sc_hd__buf_1
XANTENNA_clkbuf_3_1_0_clk_X clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout696 net697 vssd1 vssd1 vccd1 vccd1 net696 sky130_fd_sc_hd__buf_2
X_12930_ clknet_leaf_25_clk _00522_ net1012 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[13\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_198_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_161_2855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_161_2866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12861_ clknet_leaf_119_clk _00453_ net930 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[11\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_201_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_198_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_201_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11812_ _05693_ _05694_ vssd1 vssd1 vccd1 vccd1 _05695_ sky130_fd_sc_hd__or2_1
XFILLER_0_139_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12792_ clknet_leaf_125_clk _00384_ net924 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[9\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_68_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10266__A1 net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_194_3354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11743_ _01399_ _05585_ _05620_ vssd1 vssd1 vccd1 vccd1 _05626_ sky130_fd_sc_hd__and3_1
XANTENNA__10387__S net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07682__A2 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11674_ top.a1.dataIn\[10\] _05550_ _05554_ _05555_ vssd1 vssd1 vccd1 vccd1 _05557_
+ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__06166__A net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_12_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13413_ clknet_leaf_35_clk _01005_ net1041 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[28\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_10625_ net152 top.DUT.register\[21\]\[29\] net349 vssd1 vssd1 vccd1 vccd1 _00790_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__06890__B1 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_77_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10556_ net1991 net164 net355 vssd1 vssd1 vccd1 vccd1 _00723_ sky130_fd_sc_hd__mux2_1
XANTENNA__08631__A1 net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07434__A2 net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13344_ clknet_leaf_55_clk _00936_ net1072 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[26\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_134_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10487_ net1257 net175 net363 vssd1 vssd1 vccd1 vccd1 _00657_ sky130_fd_sc_hd__mux2_1
X_13275_ clknet_leaf_126_clk _00867_ net924 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[24\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_12226_ net1190 _06052_ _06066_ net978 vssd1 vssd1 vccd1 vccd1 _01316_ sky130_fd_sc_hd__o211a_1
XFILLER_0_122_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_184_Right_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12404__Q top.a1.instruction\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10850__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12157_ _06038_ _06039_ vssd1 vssd1 vccd1 vccd1 _06040_ sky130_fd_sc_hd__or2_1
XFILLER_0_75_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11108_ net906 net1286 net861 _05059_ vssd1 vssd1 vccd1 vccd1 _01205_ sky130_fd_sc_hd__a31o_1
X_12088_ top.a1.dataIn\[3\] _05948_ vssd1 vssd1 vccd1 vccd1 _05971_ sky130_fd_sc_hd__nor2_1
X_11039_ net19 net838 net816 net2051 vssd1 vssd1 vccd1 vccd1 _01151_ sky130_fd_sc_hd__o22a_1
XFILLER_0_204_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_88_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06580_ top.DUT.register\[30\]\[28\] net582 net450 top.DUT.register\[21\]\[28\] _01718_
+ vssd1 vssd1 vccd1 vccd1 _01719_ sky130_fd_sc_hd__a221o_1
XFILLER_0_87_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_188_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10297__S net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07122__A1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08275__B _02899_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08250_ net315 _03381_ vssd1 vssd1 vccd1 vccd1 _03387_ sky130_fd_sc_hd__nor2_1
XFILLER_0_28_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_31_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09939__X _04944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07673__A2 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07201_ net795 _02331_ _02335_ _02339_ vssd1 vssd1 vccd1 vccd1 _02340_ sky130_fd_sc_hd__nor4_1
XTAP_TAPCELL_ROW_119_2234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08181_ _03317_ _03318_ vssd1 vssd1 vccd1 vccd1 _03319_ sky130_fd_sc_hd__nand2_1
XFILLER_0_131_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07132_ top.DUT.register\[2\]\[11\] net559 net527 top.DUT.register\[26\]\[11\] _02270_
+ vssd1 vssd1 vccd1 vccd1 _02271_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_41_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07425__A2 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_132_2423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06633__B1 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07063_ top.DUT.register\[7\]\[22\] net662 net769 top.DUT.register\[28\]\[22\] _02200_
+ vssd1 vssd1 vccd1 vccd1 _02202_ sky130_fd_sc_hd__a221o_1
XFILLER_0_11_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_151_Right_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10760__S net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07965_ top.DUT.register\[28\]\[31\] net556 net510 top.DUT.register\[4\]\[31\] _03103_
+ vssd1 vssd1 vccd1 vccd1 _03104_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout382_A net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13035__CLK clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09704_ _04716_ _04735_ vssd1 vssd1 vccd1 vccd1 _04736_ sky130_fd_sc_hd__or2_1
X_06916_ top.DUT.register\[2\]\[21\] net562 net454 top.DUT.register\[29\]\[21\] vssd1
+ vssd1 vccd1 vccd1 _02055_ sky130_fd_sc_hd__a22o_1
XFILLER_0_156_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07896_ top.DUT.register\[20\]\[1\] net566 net538 top.DUT.register\[19\]\[1\] vssd1
+ vssd1 vccd1 vccd1 _03035_ sky130_fd_sc_hd__a22o_1
XANTENNA__09850__A top.pc\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09635_ top.pad.keyCode\[4\] top.pad.keyCode\[5\] top.pad.keyCode\[7\] top.pad.keyCode\[6\]
+ vssd1 vssd1 vccd1 vccd1 _04677_ sky130_fd_sc_hd__or4b_2
XANTENNA_clkbuf_leaf_4_clk_A clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06847_ top.DUT.register\[9\]\[19\] net764 net753 top.DUT.register\[26\]\[19\] vssd1
+ vssd1 vccd1 vccd1 _01986_ sky130_fd_sc_hd__a22o_1
XANTENNA__08737__Y _03854_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout647_A _01612_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_143_2585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_2596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06778_ net808 _01916_ net438 vssd1 vssd1 vccd1 vccd1 _01917_ sky130_fd_sc_hd__o21a_1
X_09566_ top.pc\[29\] _04605_ vssd1 vssd1 vccd1 vccd1 _04614_ sky130_fd_sc_hd__and2_1
XANTENNA__13185__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08517_ net297 _03440_ vssd1 vssd1 vccd1 vccd1 _03644_ sky130_fd_sc_hd__nand2_1
XFILLER_0_77_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09231__A_N _02502_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout814_A _01446_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09497_ _01505_ _04548_ _04549_ _04205_ vssd1 vssd1 vccd1 vccd1 _04550_ sky130_fd_sc_hd__a31o_1
XANTENNA__09996__S net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_176_3084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10000__S net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08448_ _03577_ vssd1 vssd1 vccd1 vccd1 _03578_ sky130_fd_sc_hd__inv_2
XANTENNA__11323__C top.a1.dataIn\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06872__B1 net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08379_ net430 _03508_ _03510_ _03334_ _03511_ vssd1 vssd1 vccd1 vccd1 _03512_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout602_X net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10935__S net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_288 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08913__B _03099_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_631 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10410_ net1314 net208 net370 vssd1 vssd1 vccd1 vccd1 _00582_ sky130_fd_sc_hd__mux2_1
X_11390_ _05234_ _05262_ vssd1 vssd1 vccd1 vccd1 _05273_ sky130_fd_sc_hd__xor2_2
XANTENNA__07416__A2 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_190_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_59_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10341_ net1928 net211 net377 vssd1 vssd1 vccd1 vccd1 _00517_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_59_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_563 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13060_ clknet_leaf_37_clk _00652_ net1051 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[17\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_10272_ net1456 net233 net385 vssd1 vssd1 vccd1 vccd1 _00450_ sky130_fd_sc_hd__mux2_1
X_12011_ _05883_ _05885_ _05861_ vssd1 vssd1 vccd1 vccd1 _05894_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_72_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08916__A2 _04020_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10670__S net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08129__B1 _03265_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout460 _01552_ vssd1 vssd1 vccd1 vccd1 net460 sky130_fd_sc_hd__buf_4
Xfanout471 net472 vssd1 vssd1 vccd1 vccd1 net471 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_205_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout482 _04962_ vssd1 vssd1 vccd1 vccd1 net482 sky130_fd_sc_hd__clkbuf_8
Xfanout493 _03339_ vssd1 vssd1 vccd1 vccd1 net493 sky130_fd_sc_hd__clkbuf_2
X_12913_ clknet_leaf_111_clk _00505_ net988 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[13\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_201_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_186_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_17_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12844_ clknet_leaf_63_clk _00436_ net1093 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[10\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_158_427 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_139_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12775_ clknet_leaf_6_clk _00367_ net944 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[8\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08301__B1 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_83_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11726_ _05605_ _05607_ vssd1 vssd1 vccd1 vccd1 _05609_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_83_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07655__A2 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11233__C _05123_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08852__B2 _03264_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10845__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_181_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11657_ _05492_ _05538_ vssd1 vssd1 vccd1 vccd1 _05540_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_4_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_211_3608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_211_3619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10608_ net214 net2041 net346 vssd1 vssd1 vccd1 vccd1 _00773_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_344 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_181_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11588_ _05432_ net250 vssd1 vssd1 vccd1 vccd1 _05471_ sky130_fd_sc_hd__nand2_1
X_13327_ clknet_leaf_32_clk _00919_ net1045 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[25\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold908 top.DUT.register\[11\]\[11\] vssd1 vssd1 vccd1 vccd1 net2024 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10539_ net1641 _04760_ net354 vssd1 vssd1 vccd1 vccd1 _00706_ sky130_fd_sc_hd__mux2_1
Xhold919 top.DUT.register\[6\]\[1\] vssd1 vssd1 vccd1 vccd1 net2035 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_114_2153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13258_ clknet_leaf_118_clk _00850_ net954 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[23\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08368__B1 _03495_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12209_ top.lcd.cnt_20ms\[9\] top.lcd.cnt_20ms\[7\] top.lcd.cnt_20ms\[6\] top.lcd.cnt_20ms\[8\]
+ vssd1 vssd1 vccd1 vccd1 _06055_ sky130_fd_sc_hd__or4b_1
XANTENNA__10580__S net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13189_ clknet_leaf_35_clk _00781_ net1041 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[21\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_209_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_208_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09580__A2 _04620_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07750_ _02882_ _02884_ _02886_ _02888_ vssd1 vssd1 vccd1 vccd1 _02889_ sky130_fd_sc_hd__or4_4
XFILLER_0_193_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09332__A2 top.pc\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06701_ top.DUT.register\[16\]\[25\] net543 net439 top.DUT.register\[5\]\[25\] _01839_
+ vssd1 vssd1 vccd1 vccd1 _01840_ sky130_fd_sc_hd__a221o_1
X_07681_ top.DUT.register\[5\]\[4\] net653 net756 top.DUT.register\[1\]\[4\] _02819_
+ vssd1 vssd1 vccd1 vccd1 _02820_ sky130_fd_sc_hd__a221o_1
XFILLER_0_211_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06632_ top.DUT.register\[4\]\[27\] net670 net666 top.DUT.register\[20\]\[27\] _01770_
+ vssd1 vssd1 vccd1 vccd1 _01771_ sky130_fd_sc_hd__a221o_1
X_09420_ net901 top.pc\[19\] _04477_ net891 vssd1 vssd1 vccd1 vccd1 _00099_ sky130_fd_sc_hd__o211a_1
XFILLER_0_149_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07902__B _03040_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07894__A2 net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06563_ _01701_ vssd1 vssd1 vccd1 vccd1 _01702_ sky130_fd_sc_hd__inv_2
X_09351_ _04410_ _04411_ vssd1 vssd1 vccd1 vccd1 _04412_ sky130_fd_sc_hd__or2_1
X_08302_ _03436_ vssd1 vssd1 vccd1 vccd1 _03437_ sky130_fd_sc_hd__inv_2
XFILLER_0_74_222 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09282_ top.pc\[12\] _04336_ vssd1 vssd1 vccd1 vccd1 _04347_ sky130_fd_sc_hd__and2_1
X_06494_ top.DUT.register\[8\]\[30\] net641 net756 top.DUT.register\[1\]\[30\] _01632_
+ vssd1 vssd1 vccd1 vccd1 _01633_ sky130_fd_sc_hd__a221o_1
XANTENNA__07646__A2 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08233_ _03368_ _03369_ net302 vssd1 vssd1 vccd1 vccd1 _03370_ sky130_fd_sc_hd__mux2_2
XFILLER_0_28_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06854__B1 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_195 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_96 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10755__S net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09829__B _04499_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout228_A net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08164_ _03300_ _03301_ vssd1 vssd1 vccd1 vccd1 _03302_ sky130_fd_sc_hd__nand2_1
XFILLER_0_160_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_815 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07115_ top.DUT.register\[1\]\[16\] net755 net719 top.DUT.register\[19\]\[16\] vssd1
+ vssd1 vccd1 vccd1 _02254_ sky130_fd_sc_hd__a22o_1
X_08095_ _02773_ net330 vssd1 vssd1 vccd1 vccd1 _03234_ sky130_fd_sc_hd__nand2_1
XANTENNA__06253__B net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload70 clknet_leaf_52_clk vssd1 vssd1 vccd1 vccd1 clkload70/Y sky130_fd_sc_hd__clkinv_4
X_07046_ top.DUT.register\[9\]\[22\] net470 net523 top.DUT.register\[11\]\[22\] _02184_
+ vssd1 vssd1 vccd1 vccd1 _02185_ sky130_fd_sc_hd__a221o_1
Xclkload81 clknet_leaf_43_clk vssd1 vssd1 vccd1 vccd1 clkload81/Y sky130_fd_sc_hd__inv_6
Xclkload92 clknet_leaf_79_clk vssd1 vssd1 vccd1 vccd1 clkload92/Y sky130_fd_sc_hd__clkinv_4
XANTENNA_fanout597_A _04966_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10490__S net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06540__Y _01679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07031__B1 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08997_ _03556_ _03580_ _03606_ _03632_ vssd1 vssd1 vccd1 vccd1 _04072_ sky130_fd_sc_hd__and4_1
XANTENNA_fanout764_A net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout385_X net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_2614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_2625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07948_ _02223_ _03081_ _02111_ _02132_ vssd1 vssd1 vccd1 vccd1 _03087_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA_fanout931_A net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout552_X net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07879_ _03013_ _03015_ _03017_ vssd1 vssd1 vccd1 vccd1 _03018_ sky130_fd_sc_hd__or3_1
XANTENNA__07334__A1 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_178_3113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09618_ top.a1.state\[1\] top.a1.state\[0\] top.a1.state\[2\] vssd1 vssd1 vccd1 vccd1
+ _04663_ sky130_fd_sc_hd__or3b_1
X_10890_ net1829 net264 net478 vssd1 vssd1 vccd1 vccd1 _01051_ sky130_fd_sc_hd__mux2_1
XANTENNA__07885__A2 net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09549_ top.pc\[27\] _04567_ top.pc\[28\] vssd1 vssd1 vccd1 vccd1 _04598_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_109_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_191_3313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07098__B1 net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_195_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_176_780 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12560_ clknet_leaf_29_clk _00152_ net1017 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[1\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_108_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06845__B1 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11511_ _05353_ _05381_ vssd1 vssd1 vccd1 vccd1 _05394_ sky130_fd_sc_hd__xor2_1
XFILLER_0_53_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10665__S net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_199_Left_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12491_ clknet_leaf_87_clk _00083_ net1006 vssd1 vssd1 vccd1 vccd1 top.pc\[3\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__08643__B _03760_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06715__Y _01854_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_163_463 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_156_2787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11442_ _05287_ net278 vssd1 vssd1 vccd1 vccd1 _05325_ sky130_fd_sc_hd__nand2_1
XFILLER_0_135_198 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11373_ _05220_ _05252_ vssd1 vssd1 vccd1 vccd1 _05256_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_189_3275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10324_ net156 net1772 net383 vssd1 vssd1 vccd1 vccd1 _00501_ sky130_fd_sc_hd__mux2_1
X_13112_ clknet_leaf_128_clk _00704_ net912 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[19\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_189_3286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09547__C1 net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13043_ clknet_leaf_120_clk _00635_ net932 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[17\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_10255_ net168 net1853 net389 vssd1 vssd1 vccd1 vccd1 _00434_ sky130_fd_sc_hd__mux2_1
XANTENNA__07022__B1 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13350__CLK clknet_leaf_40_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10186_ _04154_ net689 _04713_ vssd1 vssd1 vccd1 vccd1 _04966_ sky130_fd_sc_hd__or3b_4
XANTENNA__06376__A2 net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_208_3570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout290 net294 vssd1 vssd1 vccd1 vccd1 net290 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__07562__X _02701_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_202_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_85_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkload6_A clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07876__A2 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_186_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12827_ clknet_leaf_120_clk _00419_ net929 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[10\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07089__B1 net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07628__A2 net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12758_ clknet_leaf_12_clk _00350_ net942 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[8\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_139_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11709_ _05565_ _05591_ vssd1 vssd1 vccd1 vccd1 _05592_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10575__S net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12689_ clknet_leaf_111_clk _00281_ net988 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[6\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06625__Y _01764_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_614 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_642 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_141_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08589__B1 _03711_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold705 top.DUT.register\[20\]\[9\] vssd1 vssd1 vccd1 vccd1 net1821 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_203_Left_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09087__D _01607_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold716 top.DUT.register\[28\]\[30\] vssd1 vssd1 vccd1 vccd1 net1832 sky130_fd_sc_hd__dlygate4sd3_1
Xhold727 top.DUT.register\[23\]\[5\] vssd1 vssd1 vccd1 vccd1 net1843 sky130_fd_sc_hd__dlygate4sd3_1
Xhold738 top.DUT.register\[3\]\[9\] vssd1 vssd1 vccd1 vccd1 net1854 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_96_1889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07261__B1 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold749 top.DUT.register\[20\]\[8\] vssd1 vssd1 vccd1 vccd1 net1865 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07800__A2 net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08920_ _04009_ _04027_ vssd1 vssd1 vccd1 vccd1 _04029_ sky130_fd_sc_hd__or2_1
XANTENNA__06801__B _01939_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07013__B1 net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08851_ net281 _03408_ _03886_ vssd1 vssd1 vccd1 vccd1 _03963_ sky130_fd_sc_hd__o21a_1
XANTENNA__07564__A1 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07802_ top.DUT.register\[8\]\[2\] net539 net531 top.DUT.register\[12\]\[2\] vssd1
+ vssd1 vccd1 vccd1 _02941_ sky130_fd_sc_hd__a22o_1
X_08782_ net497 _03896_ vssd1 vssd1 vccd1 vccd1 _03897_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_127_2344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_127_2355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07733_ top.DUT.register\[23\]\[3\] net674 net744 top.DUT.register\[2\]\[3\] _02871_
+ vssd1 vssd1 vccd1 vccd1 _02872_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_0_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07867__A2 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07664_ _02800_ _02802_ vssd1 vssd1 vccd1 vccd1 _02803_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_140_2544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09403_ top.pc\[18\] top.pc\[19\] _04428_ vssd1 vssd1 vccd1 vccd1 _04461_ sky130_fd_sc_hd__and3_1
X_06615_ _01747_ _01749_ _01751_ _01753_ vssd1 vssd1 vccd1 vccd1 _01754_ sky130_fd_sc_hd__or4_4
XANTENNA__11154__B _05082_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07595_ top.DUT.register\[7\]\[6\] net659 net754 top.DUT.register\[1\]\[6\] _02733_
+ vssd1 vssd1 vccd1 vccd1 _02734_ sky130_fd_sc_hd__a221o_1
XFILLER_0_48_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout345_A _04992_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06248__B net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_84 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1087_A net1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06546_ top.DUT.register\[7\]\[29\] net661 net748 top.DUT.register\[17\]\[29\] _01684_
+ vssd1 vssd1 vccd1 vccd1 _01685_ sky130_fd_sc_hd__a221o_1
X_09334_ top.pc\[15\] _04386_ vssd1 vssd1 vccd1 vccd1 _04396_ sky130_fd_sc_hd__and2_1
XFILLER_0_192_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07619__A2 net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_192_547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_173_3043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06827__B1 net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06477_ net787 _01600_ _01602_ vssd1 vssd1 vccd1 vccd1 _01616_ sky130_fd_sc_hd__and3_1
X_09265_ _04329_ _04330_ vssd1 vssd1 vccd1 vccd1 _04331_ sky130_fd_sc_hd__nor2_1
XANTENNA__10485__S net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08292__A2 _03427_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout133_X net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout512_A _01559_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08216_ net884 top.pc\[1\] net695 _03353_ vssd1 vssd1 vccd1 vccd1 _03354_ sky130_fd_sc_hd__a22o_1
X_09196_ _01505_ _04265_ _04266_ _04260_ _01393_ vssd1 vssd1 vccd1 vccd1 _04267_ sky130_fd_sc_hd__a311o_1
XANTENNA__06264__A top.ramload\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08147_ _02899_ net300 vssd1 vssd1 vccd1 vccd1 _03285_ sky130_fd_sc_hd__nand2_1
XANTENNA__09241__A1 net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07252__B1 net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08078_ net291 _03216_ vssd1 vssd1 vccd1 vccd1 _03217_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout881_A net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_178_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07029_ top.DUT.register\[25\]\[20\] net781 net729 top.DUT.register\[18\]\[20\] _02165_
+ vssd1 vssd1 vccd1 vccd1 _02168_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout979_A net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07807__B _02944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07004__B1 net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10040_ net2270 net164 net621 vssd1 vssd1 vccd1 vccd1 _00243_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09862__X _04874_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold10 top.a1.dataInTemp\[2\] vssd1 vssd1 vccd1 vccd1 net1126 sky130_fd_sc_hd__dlygate4sd3_1
Xhold21 _01190_ vssd1 vssd1 vccd1 vccd1 net1137 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout767_X net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold32 _01189_ vssd1 vssd1 vccd1 vccd1 net1148 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12502__Q top.pc\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold43 top.a1.data\[1\] vssd1 vssd1 vccd1 vccd1 net1159 sky130_fd_sc_hd__dlygate4sd3_1
Xhold54 net114 vssd1 vssd1 vccd1 vccd1 net1170 sky130_fd_sc_hd__dlygate4sd3_1
Xhold65 _01171_ vssd1 vssd1 vccd1 vccd1 net1181 sky130_fd_sc_hd__dlygate4sd3_1
Xhold76 top.a1.row1\[105\] vssd1 vssd1 vccd1 vccd1 net1192 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold87 _01172_ vssd1 vssd1 vccd1 vccd1 net1203 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11991_ _05845_ _05855_ vssd1 vssd1 vccd1 vccd1 _05874_ sky130_fd_sc_hd__xnor2_1
Xhold98 net100 vssd1 vssd1 vccd1 vccd1 net1214 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_202_128 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13730_ clknet_leaf_96_clk _01301_ vssd1 vssd1 vccd1 vccd1 top.a1.dataInTemp\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_10942_ net1331 net181 net593 vssd1 vssd1 vccd1 vccd1 _01103_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_67_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_27_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13661_ clknet_leaf_91_clk _01237_ net995 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[107\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_211_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10873_ net216 net1878 net595 vssd1 vssd1 vccd1 vccd1 _01034_ sky130_fd_sc_hd__mux2_1
XANTENNA__06530__A2 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_183_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_158_2816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12612_ clknet_leaf_36_clk _00204_ net1049 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[3\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_155_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13592_ clknet_leaf_63_clk net1155 net1066 vssd1 vssd1 vccd1 vccd1 net83 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_155_227 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06818__B1 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_372 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12543_ clknet_leaf_24_clk _00135_ net1015 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[1\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_136_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09480__A1 net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08373__B _03505_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_567 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07491__B1 net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12474_ clknet_leaf_47_clk _00069_ net1067 vssd1 vssd1 vccd1 vccd1 top.ramstore\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_124_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_163_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_91_clk_A clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11425_ _05273_ _05307_ vssd1 vssd1 vccd1 vccd1 _05308_ sky130_fd_sc_hd__or2_1
XFILLER_0_22_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_7 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13425__RESET_B net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07243__B1 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09485__A top.pc\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11356_ _05207_ _05214_ _05218_ top.a1.dataIn\[27\] top.a1.dataIn\[26\] vssd1 vssd1
+ vccd1 vccd1 _05239_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_111_2112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12119__A1 top.a1.dataIn\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06597__A2 net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10307_ net219 net2227 net381 vssd1 vssd1 vccd1 vccd1 _00484_ sky130_fd_sc_hd__mux2_1
X_11287_ top.a1.row1\[11\] _05126_ _05171_ _05175_ _05176_ vssd1 vssd1 vccd1 vccd1
+ _05177_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_169_2978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13026_ clknet_leaf_10_clk _00618_ net949 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[16\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_10238_ net237 net1876 net392 vssd1 vssd1 vccd1 vccd1 _00417_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_206_3529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1030 net1032 vssd1 vssd1 vccd1 vccd1 net1030 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12412__Q top.a1.instruction\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1041 net1042 vssd1 vssd1 vccd1 vccd1 net1041 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09940__C1 _04944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1052 net1071 vssd1 vssd1 vccd1 vccd1 net1052 sky130_fd_sc_hd__buf_2
X_10169_ net1794 net176 net603 vssd1 vssd1 vccd1 vccd1 _00368_ sky130_fd_sc_hd__mux2_1
Xfanout1063 net1070 vssd1 vssd1 vccd1 vccd1 net1063 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_83_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1074 net1087 vssd1 vssd1 vccd1 vccd1 net1074 sky130_fd_sc_hd__clkbuf_4
Xfanout1085 net1086 vssd1 vssd1 vccd1 vccd1 net1085 sky130_fd_sc_hd__clkbuf_2
Xfanout1096 net1097 vssd1 vssd1 vccd1 vccd1 net1096 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_109_2074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_2085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_656 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07849__A2 net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_190_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_44_clk_A clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_199 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_122_2274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06521__A2 net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06400_ net685 _01527_ _01531_ vssd1 vssd1 vccd1 vccd1 _01539_ sky130_fd_sc_hd__and3_1
XFILLER_0_57_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07380_ top.DUT.register\[24\]\[8\] net644 net703 top.DUT.register\[3\]\[8\] _02518_
+ vssd1 vssd1 vccd1 vccd1 _02519_ sky130_fd_sc_hd__a221o_1
XFILLER_0_174_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_174_558 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06331_ top.a1.instruction\[13\] top.a1.instruction\[14\] vssd1 vssd1 vccd1 vccd1
+ _01478_ sky130_fd_sc_hd__or2_1
XFILLER_0_72_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06809__B1 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_1918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09050_ net321 _03530_ _03845_ _03855_ _04124_ vssd1 vssd1 vccd1 vccd1 _04125_ sky130_fd_sc_hd__a2111o_1
X_06262_ top.ramload\[23\] net853 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedData\[23\]
+ sky130_fd_sc_hd__and2_1
XANTENNA__07482__B1 net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08001_ _03135_ _03137_ _03139_ vssd1 vssd1 vccd1 vccd1 _03140_ sky130_fd_sc_hd__or3_1
XFILLER_0_115_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06193_ net1118 net887 net886 vssd1 vssd1 vccd1 vccd1 _00010_ sky130_fd_sc_hd__a21o_1
XANTENNA__08026__A2 _03142_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_102_clk_A clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold502 top.DUT.register\[21\]\[15\] vssd1 vssd1 vccd1 vccd1 net1618 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold513 top.ramaddr\[15\] vssd1 vssd1 vccd1 vccd1 net1629 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07234__B1 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold524 top.DUT.register\[14\]\[7\] vssd1 vssd1 vccd1 vccd1 net1640 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08503__S net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold535 top.DUT.register\[28\]\[7\] vssd1 vssd1 vccd1 vccd1 net1651 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06588__A2 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold546 top.DUT.register\[22\]\[2\] vssd1 vssd1 vccd1 vccd1 net1662 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_464 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07785__A1 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold557 top.DUT.register\[4\]\[17\] vssd1 vssd1 vccd1 vccd1 net1673 sky130_fd_sc_hd__dlygate4sd3_1
Xhold568 top.ramload\[13\] vssd1 vssd1 vccd1 vccd1 net1684 sky130_fd_sc_hd__dlygate4sd3_1
X_09952_ net1463 net247 net627 vssd1 vssd1 vccd1 vccd1 _00160_ sky130_fd_sc_hd__mux2_1
Xhold579 top.DUT.register\[10\]\[3\] vssd1 vssd1 vccd1 vccd1 net1695 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08903_ net1760 net831 net801 _04012_ vssd1 vssd1 vccd1 vccd1 _00047_ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_117_clk_A clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09883_ net827 _04569_ _04892_ vssd1 vssd1 vccd1 vccd1 _04893_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_5_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08834_ _01834_ _03092_ vssd1 vssd1 vccd1 vccd1 _03947_ sky130_fd_sc_hd__and2_1
XANTENNA__09931__C1 _04936_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10988__B net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08765_ net281 _03527_ vssd1 vssd1 vccd1 vccd1 _03881_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout462_A _01552_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06760__A2 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07716_ net820 net410 _02854_ net805 vssd1 vssd1 vccd1 vccd1 _02855_ sky130_fd_sc_hd__a31o_1
X_08696_ _02179_ _03813_ vssd1 vssd1 vccd1 vccd1 _03815_ sky130_fd_sc_hd__nor2_1
XANTENNA__06259__A top.ramload\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07647_ top.DUT.register\[23\]\[5\] net671 net639 top.DUT.register\[8\]\[5\] _02784_
+ vssd1 vssd1 vccd1 vccd1 _02786_ sky130_fd_sc_hd__a221o_1
XFILLER_0_94_114 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_339 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout727_A _01628_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout348_X net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06512__A2 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_177_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07578_ top.DUT.register\[8\]\[6\] net539 net443 top.DUT.register\[1\]\[6\] _02716_
+ vssd1 vssd1 vccd1 vccd1 _02717_ sky130_fd_sc_hd__a221o_1
XFILLER_0_82_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06169__A_N top.a1.halfData\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_165_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09317_ _04365_ _04366_ _04363_ vssd1 vssd1 vccd1 vccd1 _04380_ sky130_fd_sc_hd__o21bai_1
X_06529_ _01661_ _01663_ _01665_ _01667_ vssd1 vssd1 vccd1 vccd1 _01668_ sky130_fd_sc_hd__or4_1
XANTENNA__09289__B _02453_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout515_X net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_539 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09248_ _04314_ vssd1 vssd1 vccd1 vccd1 _04315_ sky130_fd_sc_hd__inv_2
XFILLER_0_106_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_173_591 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_153_2735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_153_2746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12763__CLK clknet_leaf_120_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09179_ net136 _04238_ _04250_ net899 vssd1 vssd1 vccd1 vccd1 _04251_ sky130_fd_sc_hd__o211ai_1
XANTENNA__10943__S net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11210_ _05111_ net1234 net471 vssd1 vssd1 vccd1 vccd1 _01255_ sky130_fd_sc_hd__mux2_1
X_12190_ net1283 net848 _05082_ vssd1 vssd1 vccd1 vccd1 _01298_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_186_3234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06579__A2 net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11141_ net63 net867 vssd1 vssd1 vccd1 vccd1 _05076_ sky130_fd_sc_hd__and2_1
Xoutput44 net44 vssd1 vssd1 vccd1 vccd1 ADR_O[13] sky130_fd_sc_hd__buf_2
Xoutput55 net55 vssd1 vssd1 vccd1 vccd1 ADR_O[23] sky130_fd_sc_hd__buf_2
XFILLER_0_9_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput66 net66 vssd1 vssd1 vccd1 vccd1 ADR_O[4] sky130_fd_sc_hd__buf_2
Xoutput77 net77 vssd1 vssd1 vccd1 vccd1 DAT_O[13] sky130_fd_sc_hd__clkbuf_4
X_11072_ net1182 net870 net834 top.ramstore\[23\] vssd1 vssd1 vccd1 vccd1 _01183_
+ sky130_fd_sc_hd__a22o_1
Xoutput88 net88 vssd1 vssd1 vccd1 vccd1 DAT_O[23] sky130_fd_sc_hd__clkbuf_4
Xoutput99 net99 vssd1 vssd1 vccd1 vccd1 DAT_O[4] sky130_fd_sc_hd__clkbuf_4
X_10023_ net1416 net233 net619 vssd1 vssd1 vccd1 vccd1 _00226_ sky130_fd_sc_hd__mux2_1
XANTENNA__10532__A0 top.DUT.register\[19\]\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_208_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input23_A DAT_I[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06751__A2 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11088__A1 net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_187_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11974_ _05846_ _05850_ _05856_ _05842_ vssd1 vssd1 vccd1 vccd1 _05857_ sky130_fd_sc_hd__a22o_1
XFILLER_0_59_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_604 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_201_3459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12400__RESET_B net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13713_ clknet_leaf_96_clk _01284_ net984 vssd1 vssd1 vccd1 vccd1 top.a1.row2\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_10925_ net1735 net251 net593 vssd1 vssd1 vccd1 vccd1 _01086_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_127_Left_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_196_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_659 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_197_3396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13644_ clknet_leaf_94_clk top.ru.next_write_i net983 vssd1 vssd1 vccd1 vccd1 top.Wen
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10856_ net147 net1969 net595 vssd1 vssd1 vccd1 vccd1 _01017_ sky130_fd_sc_hd__mux2_1
XANTENNA__08384__A _02678_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13575_ clknet_leaf_123_clk net1211 net927 vssd1 vssd1 vccd1 vccd1 net95 sky130_fd_sc_hd__dfrtp_1
XANTENNA__08256__A2 net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10787_ net2143 net161 net485 vssd1 vssd1 vccd1 vccd1 _00948_ sky130_fd_sc_hd__mux2_1
XFILLER_0_183_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12526_ clknet_leaf_71_clk _00118_ vssd1 vssd1 vccd1 vccd1 top.a1.halfData\[3\] sky130_fd_sc_hd__dfxtp_2
XANTENNA__11241__C _05128_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10853__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12457_ clknet_leaf_123_clk _00052_ net926 vssd1 vssd1 vccd1 vccd1 top.ramstore\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_78_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_291 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11408_ _05288_ _05289_ _05290_ vssd1 vssd1 vccd1 vccd1 _05291_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_10_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_136_Left_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12388_ clknet_leaf_103_clk top.ru.next_FetchedInstr\[0\] net976 vssd1 vssd1 vccd1
+ vccd1 top.a1.instruction\[0\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_93_1837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_1848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11339_ top.a1.dataIn\[20\] _05218_ top.a1.dataIn\[21\] vssd1 vssd1 vccd1 vccd1 _05222_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_10_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06990__A2 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11315__A2 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_182_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13009_ clknet_leaf_113_clk _00601_ net991 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[16\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_06880_ top.DUT.register\[7\]\[18\] net517 net514 top.DUT.register\[24\]\[18\] _02018_
+ vssd1 vssd1 vccd1 vccd1 _02019_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_124_2303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09381__C _04438_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06742__A2 net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08550_ _03576_ _03675_ net310 vssd1 vssd1 vccd1 vccd1 _03676_ sky130_fd_sc_hd__mux2_1
XFILLER_0_178_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_145_Left_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_159_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07501_ top.DUT.register\[25\]\[14\] net780 net645 top.DUT.register\[24\]\[14\] _02636_
+ vssd1 vssd1 vccd1 vccd1 _02640_ sky130_fd_sc_hd__a221o_1
XFILLER_0_194_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08481_ _03370_ _03534_ _03598_ vssd1 vssd1 vccd1 vccd1 _03610_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_193_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_175_823 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_374 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07432_ _02568_ _02570_ vssd1 vssd1 vccd1 vccd1 _02571_ sky130_fd_sc_hd__nand2_2
XFILLER_0_57_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_174_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07363_ top.a1.instruction\[29\] net805 _02499_ _02500_ vssd1 vssd1 vccd1 vccd1 _02502_
+ sky130_fd_sc_hd__o2bb2a_2
XTAP_TAPCELL_ROW_170_3002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_1977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09102_ _02349_ _02350_ _02352_ _02354_ vssd1 vssd1 vccd1 vccd1 _04177_ sky130_fd_sc_hd__and4b_1
XFILLER_0_150_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07455__B1 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_794 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06314_ _01332_ _01450_ _01460_ _01333_ vssd1 vssd1 vccd1 vccd1 _01468_ sky130_fd_sc_hd__a31o_1
X_07294_ _02409_ _02430_ vssd1 vssd1 vccd1 vccd1 _02433_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_198_Right_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_150_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06245_ net1245 net854 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedData\[6\] sky130_fd_sc_hd__and2_1
XFILLER_0_72_386 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09033_ _02801_ _02850_ _03612_ _04107_ vssd1 vssd1 vccd1 vccd1 _04108_ sky130_fd_sc_hd__or4_1
XFILLER_0_5_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10763__S net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_154_Left_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09837__B _04514_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout210_A _04780_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_2465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_2476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09747__A2 net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold310 top.DUT.register\[24\]\[23\] vssd1 vssd1 vccd1 vccd1 net1426 sky130_fd_sc_hd__dlygate4sd3_1
X_06176_ top.a1.halfData\[5\] _01416_ vssd1 vssd1 vccd1 vccd1 _01418_ sky130_fd_sc_hd__nor2_1
Xhold321 top.DUT.register\[25\]\[11\] vssd1 vssd1 vccd1 vccd1 net1437 sky130_fd_sc_hd__dlygate4sd3_1
Xhold332 top.DUT.register\[15\]\[12\] vssd1 vssd1 vccd1 vccd1 net1448 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold343 top.DUT.register\[24\]\[15\] vssd1 vssd1 vccd1 vccd1 net1459 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08955__B1 _02304_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold354 top.DUT.register\[23\]\[14\] vssd1 vssd1 vccd1 vccd1 net1470 sky130_fd_sc_hd__dlygate4sd3_1
Xhold365 top.DUT.register\[17\]\[15\] vssd1 vssd1 vccd1 vccd1 net1481 sky130_fd_sc_hd__dlygate4sd3_1
Xhold376 top.DUT.register\[8\]\[2\] vssd1 vssd1 vccd1 vccd1 net1492 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06261__B net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold387 top.DUT.register\[31\]\[3\] vssd1 vssd1 vccd1 vccd1 net1503 sky130_fd_sc_hd__dlygate4sd3_1
Xhold398 top.DUT.register\[10\]\[26\] vssd1 vssd1 vccd1 vccd1 net1514 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout801 net802 vssd1 vssd1 vccd1 vccd1 net801 sky130_fd_sc_hd__clkbuf_2
Xfanout812 _01506_ vssd1 vssd1 vccd1 vccd1 net812 sky130_fd_sc_hd__clkbuf_4
X_09935_ _04930_ _04933_ _04931_ vssd1 vssd1 vccd1 vccd1 _04940_ sky130_fd_sc_hd__a21o_1
Xfanout823 net824 vssd1 vssd1 vccd1 vccd1 net823 sky130_fd_sc_hd__clkbuf_4
Xfanout834 net835 vssd1 vssd1 vccd1 vccd1 net834 sky130_fd_sc_hd__buf_2
XFILLER_0_0_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout677_A _01548_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11306__A2 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout845 _04664_ vssd1 vssd1 vccd1 vccd1 net845 sky130_fd_sc_hd__clkbuf_2
XANTENNA__06981__A2 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout298_X net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout856 net857 vssd1 vssd1 vccd1 vccd1 net856 sky130_fd_sc_hd__buf_2
X_09866_ top.a1.instruction\[25\] net487 net401 top.a1.dataIn\[25\] net397 vssd1 vssd1
+ vccd1 vccd1 _04877_ sky130_fd_sc_hd__a221o_1
Xfanout867 net869 vssd1 vssd1 vccd1 vccd1 net867 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_181_3164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1010 top.DUT.register\[5\]\[11\] vssd1 vssd1 vccd1 vccd1 net2126 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout878 top.lcd.nextState\[2\] vssd1 vssd1 vccd1 vccd1 net878 sky130_fd_sc_hd__clkbuf_2
Xhold1021 top.DUT.register\[9\]\[3\] vssd1 vssd1 vccd1 vccd1 net2137 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout889 net892 vssd1 vssd1 vccd1 vccd1 net889 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09380__B1 _04438_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1032 top.DUT.register\[4\]\[20\] vssd1 vssd1 vccd1 vccd1 net2148 sky130_fd_sc_hd__dlygate4sd3_1
X_08817_ _03909_ _03929_ vssd1 vssd1 vccd1 vccd1 _03931_ sky130_fd_sc_hd__and2_1
Xhold1043 top.DUT.register\[19\]\[27\] vssd1 vssd1 vccd1 vccd1 net2159 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_163_Left_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1054 top.DUT.register\[23\]\[6\] vssd1 vssd1 vccd1 vccd1 net2170 sky130_fd_sc_hd__dlygate4sd3_1
X_09797_ _04453_ net486 net401 top.a1.dataIn\[18\] net397 vssd1 vssd1 vccd1 vccd1
+ _04815_ sky130_fd_sc_hd__a221o_1
XANTENNA__08188__B _03122_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1065 top.ramload\[19\] vssd1 vssd1 vccd1 vccd1 net2181 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06733__A2 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout465_X net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1076 top.DUT.register\[22\]\[9\] vssd1 vssd1 vccd1 vccd1 net2192 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09999__S net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08748_ _02222_ _03863_ vssd1 vssd1 vccd1 vccd1 _03865_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10003__S net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1087 top.DUT.register\[29\]\[31\] vssd1 vssd1 vccd1 vccd1 net2203 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1098 top.DUT.register\[6\]\[15\] vssd1 vssd1 vccd1 vccd1 net2214 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_197_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08679_ net282 _03797_ _03798_ _03793_ vssd1 vssd1 vccd1 vccd1 _03799_ sky130_fd_sc_hd__o211a_1
XFILLER_0_178_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10938__S net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09683__A1 top.a1.instruction\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout632_X net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11623__A top.a1.dataIn\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10710_ net1897 net198 net335 vssd1 vssd1 vccd1 vccd1 _00871_ sky130_fd_sc_hd__mux2_1
XANTENNA__07694__B1 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11690_ _05495_ _05540_ _05572_ _05568_ vssd1 vssd1 vccd1 vccd1 _05573_ sky130_fd_sc_hd__nor4b_1
XFILLER_0_67_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10641_ net214 net2007 net342 vssd1 vssd1 vccd1 vccd1 _00805_ sky130_fd_sc_hd__mux2_1
XANTENNA__09435__A1 net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07446__B1 net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13360_ clknet_leaf_29_clk _00952_ net1017 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[26\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_172_Left_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10572_ net1821 net233 net350 vssd1 vssd1 vccd1 vccd1 _00738_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_165_Right_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12311_ top.pad.button_control.r_counter\[4\] top.pad.button_control.r_counter\[3\]
+ _06114_ vssd1 vssd1 vccd1 vccd1 _06118_ sky130_fd_sc_hd__and3_1
XFILLER_0_63_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_161_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13291_ clknet_leaf_50_clk _00883_ net1059 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[24\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_161_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10673__S net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_263 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09199__B1 top.pc\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12242_ _06075_ _06076_ vssd1 vssd1 vccd1 vccd1 _01322_ sky130_fd_sc_hd__nor2_1
XFILLER_0_210_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06452__A top.a1.instruction\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08946__B1 _02922_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12173_ net1303 net846 net796 _06005_ vssd1 vssd1 vccd1 vccd1 _01281_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_75_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07835__X _02974_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11124_ net906 net1304 net861 _05067_ vssd1 vssd1 vccd1 vccd1 _01213_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_166_2937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11055_ net1217 net866 net837 top.ramstore\[6\] vssd1 vssd1 vccd1 vccd1 _01166_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_181_Left_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12659__CLK clknet_leaf_120_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10006_ net164 top.DUT.register\[3\]\[26\] net624 vssd1 vssd1 vccd1 vccd1 _00211_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_204_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_199_3425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_403 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_199_3436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06724__A2 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_751 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_2033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11236__C _05128_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_203_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11957_ _05831_ net127 _05839_ vssd1 vssd1 vccd1 vccd1 _05840_ sky130_fd_sc_hd__a21o_1
XANTENNA__10848__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10908_ net2266 net200 net481 vssd1 vssd1 vccd1 vccd1 _01069_ sky130_fd_sc_hd__mux2_1
XANTENNA__07685__B1 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11888_ _05734_ _05752_ vssd1 vssd1 vccd1 vccd1 _05771_ sky130_fd_sc_hd__and2_1
XFILLER_0_74_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_184_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13627_ clknet_leaf_75_clk _01214_ net1080 vssd1 vssd1 vccd1 vccd1 net54 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_15_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_692 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10839_ net1705 net191 net475 vssd1 vssd1 vccd1 vccd1 _01000_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_15_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_184_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_4_8__f_clk clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_8__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_171_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07437__B1 net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09938__A net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13558_ clknet_leaf_105_clk _01145_ net969 vssd1 vssd1 vccd1 vccd1 top.ramload\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_132_Right_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12509_ clknet_leaf_78_clk _00101_ net1074 vssd1 vssd1 vccd1 vccd1 top.pc\[21\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__10583__S net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13489_ clknet_leaf_121_clk _01081_ net934 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[31\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09729__A2 net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_2195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09673__A top.a1.instruction\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_2395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07981_ _03113_ _03115_ _03117_ _03119_ vssd1 vssd1 vccd1 vccd1 _03120_ sky130_fd_sc_hd__or4_1
XANTENNA__06963__A2 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09720_ _03548_ net403 net488 _04748_ vssd1 vssd1 vccd1 vccd1 _04749_ sky130_fd_sc_hd__o211a_4
X_06932_ top.DUT.register\[28\]\[21\] net768 net642 top.DUT.register\[8\]\[21\] vssd1
+ vssd1 vccd1 vccd1 _02071_ sky130_fd_sc_hd__a22o_1
X_09651_ _04678_ _04684_ vssd1 vssd1 vccd1 vccd1 _04692_ sky130_fd_sc_hd__nor2_1
X_06863_ _01990_ _01992_ _02001_ vssd1 vssd1 vccd1 vccd1 _02002_ sky130_fd_sc_hd__nor3_1
XANTENNA__09727__A1_N net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08602_ net1629 net833 net803 _03725_ vssd1 vssd1 vccd1 vccd1 _00033_ sky130_fd_sc_hd__a22o_1
X_09582_ _01572_ _04628_ vssd1 vssd1 vccd1 vccd1 _04629_ sky130_fd_sc_hd__and2_1
X_06794_ top.DUT.register\[10\]\[17\] net522 net507 top.DUT.register\[4\]\[17\] vssd1
+ vssd1 vccd1 vccd1 _01933_ sky130_fd_sc_hd__a22o_1
XFILLER_0_49_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08533_ _02477_ _03658_ vssd1 vssd1 vccd1 vccd1 _03660_ sky130_fd_sc_hd__and2_1
XANTENNA__10758__S net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout160_A _04906_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09665__A1 top.a1.halfData\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout258_A _04737_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08464_ _03583_ _03590_ _03593_ vssd1 vssd1 vccd1 vccd1 _03594_ sky130_fd_sc_hd__or3_4
XANTENNA__07676__B1 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_34_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07140__A2 net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12258__B net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_34_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07415_ top.DUT.register\[9\]\[9\] net762 net718 top.DUT.register\[19\]\[9\] vssd1
+ vssd1 vccd1 vccd1 _02554_ sky130_fd_sc_hd__a22o_1
XFILLER_0_174_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_2505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08395_ _03403_ _03407_ net304 vssd1 vssd1 vccd1 vccd1 _03527_ sky130_fd_sc_hd__mux2_1
XFILLER_0_190_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06256__B net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07346_ top.DUT.register\[23\]\[8\] net572 net459 top.DUT.register\[17\]\[8\] vssd1
+ vssd1 vccd1 vccd1 _02485_ sky130_fd_sc_hd__a22o_1
XANTENNA__10493__S net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09567__B _04605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07277_ top.DUT.register\[4\]\[13\] net669 net763 top.DUT.register\[9\]\[13\] _02415_
+ vssd1 vssd1 vccd1 vccd1 _02416_ sky130_fd_sc_hd__a221o_1
XFILLER_0_143_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09016_ _03805_ _04090_ _03948_ _03834_ vssd1 vssd1 vccd1 vccd1 _04091_ sky130_fd_sc_hd__or4b_1
XFILLER_0_14_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06228_ top.ramload\[22\] net858 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedInstr\[22\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_130_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_795 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06159_ top.a1.dataIn\[4\] vssd1 vssd1 vccd1 vccd1 _01402_ sky130_fd_sc_hd__inv_2
Xhold140 top.ramload\[11\] vssd1 vssd1 vccd1 vccd1 net1256 sky130_fd_sc_hd__dlygate4sd3_1
Xhold151 top.ramstore\[6\] vssd1 vssd1 vccd1 vccd1 net1267 sky130_fd_sc_hd__dlygate4sd3_1
Xhold162 top.ramload\[17\] vssd1 vssd1 vccd1 vccd1 net1278 sky130_fd_sc_hd__dlygate4sd3_1
Xhold173 top.a1.row2\[1\] vssd1 vssd1 vccd1 vccd1 net1289 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09583__A _01572_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold184 top.DUT.register\[10\]\[27\] vssd1 vssd1 vccd1 vccd1 net1300 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07600__B1 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold195 top.a1.row2\[19\] vssd1 vssd1 vccd1 vccd1 net1311 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout582_X net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout620 net622 vssd1 vssd1 vccd1 vccd1 net620 sky130_fd_sc_hd__buf_6
Xfanout631 _04714_ vssd1 vssd1 vccd1 vccd1 net631 sky130_fd_sc_hd__clkbuf_8
XANTENNA__06954__A2 net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout642 _01619_ vssd1 vssd1 vccd1 vccd1 net642 sky130_fd_sc_hd__clkbuf_4
X_09918_ _04911_ _04921_ _04924_ vssd1 vssd1 vccd1 vccd1 _04925_ sky130_fd_sc_hd__o21a_1
Xfanout653 _01610_ vssd1 vssd1 vccd1 vccd1 net653 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_148_2667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout664 _01605_ vssd1 vssd1 vccd1 vccd1 net664 sky130_fd_sc_hd__clkbuf_4
Xfanout675 _01548_ vssd1 vssd1 vccd1 vccd1 net675 sky130_fd_sc_hd__buf_4
Xfanout686 _06086_ vssd1 vssd1 vccd1 vccd1 net686 sky130_fd_sc_hd__clkbuf_2
Xfanout697 _03266_ vssd1 vssd1 vccd1 vccd1 net697 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_70_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09849_ top.pc\[23\] _01584_ vssd1 vssd1 vccd1 vccd1 _04862_ sky130_fd_sc_hd__and2_1
XFILLER_0_198_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout847_X net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06706__A2 net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_161_2856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12860_ clknet_leaf_130_clk _00452_ net909 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[11\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_161_2867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11811_ _05667_ net131 _05661_ vssd1 vssd1 vccd1 vccd1 _05694_ sky130_fd_sc_hd__a21boi_1
X_12791_ clknet_leaf_128_clk _00383_ net912 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[9\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10668__S net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09656__A1 top.a1.halfData\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_157_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_205_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11742_ _01399_ _05620_ vssd1 vssd1 vccd1 vccd1 _05625_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07667__B1 net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_194_3355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13307__CLK clknet_leaf_120_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06447__A net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07131__A2 net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11673_ _05554_ _05555_ vssd1 vssd1 vccd1 vccd1 _05556_ sky130_fd_sc_hd__and2_1
XFILLER_0_36_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08933__Y _04041_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13412_ clknet_leaf_36_clk _01004_ net1049 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[28\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_36_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10624_ net158 net1827 net349 vssd1 vssd1 vccd1 vccd1 _00789_ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_684 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13343_ clknet_leaf_19_clk _00935_ net1026 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[26\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_180_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10555_ top.DUT.register\[19\]\[25\] net168 _04988_ vssd1 vssd1 vccd1 vccd1 _00722_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_77_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08631__A2 _03750_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13274_ clknet_leaf_2_clk _00866_ net914 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[24\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_161_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10486_ net1575 net177 net362 vssd1 vssd1 vccd1 vccd1 _00656_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12225_ _06053_ _06058_ vssd1 vssd1 vccd1 vccd1 _06066_ sky130_fd_sc_hd__nand2_1
XFILLER_0_121_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12156_ _06006_ _06028_ _06034_ vssd1 vssd1 vccd1 vccd1 _06039_ sky130_fd_sc_hd__and3_1
XANTENNA__06910__A _02047_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06945__A2 net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11107_ net44 net867 vssd1 vssd1 vccd1 vccd1 _05059_ sky130_fd_sc_hd__and2_1
X_12087_ _05951_ _05968_ vssd1 vssd1 vccd1 vccd1 _05970_ sky130_fd_sc_hd__xnor2_2
X_11038_ net18 net841 net818 top.ramload\[24\] vssd1 vssd1 vccd1 vccd1 _01150_ sky130_fd_sc_hd__a22o_1
XANTENNA__11247__B _01382_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08698__A2 _03441_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09895__A1 top.a1.instruction\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06909__X _02048_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07370__A2 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_201_Right_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10578__S net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12989_ clknet_leaf_13_clk _00581_ net941 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[15\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_145_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07122__A2 net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07200_ net894 _01475_ _01478_ _02338_ vssd1 vssd1 vccd1 vccd1 _02339_ sky130_fd_sc_hd__o31ai_1
XTAP_TAPCELL_ROW_119_2224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08180_ _01809_ net329 vssd1 vssd1 vccd1 vccd1 _03318_ sky130_fd_sc_hd__nand2_1
XFILLER_0_172_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_119_2235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_41_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07131_ top.DUT.register\[6\]\[11\] net567 net563 top.DUT.register\[20\]\[11\] vssd1
+ vssd1 vccd1 vccd1 _02270_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_41_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07062_ top.DUT.register\[15\]\[22\] net707 net699 top.DUT.register\[31\]\[22\] vssd1
+ vssd1 vccd1 vccd1 _02201_ sky130_fd_sc_hd__a22o_1
XFILLER_0_112_211 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_2424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07830__B1 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_4__f_clk_A clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12503__RESET_B net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06936__A2 net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12974__CLK clknet_leaf_40_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07964_ top.DUT.register\[30\]\[31\] net581 net541 top.DUT.register\[8\]\[31\] vssd1
+ vssd1 vccd1 vccd1 _03103_ sky130_fd_sc_hd__a22o_1
XFILLER_0_4_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09690__X _04725_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09703_ top.a1.dataIn\[4\] net795 net798 top.pc\[4\] _04734_ vssd1 vssd1 vccd1 vccd1
+ _04735_ sky130_fd_sc_hd__a221o_1
X_06915_ top.DUT.register\[14\]\[21\] net586 net442 top.DUT.register\[5\]\[21\] _02053_
+ vssd1 vssd1 vccd1 vccd1 _02054_ sky130_fd_sc_hd__a221o_1
XFILLER_0_4_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07895_ top.DUT.register\[8\]\[1\] net541 net449 top.DUT.register\[21\]\[1\] _03033_
+ vssd1 vssd1 vccd1 vccd1 _03034_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout375_A _04981_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09634_ _04674_ _04675_ vssd1 vssd1 vccd1 vccd1 _04676_ sky130_fd_sc_hd__nor2_1
X_06846_ top.DUT.register\[21\]\[19\] net657 net724 top.DUT.register\[29\]\[19\] _01984_
+ vssd1 vssd1 vccd1 vccd1 _01985_ sky130_fd_sc_hd__a221o_1
XANTENNA__09850__B _01584_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07897__B1 net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_143_2586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10488__S net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09565_ top.pc\[29\] _04597_ vssd1 vssd1 vccd1 vccd1 _04613_ sky130_fd_sc_hd__xnor2_1
X_06777_ _01902_ _01906_ _01915_ vssd1 vssd1 vccd1 vccd1 _01916_ sky130_fd_sc_hd__nor3_2
XANTENNA_fanout542_A _01540_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_143_2597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08516_ net286 _03433_ _03438_ net275 vssd1 vssd1 vccd1 vccd1 _03643_ sky130_fd_sc_hd__a22o_1
XANTENNA__07649__B1 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06267__A top.ramload\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09496_ _04529_ _04546_ _04547_ vssd1 vssd1 vccd1 vccd1 _04549_ sky130_fd_sc_hd__nand3_1
XANTENNA__07113__A2 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08447_ _03475_ _03576_ net310 vssd1 vssd1 vccd1 vccd1 _03577_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_176_3085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout807_A net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11323__D top.a1.dataIn\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout428_X net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08378_ _02751_ net500 net494 _02754_ _03506_ vssd1 vssd1 vccd1 vccd1 _03511_ sky130_fd_sc_hd__a221o_1
XFILLER_0_52_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07329_ top.DUT.register\[7\]\[12\] net659 net702 top.DUT.register\[3\]\[12\] _02467_
+ vssd1 vssd1 vccd1 vccd1 _02468_ sky130_fd_sc_hd__a221o_1
XFILLER_0_116_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08613__A2 _03534_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_190_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10340_ net2241 net219 net377 vssd1 vssd1 vccd1 vccd1 _00516_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_59_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07821__B1 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_143_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout797_X net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10271_ net1433 net237 net386 vssd1 vssd1 vccd1 vccd1 _00449_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10951__S net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12010_ _05887_ _05888_ _05890_ _05891_ vssd1 vssd1 vccd1 vccd1 _05893_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_103_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_72_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout964_X net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06927__A2 net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout450 _01562_ vssd1 vssd1 vccd1 vccd1 net450 sky130_fd_sc_hd__buf_2
XANTENNA__08129__A1 net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout461 net462 vssd1 vssd1 vccd1 vccd1 net461 sky130_fd_sc_hd__clkbuf_8
XANTENNA__08129__B2 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout472 _05104_ vssd1 vssd1 vccd1 vccd1 net472 sky130_fd_sc_hd__buf_2
Xfanout483 _04962_ vssd1 vssd1 vccd1 vccd1 net483 sky130_fd_sc_hd__clkbuf_4
Xfanout494 net495 vssd1 vssd1 vccd1 vccd1 net494 sky130_fd_sc_hd__clkbuf_4
X_12912_ clknet_leaf_26_clk _00504_ net1011 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[12\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07888__B1 net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07352__A2 net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12843_ clknet_leaf_47_clk _00435_ net1069 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[10\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_17_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10398__S net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_220 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06448__Y _01587_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_439 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_562 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_4_15__f_clk_A clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12774_ clknet_leaf_33_clk _00366_ net1046 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[8\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06177__A net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07104__A2 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11725_ _05540_ _05571_ vssd1 vssd1 vccd1 vccd1 _05608_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_83_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_194_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_139_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11656_ _05492_ _05538_ vssd1 vssd1 vccd1 vccd1 _05539_ sky130_fd_sc_hd__nand2_1
XANTENNA__06464__X _01603_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10607_ net222 net2202 net346 vssd1 vssd1 vccd1 vccd1 _00772_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_211_3609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11587_ _05453_ _05460_ _05465_ vssd1 vssd1 vccd1 vccd1 _05470_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_3_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13326_ clknet_leaf_41_clk _00918_ net1047 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[25\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
Xmax_cap606 _04957_ vssd1 vssd1 vccd1 vccd1 net606 sky130_fd_sc_hd__buf_2
XFILLER_0_107_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10538_ net1596 net236 net354 vssd1 vssd1 vccd1 vccd1 _00705_ sky130_fd_sc_hd__mux2_1
Xhold909 top.DUT.register\[30\]\[1\] vssd1 vssd1 vccd1 vccd1 net2025 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_114_2154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12415__Q top.a1.instruction\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13257_ clknet_leaf_51_clk _00849_ net1058 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[23\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10861__S net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10469_ net2231 net244 net361 vssd1 vssd1 vccd1 vccd1 _00639_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12208_ _06053_ vssd1 vssd1 vccd1 vccd1 _06054_ sky130_fd_sc_hd__inv_2
X_13188_ clknet_leaf_35_clk _00780_ net1049 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[21\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06918__A2 net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12139_ _06020_ _06021_ vssd1 vssd1 vccd1 vccd1 _06022_ sky130_fd_sc_hd__and2b_1
XFILLER_0_209_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07591__A2 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_208_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09868__A1 top.pc\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_205_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06700_ top.DUT.register\[29\]\[25\] net451 net508 top.DUT.register\[4\]\[25\] vssd1
+ vssd1 vccd1 vccd1 _01839_ sky130_fd_sc_hd__a22o_1
X_07680_ top.DUT.register\[12\]\[4\] net740 net712 top.DUT.register\[11\]\[4\] vssd1
+ vssd1 vccd1 vccd1 _02819_ sky130_fd_sc_hd__a22o_1
XANTENNA__07343__A2 net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06631_ top.DUT.register\[28\]\[27\] net768 net720 top.DUT.register\[19\]\[27\] vssd1
+ vssd1 vccd1 vccd1 _01770_ sky130_fd_sc_hd__a22o_1
XANTENNA__06551__B1 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09350_ top.pc\[15\] _04377_ top.pc\[16\] vssd1 vssd1 vccd1 vccd1 _04411_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10101__S net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06562_ _01699_ _01700_ vssd1 vssd1 vccd1 vccd1 _01701_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_176_236 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08301_ net286 _03434_ _03435_ net274 _03433_ vssd1 vssd1 vccd1 vccd1 _03436_ sky130_fd_sc_hd__a32o_1
XFILLER_0_164_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_426 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_595 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09281_ _04331_ _04332_ _04329_ vssd1 vssd1 vccd1 vccd1 _04346_ sky130_fd_sc_hd__a21o_1
X_06493_ top.DUT.register\[25\]\[30\] net780 net772 top.DUT.register\[10\]\[30\] vssd1
+ vssd1 vccd1 vccd1 _01632_ sky130_fd_sc_hd__a22o_1
XFILLER_0_185_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_191_239 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08232_ net288 _03194_ vssd1 vssd1 vccd1 vccd1 _03369_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06374__X _01513_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08163_ _02112_ net329 vssd1 vssd1 vccd1 vccd1 _03301_ sky130_fd_sc_hd__or2_1
XFILLER_0_172_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12755__RESET_B net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09685__X _04721_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07114_ top.DUT.register\[26\]\[16\] net751 net711 top.DUT.register\[11\]\[16\] vssd1
+ vssd1 vccd1 vccd1 _02253_ sky130_fd_sc_hd__a22o_1
XANTENNA__07803__B1 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08094_ _02849_ net300 vssd1 vssd1 vccd1 vccd1 _03233_ sky130_fd_sc_hd__nand2_1
XFILLER_0_31_827 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_542 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload60 clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 clkload60/Y sky130_fd_sc_hd__clkinv_2
Xclkload71 clknet_leaf_30_clk vssd1 vssd1 vccd1 vccd1 clkload71/Y sky130_fd_sc_hd__clkinv_8
XANTENNA__10771__S net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07045_ top.DUT.register\[10\]\[22\] net522 net444 top.DUT.register\[1\]\[22\] vssd1
+ vssd1 vccd1 vccd1 _02184_ sky130_fd_sc_hd__a22o_1
Xclkload82 clknet_leaf_44_clk vssd1 vssd1 vccd1 vccd1 clkload82/Y sky130_fd_sc_hd__clkinv_8
XFILLER_0_30_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1032_A net1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06821__Y _01960_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload93 clknet_leaf_70_clk vssd1 vssd1 vccd1 vccd1 clkload93/Y sky130_fd_sc_hd__inv_16
XANTENNA_fanout492_A _03339_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08996_ _03920_ _03941_ _03960_ _03979_ vssd1 vssd1 vccd1 vccd1 _04071_ sky130_fd_sc_hd__or4_1
XANTENNA__07582__A2 net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09308__B1 _04370_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_2615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09861__A net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_2626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07947_ _03082_ _03085_ _02136_ vssd1 vssd1 vccd1 vccd1 _03086_ sky130_fd_sc_hd__o21ai_1
XANTENNA__06790__B1 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout378_X net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout757_A _01620_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_339 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07878_ top.DUT.register\[7\]\[1\] net660 net704 top.DUT.register\[3\]\[1\] _03016_
+ vssd1 vssd1 vccd1 vccd1 _03017_ sky130_fd_sc_hd__a221o_1
XANTENNA__08477__A net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07334__A2 _02472_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_178_3114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09617_ top.a1.state\[1\] top.a1.state\[0\] top.a1.state\[2\] vssd1 vssd1 vccd1 vccd1
+ _04662_ sky130_fd_sc_hd__nor3b_1
XANTENNA__11130__A3 net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06829_ top.DUT.register\[8\]\[19\] net542 net445 top.DUT.register\[1\]\[19\] _01967_
+ vssd1 vssd1 vccd1 vccd1 _01968_ sky130_fd_sc_hd__a221o_1
XANTENNA__06542__B1 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout545_X net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_167_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09548_ top.pc\[27\] top.pc\[28\] _04567_ vssd1 vssd1 vccd1 vccd1 _04597_ sky130_fd_sc_hd__and3_1
XANTENNA__10011__S net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_167_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_191_3314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_183_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08295__B1 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10946__S net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout712_X net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09479_ net133 _04526_ _04527_ _04532_ net811 vssd1 vssd1 vccd1 vccd1 _04533_ sky130_fd_sc_hd__o32a_1
XFILLER_0_136_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_792 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11510_ _05392_ vssd1 vssd1 vccd1 vccd1 _05393_ sky130_fd_sc_hd__inv_2
XFILLER_0_108_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12490_ clknet_leaf_86_clk _00082_ net1006 vssd1 vssd1 vccd1 vccd1 top.pc\[2\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_108_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11441_ _05306_ _05314_ _05316_ _05317_ _05323_ vssd1 vssd1 vccd1 vccd1 _05324_ sky130_fd_sc_hd__o41ai_2
XTAP_TAPCELL_ROW_22_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_156_2788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12496__RESET_B net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09795__B1 net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11372_ top.a1.dataIn\[18\] _05252_ _05253_ vssd1 vssd1 vccd1 vccd1 _05255_ sky130_fd_sc_hd__or3_1
XFILLER_0_150_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13111_ clknet_leaf_2_clk _00703_ net918 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[19\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_10323_ net160 net2021 net383 vssd1 vssd1 vccd1 vccd1 _00500_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10681__S net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_189_3276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_189_3287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13042_ clknet_leaf_23_clk _00634_ net1015 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[17\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_10254_ net172 net2175 net390 vssd1 vssd1 vccd1 vccd1 _00433_ sky130_fd_sc_hd__mux2_1
X_10185_ top.a1.instruction\[9\] _04156_ net690 _04711_ vssd1 vssd1 vccd1 vccd1 _04965_
+ sky130_fd_sc_hd__or4_4
XFILLER_0_56_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07573__A2 net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_208_3560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_208_3571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout280 _03239_ vssd1 vssd1 vccd1 vccd1 net280 sky130_fd_sc_hd__clkbuf_2
Xfanout291 net292 vssd1 vssd1 vccd1 vccd1 net291 sky130_fd_sc_hd__buf_2
XFILLER_0_89_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_202_800 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07325__A2 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12826_ clknet_leaf_5_clk _00418_ net936 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[10\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_201_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10856__S net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12757_ clknet_leaf_31_clk _00349_ net1020 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[8\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_167_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06906__Y _02045_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11708_ _05562_ _05590_ vssd1 vssd1 vccd1 vccd1 _05591_ sky130_fd_sc_hd__and2b_1
XFILLER_0_84_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12688_ clknet_leaf_28_clk _00280_ net1010 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[5\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_181_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11639_ _05503_ _05521_ vssd1 vssd1 vccd1 vccd1 _05522_ sky130_fd_sc_hd__xnor2_1
XANTENNA__13025__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_626 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08589__B2 net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_3_clk_A clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold706 top.DUT.register\[8\]\[16\] vssd1 vssd1 vccd1 vccd1 net1822 sky130_fd_sc_hd__dlygate4sd3_1
Xhold717 top.DUT.register\[17\]\[8\] vssd1 vssd1 vccd1 vccd1 net1833 sky130_fd_sc_hd__dlygate4sd3_1
X_13309_ clknet_leaf_127_clk _00901_ net930 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[25\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold728 top.DUT.register\[24\]\[16\] vssd1 vssd1 vccd1 vccd1 net1844 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_96_1879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10591__S net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold739 top.DUT.register\[27\]\[30\] vssd1 vssd1 vccd1 vccd1 net1855 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13175__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08850_ _01789_ net493 _03427_ _03922_ _03961_ vssd1 vssd1 vccd1 vccd1 _03962_ sky130_fd_sc_hd__o221a_1
X_07801_ top.DUT.register\[21\]\[2\] net447 net439 top.DUT.register\[5\]\[2\] _02939_
+ vssd1 vssd1 vccd1 vccd1 _02940_ sky130_fd_sc_hd__a221o_1
XANTENNA__09681__A net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08781_ _03894_ _03895_ vssd1 vssd1 vccd1 vccd1 _03896_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_127_2345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06772__B1 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_2356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07732_ top.DUT.register\[10\]\[3\] net772 net732 top.DUT.register\[14\]\[3\] vssd1
+ vssd1 vccd1 vccd1 _02871_ sky130_fd_sc_hd__a22o_1
XANTENNA__07316__A2 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_196_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11112__A3 net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09710__B1 net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07663_ _02801_ vssd1 vssd1 vccd1 vccd1 _02802_ sky130_fd_sc_hd__inv_2
XANTENNA__06524__B1 net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09402_ net900 top.pc\[18\] _04460_ net891 vssd1 vssd1 vccd1 vccd1 _00098_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_140_2545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06614_ top.DUT.register\[8\]\[27\] net541 net442 top.DUT.register\[5\]\[27\] _01752_
+ vssd1 vssd1 vccd1 vccd1 _01753_ sky130_fd_sc_hd__a221o_1
XFILLER_0_177_534 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07594_ top.DUT.register\[9\]\[6\] net762 net758 top.DUT.register\[30\]\[6\] vssd1
+ vssd1 vccd1 vccd1 _02733_ sky130_fd_sc_hd__a22o_1
XFILLER_0_149_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_165_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09333_ top.pc\[15\] _04377_ vssd1 vssd1 vccd1 vccd1 _04395_ sky130_fd_sc_hd__xnor2_1
X_06545_ top.DUT.register\[25\]\[29\] net780 net768 top.DUT.register\[28\]\[29\] vssd1
+ vssd1 vccd1 vccd1 _01684_ sky130_fd_sc_hd__a22o_1
XFILLER_0_165_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_96 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_126_clk clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_126_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__10766__S net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout338_A _04993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_173_3044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_559 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09264_ top.pc\[11\] _02365_ vssd1 vssd1 vccd1 vccd1 _04330_ sky130_fd_sc_hd__and2b_1
X_06476_ _01604_ _01607_ net792 vssd1 vssd1 vccd1 vccd1 _01615_ sky130_fd_sc_hd__and3b_1
XFILLER_0_47_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08215_ _03344_ _03351_ _03352_ vssd1 vssd1 vccd1 vccd1 _03353_ sky130_fd_sc_hd__or3_2
XFILLER_0_172_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09226__C1 net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09195_ _04246_ _04264_ _04263_ vssd1 vssd1 vccd1 vccd1 _04266_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout505_A net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06264__B net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11179__A3 net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08146_ _03276_ _03283_ net312 vssd1 vssd1 vccd1 vccd1 _03284_ sky130_fd_sc_hd__mux2_1
X_08077_ _03214_ _03215_ vssd1 vssd1 vccd1 vccd1 _03216_ sky130_fd_sc_hd__nand2_1
X_07028_ _02159_ _02160_ _02162_ _02164_ vssd1 vssd1 vccd1 vccd1 _02167_ sky130_fd_sc_hd__or4_1
XFILLER_0_101_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout874_A net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_80 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout495_X net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13724__RESET_B net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10006__S net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07555__A2 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold11 top.a1.dataInTemp\[1\] vssd1 vssd1 vccd1 vccd1 net1127 sky130_fd_sc_hd__dlygate4sd3_1
Xhold22 top.a1.dataInTemp\[9\] vssd1 vssd1 vccd1 vccd1 net1138 sky130_fd_sc_hd__dlygate4sd3_1
Xhold33 top.ramstore\[31\] vssd1 vssd1 vccd1 vccd1 net1149 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout662_X net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold44 top.a1.data\[10\] vssd1 vssd1 vccd1 vccd1 net1160 sky130_fd_sc_hd__dlygate4sd3_1
X_08979_ _03510_ _03522_ _04053_ vssd1 vssd1 vccd1 vccd1 _04054_ sky130_fd_sc_hd__or3b_1
XANTENNA__06763__B1 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold55 top.a1.dataInTemp\[11\] vssd1 vssd1 vccd1 vccd1 net1171 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08919__B _04027_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold66 net88 vssd1 vssd1 vccd1 vccd1 net1182 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_194_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07382__Y _02521_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold77 net74 vssd1 vssd1 vccd1 vccd1 net1193 sky130_fd_sc_hd__dlygate4sd3_1
X_11990_ _05865_ _05872_ vssd1 vssd1 vccd1 vccd1 _05873_ sky130_fd_sc_hd__nand2_1
Xhold88 top.ramload\[15\] vssd1 vssd1 vccd1 vccd1 net1204 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06279__X _01442_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold99 _01165_ vssd1 vssd1 vccd1 vccd1 net1215 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07307__A2 net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10941_ net1716 net194 net592 vssd1 vssd1 vccd1 vccd1 _01102_ sky130_fd_sc_hd__mux2_1
XFILLER_0_196_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_168_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_67_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_203_3490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13660_ clknet_leaf_91_clk _01236_ net996 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[106\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_27_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10872_ net223 net1607 net595 vssd1 vssd1 vccd1 vccd1 _01033_ sky130_fd_sc_hd__mux2_1
XFILLER_0_195_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12611_ clknet_leaf_49_clk _00203_ net1061 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[3\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_158_2817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_183_515 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13591_ clknet_leaf_63_clk net1135 net1092 vssd1 vssd1 vccd1 vccd1 net82 sky130_fd_sc_hd__dfrtp_1
XANTENNA__13048__CLK clknet_leaf_128_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_117_clk clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_117_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__10676__S net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10529__X _04989_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_210_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_239 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_111 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12542_ clknet_leaf_54_clk _00134_ net1031 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[1\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06455__A top.a1.instruction\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12473_ clknet_leaf_64_clk _00068_ net1090 vssd1 vssd1 vccd1 vccd1 top.ramstore\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_49_Left_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_191_592 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_579 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11424_ _05267_ _05285_ vssd1 vssd1 vccd1 vccd1 _05307_ sky130_fd_sc_hd__nand2_1
XFILLER_0_22_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08670__A _02007_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_8 _01513_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11355_ _05207_ _05214_ _05218_ vssd1 vssd1 vccd1 vccd1 _05238_ sky130_fd_sc_hd__a21o_1
XANTENNA__09485__B _01584_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_2113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07794__A2 net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10306_ net227 top.DUT.register\[12\]\[10\] net381 vssd1 vssd1 vccd1 vccd1 _00483_
+ sky130_fd_sc_hd__mux2_1
X_11286_ top.a1.row2\[35\] _05140_ _05149_ top.a1.row1\[123\] _05170_ vssd1 vssd1
+ vccd1 vccd1 _05176_ sky130_fd_sc_hd__a221o_1
XFILLER_0_67_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13025_ clknet_leaf_16_clk _00617_ net961 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[16\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_169_2979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10237_ net248 net2045 net389 vssd1 vssd1 vccd1 vccd1 _00416_ sky130_fd_sc_hd__mux2_1
XANTENNA__07546__A2 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1020 net1025 vssd1 vssd1 vccd1 vccd1 net1020 sky130_fd_sc_hd__buf_2
Xfanout1031 net1032 vssd1 vssd1 vccd1 vccd1 net1031 sky130_fd_sc_hd__clkbuf_4
Xfanout1042 net1043 vssd1 vssd1 vccd1 vccd1 net1042 sky130_fd_sc_hd__clkbuf_4
Xfanout1053 net1055 vssd1 vssd1 vccd1 vccd1 net1053 sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_58_Left_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10168_ net1688 net182 net603 vssd1 vssd1 vccd1 vccd1 _00367_ sky130_fd_sc_hd__mux2_1
XANTENNA__06754__B1 net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1064 net1070 vssd1 vssd1 vccd1 vccd1 net1064 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11536__A top.a1.dataIn\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1075 net1087 vssd1 vssd1 vccd1 vccd1 net1075 sky130_fd_sc_hd__clkbuf_4
Xfanout1086 net1087 vssd1 vssd1 vccd1 vccd1 net1086 sky130_fd_sc_hd__buf_2
Xfanout1097 net1098 vssd1 vssd1 vccd1 vccd1 net1097 sky130_fd_sc_hd__clkbuf_4
X_10099_ net1512 net185 net613 vssd1 vssd1 vccd1 vccd1 _00300_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_635 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_109_2075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_2086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11255__B _05128_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06506__B1 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_179_Right_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_122_2275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12809_ clknet_leaf_53_clk _00401_ net1038 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[9\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10586__S net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_108_clk clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_108_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_123_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13789_ clknet_leaf_68_clk _01358_ vssd1 vssd1 vccd1 vccd1 top.pad.button_control.r_counter\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_06330_ top.a1.instruction\[13\] net893 vssd1 vssd1 vccd1 vccd1 _01477_ sky130_fd_sc_hd__nor2_2
XFILLER_0_8_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08056__S net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_199_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_535 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_1919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06261_ top.ramload\[22\] net853 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedData\[22\]
+ sky130_fd_sc_hd__and2_1
XANTENNA__06285__A2 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08000_ top.DUT.register\[10\]\[31\] net772 net728 top.DUT.register\[18\]\[31\] _03138_
+ vssd1 vssd1 vccd1 vccd1 _03139_ sky130_fd_sc_hd__a221o_1
XANTENNA__09759__B1 _04752_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06192_ _00008_ top.a1.nextHex\[7\] vssd1 vssd1 vccd1 vccd1 top.a1.nextHex\[4\] sky130_fd_sc_hd__or2_1
XFILLER_0_40_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_787 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold503 top.DUT.register\[2\]\[13\] vssd1 vssd1 vccd1 vccd1 net1619 sky130_fd_sc_hd__dlygate4sd3_1
Xhold514 top.DUT.register\[11\]\[18\] vssd1 vssd1 vccd1 vccd1 net1630 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold525 top.DUT.register\[19\]\[9\] vssd1 vssd1 vccd1 vccd1 net1641 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08431__B1 _03560_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold536 top.DUT.register\[7\]\[12\] vssd1 vssd1 vccd1 vccd1 net1652 sky130_fd_sc_hd__dlygate4sd3_1
Xhold547 top.DUT.register\[6\]\[21\] vssd1 vssd1 vccd1 vccd1 net1663 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07785__A2 _02904_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold558 top.DUT.register\[24\]\[28\] vssd1 vssd1 vccd1 vccd1 net1674 sky130_fd_sc_hd__dlygate4sd3_1
X_09951_ net1616 net243 net627 vssd1 vssd1 vccd1 vccd1 _00159_ sky130_fd_sc_hd__mux2_1
Xhold569 top.DUT.register\[16\]\[19\] vssd1 vssd1 vccd1 vccd1 net1685 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06993__B1 net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08902_ net884 top.pc\[29\] net695 _04011_ vssd1 vssd1 vccd1 vccd1 _04012_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_51_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09882_ top.a1.instruction\[26\] net486 net402 top.a1.dataIn\[26\] _04753_ vssd1
+ vssd1 vccd1 vccd1 _04892_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_5_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07537__A2 net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08833_ net435 _03941_ _03945_ net427 _03944_ vssd1 vssd1 vccd1 vccd1 _03946_ sky130_fd_sc_hd__a221o_1
XANTENNA__07924__A _02409_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout190_A net191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06745__B1 net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout288_A net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11446__A top.a1.dataIn\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08764_ net434 _03879_ vssd1 vssd1 vccd1 vccd1 _03880_ sky130_fd_sc_hd__nor2_1
XFILLER_0_197_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07715_ top.a1.instruction\[23\] _01507_ net793 top.a1.instruction\[15\] _02853_
+ vssd1 vssd1 vccd1 vccd1 _02854_ sky130_fd_sc_hd__a221o_2
X_08695_ _02179_ _03813_ vssd1 vssd1 vccd1 vccd1 _03814_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout455_A _01553_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_196_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06259__B net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07646_ top.DUT.register\[7\]\[5\] net659 net719 top.DUT.register\[19\]\[5\] vssd1
+ vssd1 vccd1 vccd1 _02785_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_146_Right_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_24_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07577_ top.DUT.register\[28\]\[6\] net555 net439 top.DUT.register\[5\]\[6\] vssd1
+ vssd1 vccd1 vccd1 _02716_ sky130_fd_sc_hd__a22o_1
XANTENNA__10496__S net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_192_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_576 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09316_ _04377_ _04378_ vssd1 vssd1 vccd1 vccd1 _04379_ sky130_fd_sc_hd__or2_1
X_06528_ top.DUT.register\[7\]\[29\] net517 net513 top.DUT.register\[24\]\[29\] _01666_
+ vssd1 vssd1 vccd1 vccd1 _01667_ sky130_fd_sc_hd__a221o_1
XFILLER_0_146_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_192_367 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09247_ top.pc\[10\] _02547_ vssd1 vssd1 vccd1 vccd1 _04314_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_7_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06459_ top.a1.instruction\[20\] top.a1.instruction\[21\] top.a1.instruction\[24\]
+ net792 vssd1 vssd1 vccd1 vccd1 _01598_ sky130_fd_sc_hd__o31a_2
XFILLER_0_105_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout508_X net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_153_2736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_153_2747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09178_ _04245_ _04248_ _04249_ vssd1 vssd1 vccd1 vccd1 _04250_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout991_A net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08129_ net886 top.pc\[0\] _03265_ net697 vssd1 vssd1 vccd1 vccd1 _03268_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_186_3235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07776__A2 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11140_ net907 net1760 net862 _05075_ vssd1 vssd1 vccd1 vccd1 _01221_ sky130_fd_sc_hd__a31o_1
XANTENNA__08973__B2 net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout877_X net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06984__B1 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput45 net45 vssd1 vssd1 vccd1 vccd1 ADR_O[14] sky130_fd_sc_hd__buf_2
XANTENNA__12513__Q top.pc\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput56 net56 vssd1 vssd1 vccd1 vccd1 ADR_O[24] sky130_fd_sc_hd__buf_2
Xoutput67 net67 vssd1 vssd1 vccd1 vccd1 ADR_O[5] sky130_fd_sc_hd__buf_2
Xoutput78 net78 vssd1 vssd1 vccd1 vccd1 DAT_O[14] sky130_fd_sc_hd__clkbuf_4
X_11071_ net87 net872 net836 net1173 vssd1 vssd1 vccd1 vccd1 _01182_ sky130_fd_sc_hd__a22o_1
Xoutput89 net89 vssd1 vssd1 vccd1 vccd1 DAT_O[24] sky130_fd_sc_hd__clkbuf_4
XANTENNA__07528__A2 net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10022_ net1569 net236 net622 vssd1 vssd1 vccd1 vccd1 _00225_ sky130_fd_sc_hd__mux2_1
XANTENNA__07834__A net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08649__B _02049_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_208_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input16_A DAT_I[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11973_ _05845_ _05855_ vssd1 vssd1 vccd1 vccd1 _05856_ sky130_fd_sc_hd__nand2_1
XANTENNA__08489__B1 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06169__B top.a1.halfData\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_616 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10924_ net1943 net257 net592 vssd1 vssd1 vccd1 vccd1 _01085_ sky130_fd_sc_hd__mux2_1
X_13712_ clknet_leaf_96_clk _01283_ net985 vssd1 vssd1 vccd1 vccd1 top.a1.row2\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07161__B1 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_113_Right_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_197_3397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_195_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13643_ clknet_leaf_94_clk _00010_ net994 vssd1 vssd1 vccd1 vccd1 top.ru.state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_10855_ net1254 net143 net475 vssd1 vssd1 vccd1 vccd1 _01016_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_16_clk_X clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13574_ clknet_leaf_63_clk net1177 net1090 vssd1 vssd1 vccd1 vccd1 net84 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10786_ net2168 net165 net485 vssd1 vssd1 vccd1 vccd1 _00947_ sky130_fd_sc_hd__mux2_1
XFILLER_0_183_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_171_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12525_ clknet_leaf_70_clk _00117_ vssd1 vssd1 vccd1 vccd1 top.a1.halfData\[2\] sky130_fd_sc_hd__dfxtp_2
XANTENNA__11260__A2 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08661__B1 _03777_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12456_ clknet_leaf_46_clk _00051_ net1066 vssd1 vssd1 vccd1 vccd1 top.ramstore\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11407_ _05285_ _05256_ vssd1 vssd1 vccd1 vccd1 _05290_ sky130_fd_sc_hd__and2b_1
XFILLER_0_78_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12387_ clknet_leaf_110_clk top.ru.next_FetchedData\[31\] net989 vssd1 vssd1 vccd1
+ vccd1 top.a1.dataIn\[31\] sky130_fd_sc_hd__dfrtp_2
XANTENNA__09610__C1 net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_1838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07767__A2 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11338_ top.a1.dataIn\[21\] top.a1.dataIn\[20\] _05218_ vssd1 vssd1 vccd1 vccd1 _05221_
+ sky130_fd_sc_hd__or3_1
XFILLER_0_120_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06975__B1 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09943__B top.a1.instruction\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11269_ _05156_ _05157_ _05158_ _05160_ vssd1 vssd1 vccd1 vccd1 _05161_ sky130_fd_sc_hd__or4_2
XFILLER_0_94_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13008_ clknet_leaf_31_clk _00600_ net1018 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[15\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06727__B1 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_175_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_124_2304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07500_ top.DUT.register\[13\]\[14\] net777 net719 top.DUT.register\[19\]\[14\] vssd1
+ vssd1 vccd1 vccd1 _02639_ sky130_fd_sc_hd__a22o_1
XANTENNA__12528__RESET_B net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08480_ _02389_ net494 _03607_ _03608_ vssd1 vssd1 vccd1 vccd1 _03609_ sky130_fd_sc_hd__a211o_1
XANTENNA__07152__B1 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07431_ _02569_ vssd1 vssd1 vccd1 vccd1 _02570_ sky130_fd_sc_hd__inv_2
XFILLER_0_175_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_159_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06366__Y _01505_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07362_ top.a1.instruction\[29\] net789 net794 top.a1.instruction\[21\] vssd1 vssd1
+ vccd1 vccd1 _02501_ sky130_fd_sc_hd__a22o_1
XFILLER_0_73_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_170_3003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_1978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09101_ _04175_ _04174_ _04142_ vssd1 vssd1 vccd1 vccd1 _04176_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06313_ _01331_ _01463_ _01467_ _01449_ vssd1 vssd1 vccd1 vccd1 _00002_ sky130_fd_sc_hd__o22a_1
XFILLER_0_174_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_155_581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07293_ _02431_ vssd1 vssd1 vccd1 vccd1 _02432_ sky130_fd_sc_hd__inv_2
X_09032_ _02135_ _03143_ _03187_ _04064_ vssd1 vssd1 vccd1 vccd1 _04107_ sky130_fd_sc_hd__or4_1
XFILLER_0_32_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06244_ net1274 net854 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedData\[5\] sky130_fd_sc_hd__and2_1
XFILLER_0_143_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_150_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06823__A _01940_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_398 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_2466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_2477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold300 top.DUT.register\[4\]\[9\] vssd1 vssd1 vccd1 vccd1 net1416 sky130_fd_sc_hd__dlygate4sd3_1
X_06175_ top.a1.halfData\[5\] _01416_ vssd1 vssd1 vccd1 vccd1 _01417_ sky130_fd_sc_hd__or2_1
Xhold311 top.DUT.register\[19\]\[24\] vssd1 vssd1 vccd1 vccd1 net1427 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout203_A net206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold322 top.DUT.register\[30\]\[30\] vssd1 vssd1 vccd1 vccd1 net1438 sky130_fd_sc_hd__dlygate4sd3_1
Xhold333 top.DUT.register\[25\]\[17\] vssd1 vssd1 vccd1 vccd1 net1449 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07758__A2 net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08955__B2 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold344 top.DUT.register\[15\]\[14\] vssd1 vssd1 vccd1 vccd1 net1460 sky130_fd_sc_hd__dlygate4sd3_1
Xhold355 top.DUT.register\[20\]\[26\] vssd1 vssd1 vccd1 vccd1 net1471 sky130_fd_sc_hd__dlygate4sd3_1
Xhold366 top.DUT.register\[14\]\[8\] vssd1 vssd1 vccd1 vccd1 net1482 sky130_fd_sc_hd__dlygate4sd3_1
Xhold377 top.DUT.register\[17\]\[10\] vssd1 vssd1 vccd1 vccd1 net1493 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold388 top.DUT.register\[6\]\[26\] vssd1 vssd1 vccd1 vccd1 net1504 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout802 _03269_ vssd1 vssd1 vccd1 vccd1 net802 sky130_fd_sc_hd__clkbuf_2
Xhold399 top.DUT.register\[13\]\[26\] vssd1 vssd1 vccd1 vccd1 net1515 sky130_fd_sc_hd__dlygate4sd3_1
X_09934_ _04045_ net407 vssd1 vssd1 vccd1 vccd1 _04939_ sky130_fd_sc_hd__nand2_1
XANTENNA__06430__A2 net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout813 net814 vssd1 vssd1 vccd1 vccd1 net813 sky130_fd_sc_hd__clkbuf_4
Xfanout824 net825 vssd1 vssd1 vccd1 vccd1 net824 sky130_fd_sc_hd__buf_2
Xfanout835 net836 vssd1 vssd1 vccd1 vccd1 net835 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__10999__B net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout846 net847 vssd1 vssd1 vccd1 vccd1 net846 sky130_fd_sc_hd__buf_2
XANTENNA__09904__B1 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09865_ net1739 net174 net634 vssd1 vssd1 vccd1 vccd1 _00145_ sky130_fd_sc_hd__mux2_1
Xfanout857 top.ru.next_iready vssd1 vssd1 vccd1 vccd1 net857 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_input8_A DAT_I[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06718__B1 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1000 top.DUT.register\[10\]\[31\] vssd1 vssd1 vccd1 vccd1 net2116 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_181_3154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout572_A _01519_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout868 net869 vssd1 vssd1 vccd1 vccd1 net868 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_181_3165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1011 top.DUT.register\[29\]\[22\] vssd1 vssd1 vccd1 vccd1 net2127 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout879 top.lcd.nextState\[2\] vssd1 vssd1 vccd1 vccd1 net879 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09380__A1 _01930_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1022 top.a1.hexop\[2\] vssd1 vssd1 vccd1 vccd1 net2138 sky130_fd_sc_hd__dlygate4sd3_1
X_08816_ _03909_ _03929_ vssd1 vssd1 vccd1 vccd1 _03930_ sky130_fd_sc_hd__nor2_1
Xhold1033 top.DUT.register\[31\]\[30\] vssd1 vssd1 vccd1 vccd1 net2149 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1044 top.DUT.register\[7\]\[2\] vssd1 vssd1 vccd1 vccd1 net2160 sky130_fd_sc_hd__dlygate4sd3_1
X_09796_ net1562 net215 net632 vssd1 vssd1 vccd1 vccd1 _00138_ sky130_fd_sc_hd__mux2_1
XANTENNA__07391__B1 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1055 top.DUT.register\[16\]\[23\] vssd1 vssd1 vccd1 vccd1 net2171 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1066 top.DUT.register\[11\]\[6\] vssd1 vssd1 vccd1 vccd1 net2182 sky130_fd_sc_hd__dlygate4sd3_1
X_08747_ _03863_ vssd1 vssd1 vccd1 vccd1 _03864_ sky130_fd_sc_hd__inv_2
Xhold1077 top.DUT.register\[2\]\[25\] vssd1 vssd1 vccd1 vccd1 net2193 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_90_clk_A clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1088 top.pad.keyCode\[5\] vssd1 vssd1 vccd1 vccd1 net2204 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout360_X net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1099 top.DUT.register\[21\]\[24\] vssd1 vssd1 vccd1 vccd1 net2215 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout837_A _05045_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout458_X net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08678_ net274 _03629_ vssd1 vssd1 vccd1 vccd1 _03798_ sky130_fd_sc_hd__nand2_1
XANTENNA__07143__B1 net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09683__A2 top.a1.instruction\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06497__A2 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07629_ top.DUT.register\[3\]\[5\] net551 net459 top.DUT.register\[17\]\[5\] vssd1
+ vssd1 vccd1 vccd1 _02768_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_37_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10079__X _04955_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08891__B1 net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout625_X net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10640_ net221 net1931 net342 vssd1 vssd1 vccd1 vccd1 _00804_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10571_ net1865 net237 net350 vssd1 vssd1 vccd1 vccd1 _00737_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12310_ _06116_ _06117_ net790 vssd1 vssd1 vccd1 vccd1 _01355_ sky130_fd_sc_hd__and3b_1
XANTENNA__07997__A2 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13290_ clknet_leaf_118_clk _00882_ net933 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[24\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08424__S net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12241_ net2057 _06074_ net978 vssd1 vssd1 vccd1 vccd1 _06076_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_133_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07749__A2 net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08946__B2 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12172_ net1378 net846 net796 _06019_ vssd1 vssd1 vccd1 vccd1 _01280_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_75_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_662 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06957__B1 net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11123_ net53 net867 vssd1 vssd1 vccd1 vccd1 _05067_ sky130_fd_sc_hd__and2_1
XANTENNA_clkbuf_leaf_43_clk_A clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06421__A2 net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_166_2938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11054_ net1214 net865 net837 top.ramstore\[5\] vssd1 vssd1 vccd1 vccd1 _01165_ sky130_fd_sc_hd__a22o_1
XANTENNA__08012__X _03151_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06709__B1 net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10005_ net2178 net168 _04951_ vssd1 vssd1 vccd1 vccd1 _00210_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_199_3426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_199_3437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_58_clk_A clknet_4_12__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_106_2034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_763 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08666__Y _03787_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07134__B1 net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11956_ _05830_ _05838_ vssd1 vssd1 vccd1 vccd1 _05839_ sky130_fd_sc_hd__xnor2_2
XANTENNA__06467__X _01606_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06908__A _02026_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10907_ net2184 net185 net480 vssd1 vssd1 vccd1 vccd1 _01068_ sky130_fd_sc_hd__mux2_1
XFILLER_0_168_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11887_ _05768_ _05769_ _05731_ _05751_ vssd1 vssd1 vccd1 vccd1 _05770_ sky130_fd_sc_hd__a2bb2o_2
XFILLER_0_86_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_156_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09003__B _03902_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11252__C top.lcd.nextState\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10838_ net2144 net197 net475 vssd1 vssd1 vccd1 vccd1 _00999_ sky130_fd_sc_hd__mux2_1
X_13626_ clknet_leaf_75_clk _01213_ net1081 vssd1 vssd1 vccd1 vccd1 net53 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_15_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_116_clk_A clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13557_ clknet_leaf_105_clk _01144_ net968 vssd1 vssd1 vccd1 vccd1 top.ramload\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_10769_ net1352 net232 net482 vssd1 vssd1 vccd1 vccd1 _00930_ sky130_fd_sc_hd__mux2_1
XANTENNA__10864__S net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07988__A2 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12508_ clknet_leaf_78_clk _00100_ net1074 vssd1 vssd1 vccd1 vccd1 top.pc\[20\] sky130_fd_sc_hd__dfrtp_4
X_13488_ clknet_leaf_26_clk _01080_ net1011 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[30\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_12439_ clknet_leaf_87_clk _00035_ net1004 vssd1 vssd1 vccd1 vccd1 top.ramaddr\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_117_2196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08937__A1 net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_196_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06412__A2 net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07980_ top.DUT.register\[18\]\[31\] net548 net517 top.DUT.register\[7\]\[31\] _03118_
+ vssd1 vssd1 vccd1 vccd1 _03119_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_130_2396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07474__A _02590_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06931_ _02069_ vssd1 vssd1 vccd1 vccd1 _02070_ sky130_fd_sc_hd__inv_2
XFILLER_0_38_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08289__B _03421_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09650_ top.a1.halfData\[0\] _01471_ _04683_ _04691_ net1086 vssd1 vssd1 vccd1 vccd1
+ _00115_ sky130_fd_sc_hd__o221a_1
X_06862_ _01996_ _01998_ _02000_ vssd1 vssd1 vccd1 vccd1 _02001_ sky130_fd_sc_hd__or3_1
XANTENNA__10104__S net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07373__B1 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08601_ net886 top.pc\[15\] net697 _03724_ vssd1 vssd1 vccd1 vccd1 _03725_ sky130_fd_sc_hd__a22o_1
X_09581_ top.a1.instruction\[30\] net822 _04470_ vssd1 vssd1 vccd1 vccd1 _04628_ sky130_fd_sc_hd__a21o_2
X_06793_ top.DUT.register\[12\]\[17\] net532 _01931_ vssd1 vssd1 vccd1 vccd1 _01932_
+ sky130_fd_sc_hd__a21o_1
XANTENNA__09114__A1 net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08532_ _02477_ _03658_ vssd1 vssd1 vccd1 vccd1 _03659_ sky130_fd_sc_hd__nor2_1
XANTENNA__07921__B _02567_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08463_ net496 _03592_ _03574_ net423 vssd1 vssd1 vccd1 vccd1 _03593_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_46_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout153_A _04929_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07414_ top.DUT.register\[21\]\[9\] net655 net647 top.DUT.register\[22\]\[9\] _02552_
+ vssd1 vssd1 vccd1 vccd1 _02553_ sky130_fd_sc_hd__a221o_1
XANTENNA__09688__X _04724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08394_ net304 _03398_ _03525_ net286 vssd1 vssd1 vccd1 vccd1 _03526_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_137_2506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07428__A1 _02566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07345_ top.DUT.register\[30\]\[8\] net580 net440 top.DUT.register\[5\]\[8\] _02483_
+ vssd1 vssd1 vccd1 vccd1 _02484_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout320_A _02830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10774__S net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1062_A net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_30_clk clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_30_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout418_A net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07979__A2 net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07276_ top.DUT.register\[17\]\[13\] net749 net637 top.DUT.register\[6\]\[13\] vssd1
+ vssd1 vccd1 vccd1 _02415_ sky130_fd_sc_hd__a22o_1
XFILLER_0_72_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09015_ _03666_ _04083_ _04089_ _03685_ vssd1 vssd1 vccd1 vccd1 _04090_ sky130_fd_sc_hd__or4b_1
X_06227_ top.ramload\[21\] net858 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedInstr\[21\]
+ sky130_fd_sc_hd__and2_1
XANTENNA__12185__B1 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_251 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout206_X net206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold130 top.DUT.register\[26\]\[21\] vssd1 vssd1 vccd1 vccd1 net1246 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold141 top.DUT.register\[17\]\[24\] vssd1 vssd1 vccd1 vccd1 net1257 sky130_fd_sc_hd__dlygate4sd3_1
X_06158_ top.a1.dataIn\[7\] vssd1 vssd1 vccd1 vccd1 _01401_ sky130_fd_sc_hd__inv_2
Xhold152 top.DUT.register\[1\]\[18\] vssd1 vssd1 vccd1 vccd1 net1268 sky130_fd_sc_hd__dlygate4sd3_1
Xhold163 top.ramstore\[23\] vssd1 vssd1 vccd1 vccd1 net1279 sky130_fd_sc_hd__dlygate4sd3_1
Xhold174 top.a1.dataInTemp\[10\] vssd1 vssd1 vccd1 vccd1 net1290 sky130_fd_sc_hd__dlygate4sd3_1
Xhold185 top.edg2.flip1 vssd1 vssd1 vccd1 vccd1 net1301 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09583__B _04628_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout610 _04956_ vssd1 vssd1 vccd1 vccd1 net610 sky130_fd_sc_hd__buf_4
Xhold196 top.DUT.register\[11\]\[17\] vssd1 vssd1 vccd1 vccd1 net1312 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout621 net622 vssd1 vssd1 vccd1 vccd1 net621 sky130_fd_sc_hd__buf_4
XFILLER_0_186_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07384__A _02497_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout632 _04714_ vssd1 vssd1 vccd1 vccd1 net632 sky130_fd_sc_hd__clkbuf_4
X_09917_ _04918_ _04919_ _04911_ vssd1 vssd1 vccd1 vccd1 _04924_ sky130_fd_sc_hd__or3b_1
Xfanout643 _01613_ vssd1 vssd1 vccd1 vccd1 net643 sky130_fd_sc_hd__clkbuf_8
Xfanout654 _01610_ vssd1 vssd1 vccd1 vccd1 net654 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout575_X net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout954_A net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_148_2668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_97_clk clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_97_clk
+ sky130_fd_sc_hd__clkbuf_8
Xfanout665 _01605_ vssd1 vssd1 vccd1 vccd1 net665 sky130_fd_sc_hd__clkbuf_8
Xfanout676 _01548_ vssd1 vssd1 vccd1 vccd1 net676 sky130_fd_sc_hd__buf_2
XANTENNA__10014__S net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout687 _06086_ vssd1 vssd1 vccd1 vccd1 net687 sky130_fd_sc_hd__buf_1
X_09848_ top.pc\[22\] _04514_ _04853_ vssd1 vssd1 vccd1 vccd1 _04861_ sky130_fd_sc_hd__a21o_1
Xfanout698 _01643_ vssd1 vssd1 vccd1 vccd1 net698 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_70_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07364__B1 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10949__S net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout742_X net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_161_2857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09779_ _04798_ _04797_ vssd1 vssd1 vccd1 vccd1 _04799_ sky130_fd_sc_hd__and2b_1
XFILLER_0_198_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_161_2868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11810_ _05661_ _05667_ net131 vssd1 vssd1 vccd1 vccd1 _05693_ sky130_fd_sc_hd__and3b_1
X_12790_ clknet_leaf_12_clk _00382_ net942 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[9\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07116__B1 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11741_ top.a1.dataIn\[9\] _05620_ vssd1 vssd1 vccd1 vccd1 _05624_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07667__A1 top.a1.instruction\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_194_3356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06447__B _01585_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09598__X _04644_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11672_ top.a1.dataIn\[11\] _05525_ _05549_ vssd1 vssd1 vccd1 vccd1 _05555_ sky130_fd_sc_hd__or3b_1
XANTENNA__08943__A net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_518 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10623_ net159 net2110 net349 vssd1 vssd1 vccd1 vccd1 _00788_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13411_ clknet_leaf_54_clk _01003_ net1037 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[28\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_12_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10684__S net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06890__A2 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_21_clk clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_21_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_91_460 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13342_ clknet_leaf_55_clk _00934_ net1032 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[26\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_64_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10554_ net1427 net172 net355 vssd1 vssd1 vccd1 vccd1 _00721_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06642__A2 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13273_ clknet_leaf_14_clk _00865_ net959 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[24\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_10485_ net1495 net183 net362 vssd1 vssd1 vccd1 vccd1 _00655_ sky130_fd_sc_hd__mux2_1
X_12224_ _06059_ _06065_ net980 vssd1 vssd1 vccd1 vccd1 _01315_ sky130_fd_sc_hd__o21a_1
XFILLER_0_20_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12155_ _06006_ _06034_ _06028_ vssd1 vssd1 vccd1 vccd1 _06038_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_209_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06910__B _02048_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11106_ net907 top.ramaddr\[12\] net861 _05058_ vssd1 vssd1 vccd1 vccd1 _01204_ sky130_fd_sc_hd__a31o_1
XANTENNA__07294__A _02409_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12873__RESET_B net1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12086_ _05951_ _05968_ vssd1 vssd1 vccd1 vccd1 _05969_ sky130_fd_sc_hd__nor2_1
XFILLER_0_75_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_88_clk clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_88_clk
+ sky130_fd_sc_hd__clkbuf_8
X_11037_ net17 net838 net816 top.ramload\[23\] vssd1 vssd1 vccd1 vccd1 _01149_ sky130_fd_sc_hd__o22a_1
XANTENNA__07355__B1 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08552__C1 net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10859__S net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_182_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06197__X _01428_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07107__B1 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12988_ clknet_leaf_2_clk _00580_ net914 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[15\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11939_ net128 _05818_ _05820_ _05783_ vssd1 vssd1 vccd1 vccd1 _05822_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_87_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08853__A _01790_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13609_ clknet_leaf_73_clk _01196_ net1078 vssd1 vssd1 vccd1 vccd1 net66 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_119_2225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10594__S net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_184_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_2236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06881__A2 net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_12_clk clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_12_clk
+ sky130_fd_sc_hd__clkbuf_8
X_07130_ top.DUT.register\[30\]\[11\] net579 net463 top.DUT.register\[13\]\[11\] _02268_
+ vssd1 vssd1 vccd1 vccd1 _02269_ sky130_fd_sc_hd__a221o_1
XFILLER_0_40_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07061_ top.DUT.register\[20\]\[22\] net664 net771 top.DUT.register\[10\]\[22\] vssd1
+ vssd1 vccd1 vccd1 _02200_ sky130_fd_sc_hd__a22o_1
XANTENNA__06633__A2 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_2425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_152_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09684__A _04712_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10182__X _04962_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07594__B1 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_276 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07963_ _01572_ _01656_ _03101_ vssd1 vssd1 vccd1 vccd1 _03102_ sky130_fd_sc_hd__a21boi_1
Xclkbuf_leaf_79_clk clknet_4_12__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_79_clk
+ sky130_fd_sc_hd__clkbuf_8
X_06914_ top.DUT.register\[28\]\[21\] net557 net518 top.DUT.register\[7\]\[21\] vssd1
+ vssd1 vccd1 vccd1 _02053_ sky130_fd_sc_hd__a22o_1
XFILLER_0_4_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09702_ net828 _04223_ vssd1 vssd1 vccd1 vccd1 _04734_ sky130_fd_sc_hd__nor2_1
X_07894_ top.DUT.register\[14\]\[1\] net585 net446 top.DUT.register\[1\]\[1\] vssd1
+ vssd1 vccd1 vccd1 _03033_ sky130_fd_sc_hd__a22o_1
XANTENNA__07346__B1 net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11142__A1 net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06845_ top.DUT.register\[16\]\[19\] net735 net712 top.DUT.register\[11\]\[19\] vssd1
+ vssd1 vccd1 vccd1 _01984_ sky130_fd_sc_hd__a22o_1
X_09633_ top.pad.keyCode\[4\] top.pad.keyCode\[6\] top.pad.keyCode\[7\] top.pad.keyCode\[5\]
+ vssd1 vssd1 vccd1 vccd1 _04675_ sky130_fd_sc_hd__or4b_2
XANTENNA__10769__S net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout270_A _04726_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09564_ _04204_ _04612_ top.pc\[28\] _04051_ vssd1 vssd1 vccd1 vccd1 _00108_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_143_2587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06776_ _01910_ _01912_ _01914_ vssd1 vssd1 vccd1 vccd1 _01915_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_143_2598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08515_ _02476_ _03641_ vssd1 vssd1 vccd1 vccd1 _03642_ sky130_fd_sc_hd__xnor2_1
X_09495_ _04529_ _04547_ _04546_ vssd1 vssd1 vccd1 vccd1 _04548_ sky130_fd_sc_hd__a21o_1
XFILLER_0_194_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout535_A _01541_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06267__B net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout156_X net156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08446_ _03540_ _03575_ net293 vssd1 vssd1 vccd1 vccd1 _03576_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_176_3086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06872__A2 net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08377_ _02754_ _03509_ vssd1 vssd1 vccd1 vccd1 _03510_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_190_432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout702_A _01642_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_471 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07328_ top.DUT.register\[10\]\[12\] net770 net722 top.DUT.register\[29\]\[12\] vssd1
+ vssd1 vccd1 vccd1 _02467_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_12_Left_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_178 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_59_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07259_ top.DUT.register\[7\]\[13\] net517 net441 top.DUT.register\[5\]\[13\] _02397_
+ vssd1 vssd1 vccd1 vccd1 _02398_ sky130_fd_sc_hd__a221o_1
XANTENNA__10009__S net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10270_ net2048 net245 net385 vssd1 vssd1 vccd1 vccd1 _00448_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout692_X net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_72_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06388__A1 top.a1.instruction\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout440 _01566_ vssd1 vssd1 vccd1 vccd1 net440 sky130_fd_sc_hd__clkbuf_4
Xfanout451 _01561_ vssd1 vssd1 vccd1 vccd1 net451 sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_21_Left_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout462 _01552_ vssd1 vssd1 vccd1 vccd1 net462 sky130_fd_sc_hd__buf_4
Xfanout473 _05098_ vssd1 vssd1 vccd1 vccd1 net473 sky130_fd_sc_hd__buf_2
Xfanout484 _04962_ vssd1 vssd1 vccd1 vccd1 net484 sky130_fd_sc_hd__buf_6
Xfanout495 _03338_ vssd1 vssd1 vccd1 vccd1 net495 sky130_fd_sc_hd__buf_2
X_12911_ clknet_leaf_41_clk _00503_ net1045 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[12\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10679__S net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_543 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12842_ clknet_leaf_118_clk _00434_ net953 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[10\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_198_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_232 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11083__B net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12773_ clknet_leaf_34_clk _00365_ net1040 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[8\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_96_574 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10644__A0 net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_185_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11724_ _05540_ _05572_ vssd1 vssd1 vccd1 vccd1 _05607_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_83_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_30_Left_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11655_ _05507_ _05510_ _05515_ vssd1 vssd1 vccd1 vccd1 _05538_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_193_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10606_ net229 net2053 net346 vssd1 vssd1 vccd1 vccd1 _00771_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11586_ _05410_ _05464_ _05465_ _05467_ vssd1 vssd1 vccd1 vccd1 _05469_ sky130_fd_sc_hd__nor4b_1
XFILLER_0_107_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13325_ clknet_leaf_42_clk _00917_ net1064 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[25\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_10537_ net1907 net246 net354 vssd1 vssd1 vccd1 vccd1 _00704_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_143 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_2155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10468_ net1926 net252 net361 vssd1 vssd1 vccd1 vccd1 _00638_ sky130_fd_sc_hd__mux2_1
X_13256_ clknet_leaf_8_clk _00848_ net947 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[23\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_12207_ top.lcd.cnt_20ms\[5\] _06052_ vssd1 vssd1 vccd1 vccd1 _06053_ sky130_fd_sc_hd__and2_1
X_13187_ clknet_leaf_57_clk _00779_ net1076 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[21\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_10399_ net1306 net266 _04982_ vssd1 vssd1 vccd1 vccd1 _00571_ sky130_fd_sc_hd__mux2_1
X_12138_ _06017_ _06018_ vssd1 vssd1 vccd1 vccd1 _06021_ sky130_fd_sc_hd__nand2_1
XANTENNA__09009__A net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12069_ _05930_ _05935_ _05937_ vssd1 vssd1 vccd1 vccd1 _05952_ sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_1_clk clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_1_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__11124__A1 net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07328__B1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09868__A2 _04543_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10589__S net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06630_ top.DUT.register\[30\]\[27\] net761 net716 top.DUT.register\[27\]\[27\] _01768_
+ vssd1 vssd1 vccd1 vccd1 _01769_ sky130_fd_sc_hd__a221o_1
XFILLER_0_177_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06561_ _01678_ _01698_ vssd1 vssd1 vccd1 vccd1 _01700_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_714 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08300_ net305 _03254_ vssd1 vssd1 vccd1 vccd1 _03435_ sky130_fd_sc_hd__nand2_1
XFILLER_0_176_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_192_708 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09280_ top.pc\[12\] _04326_ vssd1 vssd1 vccd1 vccd1 _04345_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_47_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06492_ top.DUT.register\[7\]\[30\] net660 net637 top.DUT.register\[6\]\[30\] vssd1
+ vssd1 vccd1 vccd1 _01631_ sky130_fd_sc_hd__a22o_1
XFILLER_0_47_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07500__B1 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_602 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08231_ _03191_ _03199_ net293 vssd1 vssd1 vccd1 vccd1 _03368_ sky130_fd_sc_hd__mux2_1
XANTENNA__06854__A2 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08162_ _01897_ net329 vssd1 vssd1 vccd1 vccd1 _03300_ sky130_fd_sc_hd__nand2_1
XFILLER_0_83_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_498 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07113_ top.DUT.register\[13\]\[16\] net775 net731 top.DUT.register\[14\]\[16\] vssd1
+ vssd1 vccd1 vccd1 _02252_ sky130_fd_sc_hd__a22o_1
XANTENNA__11060__B1 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08093_ _03230_ _03231_ vssd1 vssd1 vccd1 vccd1 _03232_ sky130_fd_sc_hd__and2_1
XFILLER_0_141_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload50 clknet_leaf_84_clk vssd1 vssd1 vccd1 vccd1 clkload50/Y sky130_fd_sc_hd__inv_12
XFILLER_0_30_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07044_ top.DUT.register\[22\]\[22\] net575 net552 top.DUT.register\[3\]\[22\] _02182_
+ vssd1 vssd1 vccd1 vccd1 _02183_ sky130_fd_sc_hd__a221o_1
XFILLER_0_113_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkload61 clknet_leaf_25_clk vssd1 vssd1 vccd1 vccd1 clkload61/X sky130_fd_sc_hd__clkbuf_8
Xclkload72 clknet_leaf_32_clk vssd1 vssd1 vccd1 vccd1 clkload72/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_2_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload83 clknet_leaf_45_clk vssd1 vssd1 vccd1 vccd1 clkload83/Y sky130_fd_sc_hd__inv_6
XFILLER_0_23_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload94 clknet_leaf_71_clk vssd1 vssd1 vccd1 vccd1 clkload94/Y sky130_fd_sc_hd__inv_8
XANTENNA__07567__B1 net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1025_A net1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07031__A2 net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08995_ _03999_ _04020_ _04038_ vssd1 vssd1 vccd1 vccd1 _04070_ sky130_fd_sc_hd__or3_1
XANTENNA_fanout485_A _04962_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09308__A1 _02399_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_2616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07946_ _03083_ _03084_ _02222_ vssd1 vssd1 vccd1 vccd1 _03085_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_145_2627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07319__B1 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07662__A _02773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07877_ top.DUT.register\[5\]\[1\] net653 net641 top.DUT.register\[8\]\[1\] vssd1
+ vssd1 vccd1 vccd1 _03016_ sky130_fd_sc_hd__a22o_1
XANTENNA__10499__S net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout652_A _01610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09616_ _04660_ vssd1 vssd1 vccd1 vccd1 _04661_ sky130_fd_sc_hd__inv_2
X_06828_ top.DUT.register\[9\]\[19\] net469 net549 top.DUT.register\[18\]\[19\] vssd1
+ vssd1 vccd1 vccd1 _01967_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_178_3115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_195_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_738 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06759_ top.DUT.register\[18\]\[24\] net729 net638 top.DUT.register\[6\]\[24\] vssd1
+ vssd1 vccd1 vccd1 _01898_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout440_X net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09547_ net902 top.pc\[27\] _04595_ _04596_ net890 vssd1 vssd1 vccd1 vccd1 _00107_
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_167_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout917_A net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout538_X net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_191_3304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_183_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_191_3315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08295__A1 net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07098__A2 net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08295__B2 _03430_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09478_ _04528_ _04531_ vssd1 vssd1 vccd1 vccd1 _04532_ sky130_fd_sc_hd__xor2_1
XFILLER_0_148_462 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08429_ net325 _03559_ _03558_ vssd1 vssd1 vccd1 vccd1 _03560_ sky130_fd_sc_hd__o21a_2
XANTENNA__06845__A2 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout705_X net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10528__A _04712_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11440_ _05286_ _05320_ _05322_ vssd1 vssd1 vccd1 vccd1 _05323_ sky130_fd_sc_hd__and3_1
Xclkload0 clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clkload0/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_151_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_156_2789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_22_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_655 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11051__B1 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09795__A1 _03765_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11371_ _05252_ _05253_ vssd1 vssd1 vccd1 vccd1 _05254_ sky130_fd_sc_hd__or2_1
X_10322_ net166 net2282 net383 vssd1 vssd1 vccd1 vccd1 _00499_ sky130_fd_sc_hd__mux2_1
X_13110_ clknet_leaf_4_clk _00702_ net942 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[19\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_189_3277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_189_3288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13041_ clknet_leaf_115_clk _00633_ net963 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[17\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_10253_ net178 net2164 net390 vssd1 vssd1 vccd1 vccd1 _00432_ sky130_fd_sc_hd__mux2_1
XANTENNA__07558__B1 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07022__A2 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10184_ _04963_ vssd1 vssd1 vccd1 vccd1 _04964_ sky130_fd_sc_hd__clkinv_4
XTAP_TAPCELL_ROW_208_3561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_208_3572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout270 _04726_ vssd1 vssd1 vccd1 vccd1 net270 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout281 net282 vssd1 vssd1 vccd1 vccd1 net281 sky130_fd_sc_hd__buf_2
Xfanout292 net294 vssd1 vssd1 vccd1 vccd1 net292 sky130_fd_sc_hd__buf_2
XFILLER_0_199_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09180__C1 net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10202__S net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07730__B1 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12825_ clknet_leaf_11_clk _00417_ net948 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[10\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07089__A2 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09499__A top.pc\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06475__X _01614_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12756_ clknet_leaf_56_clk _00348_ net1075 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[8\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11707_ _05553_ _05581_ _05561_ vssd1 vssd1 vccd1 vccd1 _05590_ sky130_fd_sc_hd__a21boi_1
XANTENNA__11290__B1 _05136_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06836__A2 net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12687_ clknet_leaf_22_clk _00279_ net1024 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[5\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_11638_ _05514_ _05515_ _05506_ vssd1 vssd1 vccd1 vccd1 _05521_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_112_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_142_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08589__A2 net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10872__S net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11569_ _05448_ _05449_ _05451_ top.a1.dataIn\[13\] vssd1 vssd1 vccd1 vccd1 _05452_
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_97_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold707 top.DUT.register\[16\]\[1\] vssd1 vssd1 vccd1 vccd1 net1823 sky130_fd_sc_hd__dlygate4sd3_1
Xhold718 top.DUT.register\[16\]\[26\] vssd1 vssd1 vccd1 vccd1 net1834 sky130_fd_sc_hd__dlygate4sd3_1
X_13308_ clknet_leaf_2_clk _00900_ net915 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[25\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold729 top.DUT.register\[5\]\[14\] vssd1 vssd1 vccd1 vccd1 net1845 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07261__A2 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13239_ clknet_leaf_129_clk _00831_ net912 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[23\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06370__B net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07549__B1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07013__A2 net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07800_ top.DUT.register\[30\]\[2\] net579 net563 top.DUT.register\[20\]\[2\] vssd1
+ vssd1 vccd1 vccd1 _02939_ sky130_fd_sc_hd__a22o_1
X_08780_ _01920_ _03893_ vssd1 vssd1 vccd1 vccd1 _03895_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_127_Right_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_2346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07731_ top.DUT.register\[9\]\[3\] net763 net728 top.DUT.register\[18\]\[3\] _02859_
+ vssd1 vssd1 vccd1 vccd1 _02870_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_127_2357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10856__A0 net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09710__A1 _03488_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07662_ _02773_ _02798_ vssd1 vssd1 vccd1 vccd1 _02801_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_0_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07721__B1 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06613_ top.DUT.register\[9\]\[27\] net469 net549 top.DUT.register\[18\]\[27\] vssd1
+ vssd1 vccd1 vccd1 _01752_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_0_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09401_ net137 _04446_ _04459_ vssd1 vssd1 vccd1 vccd1 _04460_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_140_2546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_189_395 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07593_ top.DUT.register\[25\]\[6\] net778 net750 top.DUT.register\[26\]\[6\] vssd1
+ vssd1 vccd1 vccd1 _02732_ sky130_fd_sc_hd__a22o_1
XANTENNA__08584__Y _03708_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06544_ top.DUT.register\[10\]\[29\] net772 net637 top.DUT.register\[6\]\[29\] _01682_
+ vssd1 vssd1 vccd1 vccd1 _01683_ sky130_fd_sc_hd__a221o_1
X_09332_ net897 top.pc\[14\] _04394_ net889 vssd1 vssd1 vccd1 vccd1 _00094_ sky130_fd_sc_hd__o211a_1
XFILLER_0_75_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_173_3034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09263_ _02365_ top.pc\[11\] vssd1 vssd1 vccd1 vccd1 _04329_ sky130_fd_sc_hd__and2b_1
XANTENNA__09202__A top.pc\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06827__A2 net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_173_3045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06475_ net787 _01600_ _01611_ vssd1 vssd1 vccd1 vccd1 _01614_ sky130_fd_sc_hd__and3_4
XFILLER_0_173_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13720__Q top.a1.row2\[34\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout233_A _04760_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08214_ _03045_ _03340_ net425 net426 _03330_ vssd1 vssd1 vccd1 vccd1 _03352_ sky130_fd_sc_hd__a32o_1
XFILLER_0_16_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_238 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09194_ _04246_ _04263_ _04264_ vssd1 vssd1 vccd1 vccd1 _04265_ sky130_fd_sc_hd__nand3_1
XFILLER_0_173_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08145_ _03279_ _03282_ net293 vssd1 vssd1 vccd1 vccd1 _03283_ sky130_fd_sc_hd__mux2_1
XANTENNA__10782__S net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07788__B1 net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08076_ _01983_ net300 vssd1 vssd1 vccd1 vccd1 _03215_ sky130_fd_sc_hd__or2_1
XANTENNA__07252__A2 net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06561__A _01678_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07027_ top.DUT.register\[15\]\[20\] net709 net701 top.DUT.register\[31\]\[20\] vssd1
+ vssd1 vccd1 vccd1 _02166_ sky130_fd_sc_hd__a22o_1
XFILLER_0_30_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07004__A2 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout390_X net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout488_X net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout867_A net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold12 top.ru.state\[1\] vssd1 vssd1 vccd1 vccd1 net1128 sky130_fd_sc_hd__dlygate4sd3_1
Xhold23 top.ramstore\[17\] vssd1 vssd1 vccd1 vccd1 net1139 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09591__B _04620_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold34 _01191_ vssd1 vssd1 vccd1 vccd1 net1150 sky130_fd_sc_hd__dlygate4sd3_1
X_08978_ _04052_ _03487_ _03446_ _03423_ vssd1 vssd1 vccd1 vccd1 _04053_ sky130_fd_sc_hd__and4b_1
Xhold45 top.a1.row1\[104\] vssd1 vssd1 vccd1 vccd1 net1161 sky130_fd_sc_hd__dlygate4sd3_1
Xhold56 top.a1.data\[8\] vssd1 vssd1 vccd1 vccd1 net1172 sky130_fd_sc_hd__dlygate4sd3_1
Xhold67 _01183_ vssd1 vssd1 vccd1 vccd1 net1183 sky130_fd_sc_hd__dlygate4sd3_1
Xhold78 _01170_ vssd1 vssd1 vccd1 vccd1 net1194 sky130_fd_sc_hd__dlygate4sd3_1
X_07929_ _02390_ _03062_ _03067_ vssd1 vssd1 vccd1 vccd1 _03068_ sky130_fd_sc_hd__o21a_1
XANTENNA__08827__A1_N net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold89 top.ramstore\[16\] vssd1 vssd1 vccd1 vccd1 net1205 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout655_X net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10940_ net1566 net202 net592 vssd1 vssd1 vccd1 vccd1 _01101_ sky130_fd_sc_hd__mux2_1
XANTENNA__10022__S net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_196_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_203_3491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10871_ net189 net1906 net595 vssd1 vssd1 vccd1 vccd1 _01032_ sky130_fd_sc_hd__mux2_1
XFILLER_0_210_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12610_ clknet_leaf_11_clk _00202_ net948 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[3\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_211_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_158_2818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13590_ clknet_leaf_46_clk net1140 net1066 vssd1 vssd1 vccd1 vccd1 net81 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_183_527 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12541_ clknet_leaf_3_clk _00133_ net941 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[1\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06818__A2 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_164_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_6__f_clk_X clknet_4_6__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12472_ clknet_leaf_46_clk _00067_ net1066 vssd1 vssd1 vccd1 vccd1 top.ramstore\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07491__A2 net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09768__A1 top.pc\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11423_ _05291_ _05298_ _05303_ _05304_ _05302_ vssd1 vssd1 vccd1 vccd1 _05306_ sky130_fd_sc_hd__a221oi_4
XANTENNA__10692__S net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07779__B1 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_9 _03868_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11354_ _05224_ _05226_ _05235_ vssd1 vssd1 vccd1 vccd1 _05237_ sky130_fd_sc_hd__a21o_1
XANTENNA__07243__A2 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_111_2114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10305_ net231 net2047 net381 vssd1 vssd1 vccd1 vccd1 _00482_ sky130_fd_sc_hd__mux2_1
XANTENNA__06451__B1 _01589_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11285_ top.a1.row1\[59\] _05136_ _05143_ top.a1.row2\[3\] _05174_ vssd1 vssd1 vccd1
+ vccd1 _05175_ sky130_fd_sc_hd__a221o_1
XANTENNA__07854__X _02993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10236_ net243 net1754 net389 vssd1 vssd1 vccd1 vccd1 _00415_ sky130_fd_sc_hd__mux2_1
X_13024_ clknet_leaf_55_clk _00616_ net1031 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[16\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1010 net1011 vssd1 vssd1 vccd1 vccd1 net1010 sky130_fd_sc_hd__clkbuf_4
Xfanout1021 net1025 vssd1 vssd1 vccd1 vccd1 net1021 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09940__A1 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10167_ net1521 net192 net605 vssd1 vssd1 vccd1 vccd1 _00366_ sky130_fd_sc_hd__mux2_1
Xfanout1032 net1039 vssd1 vssd1 vccd1 vccd1 net1032 sky130_fd_sc_hd__clkbuf_2
Xfanout1043 net1048 vssd1 vssd1 vccd1 vccd1 net1043 sky130_fd_sc_hd__clkbuf_2
Xfanout1054 net1055 vssd1 vssd1 vccd1 vccd1 net1054 sky130_fd_sc_hd__clkbuf_4
Xfanout1065 net1068 vssd1 vssd1 vccd1 vccd1 net1065 sky130_fd_sc_hd__clkbuf_4
Xfanout1076 net1087 vssd1 vssd1 vccd1 vccd1 net1076 sky130_fd_sc_hd__clkbuf_4
X_10098_ net1714 net205 net613 vssd1 vssd1 vccd1 vccd1 _00299_ sky130_fd_sc_hd__mux2_1
Xfanout1087 net1098 vssd1 vssd1 vccd1 vccd1 net1087 sky130_fd_sc_hd__clkbuf_4
Xfanout1098 net39 vssd1 vssd1 vccd1 vccd1 net1098 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_109_2076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_2087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_199_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07703__B1 net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_682 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09721__S net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10867__S net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_202_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_122_2276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12808_ clknet_leaf_27_clk _00400_ net1008 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[9\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13788_ clknet_leaf_68_clk _01357_ vssd1 vssd1 vccd1 vccd1 top.pad.button_control.r_counter\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__06809__A2 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12739_ clknet_leaf_58_clk _00331_ net1088 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[7\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_139_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_216 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_0_clk_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_98_1909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06260_ top.ramload\[21\] net853 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedData\[21\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_199_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07482__A2 net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_170_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11015__B1 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09759__B2 top.a1.dataIn\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06191_ _01420_ _01426_ vssd1 vssd1 vccd1 vccd1 top.a1.nextHex\[3\] sky130_fd_sc_hd__or2_1
XFILLER_0_170_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_142_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold504 top.DUT.register\[4\]\[13\] vssd1 vssd1 vccd1 vccd1 net1620 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_170_799 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07234__A2 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold515 top.ramaddr\[8\] vssd1 vssd1 vccd1 vccd1 net1631 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08431__B2 net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold526 top.DUT.register\[30\]\[31\] vssd1 vssd1 vccd1 vccd1 net1642 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold537 top.DUT.register\[5\]\[13\] vssd1 vssd1 vccd1 vccd1 net1653 sky130_fd_sc_hd__dlygate4sd3_1
Xhold548 top.DUT.register\[27\]\[31\] vssd1 vssd1 vccd1 vccd1 net1664 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13292__CLK clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09950_ net1372 net253 net627 vssd1 vssd1 vccd1 vccd1 _00158_ sky130_fd_sc_hd__mux2_1
Xhold559 top.DUT.register\[21\]\[31\] vssd1 vssd1 vccd1 vccd1 net1675 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10107__S net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xmax_cap278 _05324_ vssd1 vssd1 vccd1 vccd1 net278 sky130_fd_sc_hd__clkbuf_2
XANTENNA__06993__A1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08901_ _04009_ _04010_ vssd1 vssd1 vccd1 vccd1 _04011_ sky130_fd_sc_hd__nand2_1
X_09881_ _04889_ _04890_ vssd1 vssd1 vccd1 vccd1 _04891_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_148_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_51_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09931__A1 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08832_ net281 _03372_ vssd1 vssd1 vccd1 vccd1 _03945_ sky130_fd_sc_hd__nor2_1
X_08763_ _03534_ _03542_ _03716_ net279 _03878_ vssd1 vssd1 vccd1 vccd1 _03879_ sky130_fd_sc_hd__o221a_1
XANTENNA__08101__A _02633_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout183_A _04858_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07714_ top.a1.instruction\[10\] _01474_ vssd1 vssd1 vccd1 vccd1 _02853_ sky130_fd_sc_hd__and2_1
XANTENNA__08498__A1 net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08694_ _02050_ _03761_ _03079_ vssd1 vssd1 vccd1 vccd1 _03813_ sky130_fd_sc_hd__o21ai_1
XANTENNA__09695__B1 net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07645_ top.DUT.register\[14\]\[5\] net730 net722 top.DUT.register\[29\]\[5\] vssd1
+ vssd1 vccd1 vccd1 _02784_ sky130_fd_sc_hd__a22o_1
XANTENNA__10777__S net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout350_A net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1092_A net1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout448_A _01562_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07576_ top.DUT.register\[30\]\[6\] net579 _02714_ vssd1 vssd1 vccd1 vccd1 _02715_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_48_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_165_538 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10057__A1 net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06527_ top.DUT.register\[22\]\[29\] net577 net528 top.DUT.register\[26\]\[29\] vssd1
+ vssd1 vccd1 vccd1 _01666_ sky130_fd_sc_hd__a22o_1
X_09315_ top.pc\[14\] _04360_ vssd1 vssd1 vccd1 vccd1 _04378_ sky130_fd_sc_hd__nor2_1
XFILLER_0_63_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout615_A _04954_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_192_379 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06458_ _01591_ _01594_ _01596_ vssd1 vssd1 vccd1 vccd1 _01597_ sky130_fd_sc_hd__and3_2
X_09246_ _04298_ _04301_ _04299_ vssd1 vssd1 vccd1 vccd1 _04313_ sky130_fd_sc_hd__a21o_1
XFILLER_0_8_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_153_2737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09813__B1_N _04829_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06681__B1 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_153_2748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09177_ _04245_ _04248_ net812 vssd1 vssd1 vccd1 vccd1 _04249_ sky130_fd_sc_hd__a21oi_1
X_06389_ net684 _01516_ _01527_ vssd1 vssd1 vccd1 vccd1 _01528_ sky130_fd_sc_hd__and3_4
XANTENNA_fanout403_X net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08128_ top.ru.state\[0\] _01481_ vssd1 vssd1 vccd1 vccd1 _03267_ sky130_fd_sc_hd__nand2_1
XFILLER_0_121_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08751__A1_N net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08059_ _01810_ net328 vssd1 vssd1 vccd1 vccd1 _03198_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_186_3236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10017__S net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput46 net46 vssd1 vssd1 vccd1 vccd1 ADR_O[15] sky130_fd_sc_hd__buf_2
XANTENNA__09806__S net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11070_ net86 net870 net834 net1152 vssd1 vssd1 vccd1 vccd1 _01181_ sky130_fd_sc_hd__a22o_1
Xoutput57 net57 vssd1 vssd1 vccd1 vccd1 ADR_O[25] sky130_fd_sc_hd__buf_2
Xoutput68 net68 vssd1 vssd1 vccd1 vccd1 ADR_O[6] sky130_fd_sc_hd__buf_2
Xoutput79 net79 vssd1 vssd1 vccd1 vccd1 DAT_O[15] sky130_fd_sc_hd__buf_2
XANTENNA_fanout772_X net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10021_ net1220 net248 net619 vssd1 vssd1 vccd1 vccd1 _00224_ sky130_fd_sc_hd__mux2_1
XANTENNA__09383__C1 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_205_3520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_203_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_164_2899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08489__A1 net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_811 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11972_ _05847_ _05849_ _05841_ vssd1 vssd1 vccd1 vccd1 _05855_ sky130_fd_sc_hd__a21boi_1
XANTENNA__08489__B2 _03617_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11088__A3 net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_455 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_2_clk_A clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13711_ clknet_leaf_96_clk _01282_ net984 vssd1 vssd1 vccd1 vccd1 top.a1.row2\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_168_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10923_ net1503 net259 net591 vssd1 vssd1 vccd1 vccd1 _01084_ sky130_fd_sc_hd__mux2_1
XANTENNA__10687__S net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_19_Right_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11372__A top.a1.dataIn\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_197_3398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13642_ clknet_leaf_94_clk _00006_ net982 vssd1 vssd1 vccd1 vccd1 top.ru.state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_156_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10854_ net1832 net148 net475 vssd1 vssd1 vccd1 vccd1 _01015_ sky130_fd_sc_hd__mux2_1
XFILLER_0_183_313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_4_Left_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13573_ clknet_leaf_66_clk net1243 net1094 vssd1 vssd1 vccd1 vccd1 net73 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_66_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10785_ net1699 net169 net482 vssd1 vssd1 vccd1 vccd1 _00946_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12524_ clknet_leaf_71_clk _00116_ vssd1 vssd1 vccd1 vccd1 top.a1.halfData\[1\] sky130_fd_sc_hd__dfxtp_2
XANTENNA__08661__A1 _03264_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07464__A2 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08661__B2 _03169_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06672__B1 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12455_ clknet_leaf_66_clk _00050_ net1094 vssd1 vssd1 vccd1 vccd1 top.ramstore\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_191_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11406_ _05220_ _05255_ vssd1 vssd1 vccd1 vccd1 _05289_ sky130_fd_sc_hd__or2_1
XFILLER_0_151_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08413__A1 net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12386_ clknet_leaf_110_clk top.ru.next_FetchedData\[30\] net977 vssd1 vssd1 vccd1
+ vccd1 top.a1.dataIn\[30\] sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_28_Right_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_1839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06424__B1 net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12353__D net1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11337_ top.a1.dataIn\[20\] _05218_ vssd1 vssd1 vccd1 vccd1 _05220_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_120_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09716__S net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09943__C _04708_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11268_ top.a1.row1\[9\] _05126_ _05140_ top.a1.row2\[33\] _05159_ vssd1 vssd1 vccd1
+ vccd1 _05160_ sky130_fd_sc_hd__a221o_1
XFILLER_0_94_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13007_ clknet_leaf_51_clk _00599_ net1056 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[15\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_10219_ net182 net2235 net396 vssd1 vssd1 vccd1 vccd1 _00399_ sky130_fd_sc_hd__mux2_1
X_11199_ net845 _05007_ _05021_ vssd1 vssd1 vccd1 vccd1 _05106_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_124_2305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_168_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_37_Right_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_wire416_A net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10597__S net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07430_ _02544_ _02567_ vssd1 vssd1 vccd1 vccd1 _02569_ sky130_fd_sc_hd__nor2_1
XFILLER_0_147_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06360__C1 net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07361_ _02330_ net410 net794 vssd1 vssd1 vccd1 vccd1 _02500_ sky130_fd_sc_hd__a21o_1
XFILLER_0_128_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09100_ _02357_ _04149_ _04172_ vssd1 vssd1 vccd1 vccd1 _04175_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_102_1979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06312_ _01451_ _01453_ _01456_ _01448_ vssd1 vssd1 vccd1 vccd1 _01467_ sky130_fd_sc_hd__o31a_1
XANTENNA__07455__A2 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07292_ _02409_ _02430_ vssd1 vssd1 vccd1 vccd1 _02431_ sky130_fd_sc_hd__nand2_2
XFILLER_0_17_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09031_ _03657_ _03699_ _03726_ _03767_ vssd1 vssd1 vccd1 vccd1 _04106_ sky130_fd_sc_hd__or4b_1
XANTENNA__06663__B1 net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06243_ net1224 net854 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedData\[4\] sky130_fd_sc_hd__and2_1
XANTENNA__10185__X _04965_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_46_Right_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_135_2467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_2478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06174_ _01413_ _01415_ vssd1 vssd1 vccd1 vccd1 _01416_ sky130_fd_sc_hd__and2_1
Xhold301 top.DUT.register\[15\]\[21\] vssd1 vssd1 vccd1 vccd1 net1417 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold312 top.DUT.register\[19\]\[31\] vssd1 vssd1 vccd1 vccd1 net1428 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_287 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold323 top.DUT.register\[20\]\[15\] vssd1 vssd1 vccd1 vccd1 net1439 sky130_fd_sc_hd__dlygate4sd3_1
Xhold334 top.DUT.register\[15\]\[16\] vssd1 vssd1 vccd1 vccd1 net1450 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08955__A2 net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold345 top.DUT.register\[12\]\[0\] vssd1 vssd1 vccd1 vccd1 net1461 sky130_fd_sc_hd__dlygate4sd3_1
Xhold356 top.DUT.register\[11\]\[12\] vssd1 vssd1 vccd1 vccd1 net1472 sky130_fd_sc_hd__dlygate4sd3_1
Xhold367 top.DUT.register\[14\]\[22\] vssd1 vssd1 vccd1 vccd1 net1483 sky130_fd_sc_hd__dlygate4sd3_1
Xhold378 top.DUT.register\[27\]\[25\] vssd1 vssd1 vccd1 vccd1 net1494 sky130_fd_sc_hd__dlygate4sd3_1
Xhold389 top.DUT.register\[2\]\[24\] vssd1 vssd1 vccd1 vccd1 net1505 sky130_fd_sc_hd__dlygate4sd3_1
X_09933_ net1871 net150 net633 vssd1 vssd1 vccd1 vccd1 _00151_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout803 _03269_ vssd1 vssd1 vccd1 vccd1 net803 sky130_fd_sc_hd__buf_2
XFILLER_0_111_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout814 _01446_ vssd1 vssd1 vccd1 vccd1 net814 sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_209_Left_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout825 _01575_ vssd1 vssd1 vccd1 vccd1 net825 sky130_fd_sc_hd__buf_4
XANTENNA__08707__A2 net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09365__C1 net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout836 net837 vssd1 vssd1 vccd1 vccd1 net836 sky130_fd_sc_hd__buf_2
Xfanout847 net848 vssd1 vssd1 vccd1 vccd1 net847 sky130_fd_sc_hd__buf_2
X_09864_ _03909_ net404 net489 _04875_ vssd1 vssd1 vccd1 vccd1 _04876_ sky130_fd_sc_hd__o211a_2
Xfanout858 net859 vssd1 vssd1 vccd1 vccd1 net858 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_181_3155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1001 top.DUT.register\[13\]\[0\] vssd1 vssd1 vccd1 vccd1 net2117 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout869 _01427_ vssd1 vssd1 vccd1 vccd1 net869 sky130_fd_sc_hd__clkbuf_2
Xhold1012 top.DUT.register\[17\]\[16\] vssd1 vssd1 vccd1 vccd1 net2128 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_181_3166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08815_ net424 _03928_ _03926_ _03914_ vssd1 vssd1 vccd1 vccd1 _03929_ sky130_fd_sc_hd__a211o_2
XANTENNA__09380__A2 _01939_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1023 top.DUT.register\[1\]\[10\] vssd1 vssd1 vccd1 vccd1 net2139 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1034 top.DUT.register\[22\]\[19\] vssd1 vssd1 vccd1 vccd1 net2150 sky130_fd_sc_hd__dlygate4sd3_1
X_09795_ _03765_ net404 net490 _04813_ vssd1 vssd1 vccd1 vccd1 _04814_ sky130_fd_sc_hd__o211a_1
XFILLER_0_99_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout565_A net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_55_Right_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1045 top.DUT.register\[9\]\[23\] vssd1 vssd1 vccd1 vccd1 net2161 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1056 top.DUT.register\[7\]\[29\] vssd1 vssd1 vccd1 vccd1 net2172 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1067 top.DUT.register\[3\]\[27\] vssd1 vssd1 vccd1 vccd1 net2183 sky130_fd_sc_hd__dlygate4sd3_1
X_08746_ _02092_ _03833_ _03083_ vssd1 vssd1 vccd1 vccd1 _03863_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_197_427 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1078 top.DUT.register\[2\]\[22\] vssd1 vssd1 vccd1 vccd1 net2194 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1089 top.DUT.register\[27\]\[3\] vssd1 vssd1 vccd1 vccd1 net2205 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_197_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09132__A2 _04051_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08677_ net306 _03796_ _03794_ vssd1 vssd1 vccd1 vccd1 _03797_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout353_X net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout732_A _01627_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_77_Left_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_200_3450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09683__A3 top.a1.instruction\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10300__S net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07628_ top.DUT.register\[30\]\[5\] net579 _02764_ _02766_ vssd1 vssd1 vccd1 vccd1
+ _02767_ sky130_fd_sc_hd__a211o_1
XFILLER_0_95_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07694__A2 net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_165_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout520_X net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07559_ top.DUT.register\[26\]\[7\] net750 net742 top.DUT.register\[2\]\[7\] vssd1
+ vssd1 vccd1 vccd1 _02698_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout618_X net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_181_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10570_ net1528 net247 net350 vssd1 vssd1 vccd1 vccd1 _00736_ sky130_fd_sc_hd__mux2_1
XANTENNA__07446__A2 net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09840__B1 _04151_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_64_Right_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06654__B1 net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09229_ top.pc\[9\] _04284_ vssd1 vssd1 vccd1 vccd1 _04297_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_134_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12240_ top.lcd.cnt_20ms\[11\] _06074_ vssd1 vssd1 vccd1 vccd1 _06075_ sky130_fd_sc_hd__and2_1
XFILLER_0_121_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout987_X net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_86_Left_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12524__Q top.a1.halfData\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08946__A2 net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12171_ net1362 net846 net796 _06025_ vssd1 vssd1 vccd1 vccd1 _01279_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_75_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_674 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11122_ net907 net1703 net862 _05066_ vssd1 vssd1 vccd1 vccd1 _01212_ sky130_fd_sc_hd__a31o_1
Xhold890 top.DUT.register\[3\]\[15\] vssd1 vssd1 vccd1 vccd1 net2006 sky130_fd_sc_hd__dlygate4sd3_1
X_11053_ net99 net870 net834 net1222 vssd1 vssd1 vccd1 vccd1 _01164_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_166_2939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13097__RESET_B net1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10004_ net174 net1809 net624 vssd1 vssd1 vccd1 vccd1 _00209_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_73_Right_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_199_3427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_199_3438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06748__X _01887_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11955_ _05770_ _05776_ _05788_ _05837_ vssd1 vssd1 vccd1 vccd1 _05838_ sky130_fd_sc_hd__o31a_1
X_10906_ net1792 net204 net480 vssd1 vssd1 vccd1 vccd1 _01067_ sky130_fd_sc_hd__mux2_1
XANTENNA__10210__S net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07685__A2 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11886_ _05699_ _05730_ vssd1 vssd1 vccd1 vccd1 _05769_ sky130_fd_sc_hd__nor2_1
XANTENNA__06893__B1 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13625_ clknet_leaf_72_clk _01212_ net1082 vssd1 vssd1 vccd1 vccd1 net52 sky130_fd_sc_hd__dfrtp_1
X_10837_ net1453 net207 net475 vssd1 vssd1 vccd1 vccd1 _00998_ sky130_fd_sc_hd__mux2_1
XFILLER_0_172_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11252__D _05118_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12661__RESET_B net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_82_Right_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_15_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06483__X _01622_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13556_ clknet_leaf_105_clk _01143_ net969 vssd1 vssd1 vccd1 vccd1 top.ramload\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07437__A2 net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10768_ net1329 net237 net483 vssd1 vssd1 vccd1 vccd1 _00929_ sky130_fd_sc_hd__mux2_1
XANTENNA__09831__B1 _04151_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09300__A top.pc\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06645__B1 net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12507_ clknet_leaf_78_clk _00099_ net1074 vssd1 vssd1 vccd1 vccd1 top.pc\[19\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_82_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13487_ clknet_leaf_22_clk _01079_ net1033 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[30\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_10699_ net1573 net261 net335 vssd1 vssd1 vccd1 vccd1 _00860_ sky130_fd_sc_hd__mux2_1
X_12438_ clknet_leaf_88_clk _00034_ net1001 vssd1 vssd1 vccd1 vccd1 top.ramaddr\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_799 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_2197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12434__Q top.ramaddr\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08937__A2 _04041_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10880__S net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12369_ clknet_leaf_103_clk top.ru.next_FetchedData\[13\] net974 vssd1 vssd1 vccd1
+ vccd1 top.a1.dataIn\[13\] sky130_fd_sc_hd__dfrtp_2
XANTENNA__06930__Y _02069_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07070__B1 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_91_Right_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_130_2397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09347__C1 net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06930_ _02059_ _02068_ vssd1 vssd1 vccd1 vccd1 _02069_ sky130_fd_sc_hd__nor2_4
XFILLER_0_38_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06861_ top.DUT.register\[1\]\[19\] net756 net745 top.DUT.register\[2\]\[19\] _01999_
+ vssd1 vssd1 vccd1 vccd1 _02000_ sky130_fd_sc_hd__a221o_1
X_08600_ _03713_ _03720_ _03723_ vssd1 vssd1 vccd1 vccd1 _03724_ sky130_fd_sc_hd__or3b_2
XFILLER_0_179_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06792_ top.DUT.register\[15\]\[17\] net680 net676 top.DUT.register\[31\]\[17\] vssd1
+ vssd1 vccd1 vccd1 _01931_ sky130_fd_sc_hd__a22o_1
X_09580_ _01679_ _04620_ _04622_ _04623_ vssd1 vssd1 vccd1 vccd1 _04627_ sky130_fd_sc_hd__a211o_1
XFILLER_0_145_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09114__A2 net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08531_ _03614_ _03657_ _02307_ vssd1 vssd1 vccd1 vccd1 _03658_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_54_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_194_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10120__S net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08462_ _02571_ _03591_ vssd1 vssd1 vccd1 vccd1 _03592_ sky130_fd_sc_hd__xnor2_1
XANTENNA__08873__A1 net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07676__A2 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07413_ top.DUT.register\[28\]\[9\] net766 net738 top.DUT.register\[12\]\[9\] vssd1
+ vssd1 vccd1 vccd1 _02552_ sky130_fd_sc_hd__a22o_1
XANTENNA__10680__A1 net206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08393_ net312 _03394_ vssd1 vssd1 vccd1 vccd1 _03525_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_34_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06884__B1 net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_137_2507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout146_A net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07344_ top.DUT.register\[26\]\[8\] net527 net524 top.DUT.register\[11\]\[8\] vssd1
+ vssd1 vccd1 vccd1 _02483_ sky130_fd_sc_hd__a22o_1
XANTENNA__06393__X _01532_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08525__S net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_95 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06636__B1 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07275_ top.DUT.register\[21\]\[13\] net657 net741 top.DUT.register\[12\]\[13\] _02413_
+ vssd1 vssd1 vccd1 vccd1 _02414_ sky130_fd_sc_hd__a221o_1
XFILLER_0_45_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout313_A net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_120_clk_X clknet_leaf_120_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1055_A net1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06226_ top.ramload\[20\] net858 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedInstr\[20\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_103_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09014_ _03642_ _03763_ _03907_ _04088_ vssd1 vssd1 vccd1 vccd1 _04089_ sky130_fd_sc_hd__or4_1
XFILLER_0_5_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12185__A1 top.a1.row2\[40\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold120 _01188_ vssd1 vssd1 vccd1 vccd1 net1236 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10790__S net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06157_ top.a1.dataIn\[8\] vssd1 vssd1 vccd1 vccd1 _01400_ sky130_fd_sc_hd__inv_2
XFILLER_0_13_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold131 top.ramstore\[2\] vssd1 vssd1 vccd1 vccd1 net1247 sky130_fd_sc_hd__dlygate4sd3_1
Xhold142 top.a1.row2\[25\] vssd1 vssd1 vccd1 vccd1 net1258 sky130_fd_sc_hd__dlygate4sd3_1
Xhold153 net122 vssd1 vssd1 vccd1 vccd1 net1269 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07665__A top.a1.instruction\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07061__B1 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold164 top.DUT.register\[4\]\[1\] vssd1 vssd1 vccd1 vccd1 net1280 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07600__A2 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold175 top.ramaddr\[3\] vssd1 vssd1 vccd1 vccd1 net1291 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout682_A _01547_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold186 top.a1.row1\[13\] vssd1 vssd1 vccd1 vccd1 net1302 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout600 net601 vssd1 vssd1 vccd1 vccd1 net600 sky130_fd_sc_hd__clkbuf_8
Xhold197 top.DUT.register\[24\]\[10\] vssd1 vssd1 vccd1 vccd1 net1313 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout611 net612 vssd1 vssd1 vccd1 vccd1 net611 sky130_fd_sc_hd__clkbuf_8
Xfanout622 _04953_ vssd1 vssd1 vccd1 vccd1 net622 sky130_fd_sc_hd__buf_6
X_09916_ _04151_ _04922_ vssd1 vssd1 vccd1 vccd1 _04923_ sky130_fd_sc_hd__nor2_1
XANTENNA__07384__B _02522_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout633 _04714_ vssd1 vssd1 vccd1 vccd1 net633 sky130_fd_sc_hd__buf_6
XFILLER_0_186_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout644 _01613_ vssd1 vssd1 vccd1 vccd1 net644 sky130_fd_sc_hd__clkbuf_4
XANTENNA_clkbuf_3_6_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout655 _01609_ vssd1 vssd1 vccd1 vccd1 net655 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_95_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_148_2669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout666 _01605_ vssd1 vssd1 vccd1 vccd1 net666 sky130_fd_sc_hd__clkbuf_4
X_09847_ net827 _04523_ _04859_ vssd1 vssd1 vccd1 vccd1 _04860_ sky130_fd_sc_hd__o21ba_1
Xfanout677 _01548_ vssd1 vssd1 vccd1 vccd1 net677 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout470_X net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout688 _06049_ vssd1 vssd1 vccd1 vccd1 net688 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout947_A net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout699 _01643_ vssd1 vssd1 vccd1 vccd1 net699 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_70_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout568_X net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09778_ top.pc\[16\] _04420_ vssd1 vssd1 vccd1 vccd1 _04798_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_161_2858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_198_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_197_246 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08729_ net430 _03845_ _03846_ net427 _03844_ vssd1 vssd1 vccd1 vccd1 _03847_ sky130_fd_sc_hd__a221o_1
XFILLER_0_96_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_201_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_200_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout735_X net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08313__B1 net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11740_ _05587_ _05621_ _05622_ _05588_ vssd1 vssd1 vccd1 vccd1 _05623_ sky130_fd_sc_hd__a22oi_4
XANTENNA__10030__S net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_205_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_194_3357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06875__B1 net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11671_ _01398_ _05549_ _05525_ vssd1 vssd1 vccd1 vccd1 _05554_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_166_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_153_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13410_ clknet_leaf_10_clk _01002_ net950 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[28\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_10622_ net164 net1517 net349 vssd1 vssd1 vccd1 vccd1 _00787_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_12_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_582 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06627__B1 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09120__A _02904_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13341_ clknet_leaf_127_clk _00933_ net930 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[26\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_91_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10553_ net1666 net176 net356 vssd1 vssd1 vccd1 vccd1 _00720_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_94_Left_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13272_ clknet_leaf_127_clk _00864_ net929 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[24\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_10484_ net1970 net192 net363 vssd1 vssd1 vccd1 vccd1 _00654_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_596 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12176__B2 net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12223_ _06052_ _06064_ vssd1 vssd1 vccd1 vccd1 _06065_ sky130_fd_sc_hd__nor2_1
XFILLER_0_121_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07052__B1 net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12154_ _01403_ _06036_ vssd1 vssd1 vccd1 vccd1 _06037_ sky130_fd_sc_hd__and2_1
X_11105_ net43 net869 vssd1 vssd1 vccd1 vccd1 _05058_ sky130_fd_sc_hd__and2_1
XANTENNA__10205__S net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12085_ _05958_ _05959_ _05962_ _05967_ vssd1 vssd1 vccd1 vccd1 _05968_ sky130_fd_sc_hd__or4bb_4
XANTENNA__12516__SET_B net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11036_ net16 net838 net816 top.ramload\[22\] vssd1 vssd1 vccd1 vccd1 _01148_ sky130_fd_sc_hd__o22a_1
XANTENNA__06478__X _01617_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12987_ clknet_leaf_125_clk _00579_ net924 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[15\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_176_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11938_ _05783_ _05820_ vssd1 vssd1 vccd1 vccd1 _05821_ sky130_fd_sc_hd__nor2_1
XFILLER_0_59_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08855__B2 net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10875__S net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_200_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11869_ _05740_ _05748_ _05750_ vssd1 vssd1 vccd1 vccd1 _05752_ sky130_fd_sc_hd__a21o_1
XFILLER_0_7_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_31_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13608_ clknet_leaf_74_clk _01195_ net1078 vssd1 vssd1 vccd1 vccd1 net65 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_172_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_119_2226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_119_2237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06618__B1 net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13539_ clknet_leaf_104_clk _01126_ net973 vssd1 vssd1 vccd1 vccd1 top.ramload\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_41_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_41_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06373__B top.a1.instruction\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_200_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07060_ _02198_ vssd1 vssd1 vccd1 vccd1 _02199_ sky130_fd_sc_hd__inv_2
XANTENNA__07830__A2 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_2426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_140_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07043__B1 net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07962_ _01659_ _03100_ vssd1 vssd1 vccd1 vccd1 _03101_ sky130_fd_sc_hd__nand2_1
XANTENNA__10115__S net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09701_ net2242 net261 net633 vssd1 vssd1 vccd1 vccd1 _00124_ sky130_fd_sc_hd__mux2_1
XANTENNA__08535__A1_N net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06913_ top.DUT.register\[22\]\[21\] net577 net509 top.DUT.register\[4\]\[21\] _02051_
+ vssd1 vssd1 vccd1 vccd1 _02052_ sky130_fd_sc_hd__a221o_1
XFILLER_0_4_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07893_ top.DUT.register\[17\]\[1\] net462 _03031_ vssd1 vssd1 vccd1 vccd1 _03032_
+ sky130_fd_sc_hd__a21o_1
XANTENNA__08587__Y _03711_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09632_ top.pad.keyCode\[1\] top.pad.keyCode\[0\] top.pad.keyCode\[2\] top.pad.keyCode\[3\]
+ vssd1 vssd1 vccd1 vccd1 _04674_ sky130_fd_sc_hd__or4b_2
X_06844_ _01973_ _01982_ vssd1 vssd1 vccd1 vccd1 _01983_ sky130_fd_sc_hd__or2_4
XANTENNA__07897__A2 net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09563_ net138 _04599_ _04604_ net134 _04611_ vssd1 vssd1 vccd1 vccd1 _04612_ sky130_fd_sc_hd__o221a_1
X_06775_ top.DUT.register\[24\]\[24\] net645 net752 top.DUT.register\[26\]\[24\] _01913_
+ vssd1 vssd1 vccd1 vccd1 _01914_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_143_2588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08514_ _03067_ _03640_ vssd1 vssd1 vccd1 vccd1 _03641_ sky130_fd_sc_hd__nand2_1
XFILLER_0_194_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_188_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07649__A2 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09494_ _04528_ _04530_ vssd1 vssd1 vccd1 vccd1 _04547_ sky130_fd_sc_hd__nand2_1
XFILLER_0_172_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08445_ _02498_ net300 _03280_ vssd1 vssd1 vccd1 vccd1 _03575_ sky130_fd_sc_hd__o21ai_1
XANTENNA__10785__S net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_42_clk_A clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_176_3087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout528_A net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08376_ _02801_ _03486_ _02800_ vssd1 vssd1 vccd1 vccd1 _03509_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_34_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_190_444 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06609__B1 net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07327_ top.DUT.register\[6\]\[12\] net636 _02454_ _02465_ vssd1 vssd1 vccd1 vccd1
+ _02466_ sky130_fd_sc_hd__a211o_1
XFILLER_0_151_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_483 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout316_X net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_59_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07258_ top.DUT.register\[6\]\[13\] net569 net520 top.DUT.register\[10\]\[13\] vssd1
+ vssd1 vccd1 vccd1 _02397_ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_57_clk_A clknet_4_12__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07821__A2 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout897_A net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06209_ net1284 net859 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedInstr\[3\] sky130_fd_sc_hd__and2_1
X_07189_ _02321_ _02323_ _02325_ _02327_ vssd1 vssd1 vccd1 vccd1 _02328_ sky130_fd_sc_hd__or4_4
XANTENNA_clkbuf_leaf_100_clk_A clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07034__B1 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_72_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06388__A2 top.a1.instruction\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10025__S net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout430 _03257_ vssd1 vssd1 vccd1 vccd1 net430 sky130_fd_sc_hd__buf_2
Xfanout441 _01566_ vssd1 vssd1 vccd1 vccd1 net441 sky130_fd_sc_hd__buf_6
Xfanout452 _01561_ vssd1 vssd1 vccd1 vccd1 net452 sky130_fd_sc_hd__clkbuf_4
Xfanout463 net466 vssd1 vssd1 vccd1 vccd1 net463 sky130_fd_sc_hd__clkbuf_8
XANTENNA_clkbuf_leaf_115_clk_A clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout852_X net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout474 net477 vssd1 vssd1 vccd1 vccd1 net474 sky130_fd_sc_hd__buf_6
Xfanout485 _04962_ vssd1 vssd1 vccd1 vccd1 net485 sky130_fd_sc_hd__buf_4
XANTENNA__08938__B _04045_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12910_ clknet_leaf_39_clk _00502_ net1055 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[12\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout496 net498 vssd1 vssd1 vccd1 vccd1 net496 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07888__A2 net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06739__A _01877_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09115__A _03000_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_555 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12841_ clknet_leaf_51_clk _00433_ net1035 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[10\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_17_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_408 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12772_ clknet_leaf_36_clk _00364_ net1051 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[8\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08837__A1 net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_169_Left_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_255 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06848__B1 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11723_ _05568_ _05604_ vssd1 vssd1 vccd1 vccd1 _05606_ sky130_fd_sc_hd__xnor2_2
XANTENNA__09769__B _04403_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11654_ _05507_ _05510_ _05517_ _05536_ vssd1 vssd1 vccd1 vccd1 _05537_ sky130_fd_sc_hd__a31o_1
XANTENNA__08018__X _03157_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10605_ net231 net2039 net346 vssd1 vssd1 vccd1 vccd1 _00770_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_181_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11585_ _05467_ vssd1 vssd1 vccd1 vccd1 _05468_ sky130_fd_sc_hd__inv_2
XFILLER_0_181_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_291 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13324_ clknet_leaf_62_clk _00916_ net1089 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[25\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07273__B1 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10536_ net1831 net243 net354 vssd1 vssd1 vccd1 vccd1 _00703_ sky130_fd_sc_hd__mux2_1
XANTENNA__08470__C1 _03598_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13255_ clknet_leaf_8_clk _00847_ net945 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[23\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_108_Right_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_178_Left_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10467_ net1346 net257 net363 vssd1 vssd1 vccd1 vccd1 _00637_ sky130_fd_sc_hd__mux2_1
XANTENNA__06480__Y _01619_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_114_2156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07025__B1 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12206_ top.lcd.cnt_20ms\[4\] top.lcd.cnt_20ms\[3\] _06051_ vssd1 vssd1 vccd1 vccd1
+ _06052_ sky130_fd_sc_hd__and3_1
X_13186_ clknet_leaf_9_clk _00778_ net947 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[21\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_10398_ net1798 net267 net370 vssd1 vssd1 vccd1 vccd1 _00570_ sky130_fd_sc_hd__mux2_1
X_12137_ _06014_ _06017_ _06018_ vssd1 vssd1 vccd1 vccd1 _06020_ sky130_fd_sc_hd__nor3_1
X_12068_ _05940_ _05949_ vssd1 vssd1 vccd1 vccd1 _05951_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_205_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11019_ net29 net842 net819 net1274 vssd1 vssd1 vccd1 vccd1 _01131_ sky130_fd_sc_hd__a22o_1
XANTENNA__06649__A _01764_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_200 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06551__A2 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06368__B net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13249__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_408 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08828__A1 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06560_ _01678_ _01698_ vssd1 vssd1 vccd1 vccd1 _01699_ sky130_fd_sc_hd__nor2_1
XFILLER_0_176_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06839__B1 net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06491_ net788 _01602_ _01607_ vssd1 vssd1 vccd1 vccd1 _01630_ sky130_fd_sc_hd__and3_4
XFILLER_0_118_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08230_ net315 _03366_ vssd1 vssd1 vccd1 vccd1 _03367_ sky130_fd_sc_hd__or2_1
XFILLER_0_145_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_157_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_184_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08161_ net285 _03298_ _03284_ net280 vssd1 vssd1 vccd1 vccd1 _03299_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_172_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_656 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07112_ top.DUT.register\[28\]\[16\] net767 net714 top.DUT.register\[27\]\[16\] vssd1
+ vssd1 vccd1 vccd1 _02251_ sky130_fd_sc_hd__a22o_1
X_08092_ _02678_ net300 vssd1 vssd1 vccd1 vccd1 _03231_ sky130_fd_sc_hd__or2_1
XANTENNA__07264__B1 net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07803__A2 net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload40 clknet_leaf_97_clk vssd1 vssd1 vccd1 vccd1 clkload40/Y sky130_fd_sc_hd__inv_16
X_07043_ top.DUT.register\[6\]\[22\] net568 net564 top.DUT.register\[20\]\[22\] vssd1
+ vssd1 vccd1 vccd1 _02182_ sky130_fd_sc_hd__a22o_1
Xclkload51 clknet_leaf_85_clk vssd1 vssd1 vccd1 vccd1 clkload51/Y sky130_fd_sc_hd__inv_12
Xclkload62 clknet_leaf_26_clk vssd1 vssd1 vccd1 vccd1 clkload62/Y sky130_fd_sc_hd__inv_8
XANTENNA__07927__B _02385_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload73 clknet_leaf_34_clk vssd1 vssd1 vccd1 vccd1 clkload73/Y sky130_fd_sc_hd__clkinv_8
Xclkload84 clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 clkload84/X sky130_fd_sc_hd__clkbuf_4
Xclkload95 clknet_leaf_72_clk vssd1 vssd1 vccd1 vccd1 clkload95/Y sky130_fd_sc_hd__inv_8
XFILLER_0_55_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08994_ _03691_ _03718_ _04066_ _04068_ vssd1 vssd1 vccd1 vccd1 _04069_ sky130_fd_sc_hd__or4_1
XFILLER_0_76_61 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1018_A net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09308__A2 _02408_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07945_ _02090_ _02091_ _02156_ _02176_ vssd1 vssd1 vccd1 vccd1 _03084_ sky130_fd_sc_hd__o211a_1
XFILLER_0_167_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_145_2617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_2628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout478_A _04964_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06790__A2 net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07662__B _02798_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07876_ top.DUT.register\[21\]\[1\] net657 net637 top.DUT.register\[6\]\[1\] _03014_
+ vssd1 vssd1 vccd1 vccd1 _03015_ sky130_fd_sc_hd__a221o_1
XFILLER_0_183_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09615_ top.a1.state\[2\] _04657_ top.a1.state\[1\] top.a1.state\[0\] vssd1 vssd1
+ vccd1 vccd1 _04660_ sky130_fd_sc_hd__or4bb_2
X_06827_ top.DUT.register\[28\]\[19\] net557 net449 top.DUT.register\[21\]\[19\] _01965_
+ vssd1 vssd1 vccd1 vccd1 _01966_ sky130_fd_sc_hd__a221o_1
XFILLER_0_211_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_178_3116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout645_A _01613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06542__A2 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09546_ net138 _04589_ net902 vssd1 vssd1 vccd1 vccd1 _04596_ sky130_fd_sc_hd__o21ai_1
X_06758_ _01887_ _01896_ vssd1 vssd1 vccd1 vccd1 _01897_ sky130_fd_sc_hd__nor2_2
XFILLER_0_210_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_195_547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_191_3305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09477_ _04529_ _04530_ vssd1 vssd1 vccd1 vccd1 _04531_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_191_3316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06689_ _01823_ _01825_ _01827_ vssd1 vssd1 vccd1 vccd1 _01828_ sky130_fd_sc_hd__or3_1
XFILLER_0_176_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout433_X net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_148_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08428_ net315 _03204_ vssd1 vssd1 vccd1 vccd1 _03559_ sky130_fd_sc_hd__nor2_1
XFILLER_0_109_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkload1 clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 clkload1/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_18_163 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08359_ _03355_ _03365_ net304 vssd1 vssd1 vccd1 vccd1 _03492_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout600_X net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_156_2779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07255__B1 net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_210_3600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_190_285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11370_ top.a1.dataIn\[19\] _05249_ _05250_ vssd1 vssd1 vccd1 vccd1 _05253_ sky130_fd_sc_hd__and3_1
XANTENNA__09795__A2 net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10321_ net168 net2113 net381 vssd1 vssd1 vccd1 vccd1 _00498_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_189_3278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_363 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07007__B1 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13040_ clknet_leaf_29_clk _00632_ net1017 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[16\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_10252_ net180 net1806 net392 vssd1 vssd1 vccd1 vccd1 _00431_ sky130_fd_sc_hd__mux2_1
X_10183_ _04154_ net689 _04947_ vssd1 vssd1 vccd1 vccd1 _04963_ sky130_fd_sc_hd__or3b_2
XTAP_TAPCELL_ROW_208_3562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input39_A nrst vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_208_3573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout260 net262 vssd1 vssd1 vccd1 vccd1 net260 sky130_fd_sc_hd__clkbuf_2
XANTENNA__11106__A2 top.ramaddr\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout282 _03171_ vssd1 vssd1 vccd1 vccd1 net282 sky130_fd_sc_hd__buf_2
Xfanout293 net294 vssd1 vssd1 vccd1 vccd1 net293 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_202_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_85_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06533__A2 net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12824_ clknet_leaf_127_clk _00416_ net918 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[10\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_186_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12755_ clknet_leaf_122_clk _00347_ net928 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[8\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09499__B _04543_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_761 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11706_ _05586_ _05587_ vssd1 vssd1 vccd1 vccd1 _05589_ sky130_fd_sc_hd__nand2_1
XANTENNA__11290__A1 net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_794 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12686_ clknet_leaf_43_clk _00278_ net1062 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[5\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_166_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11637_ _05480_ _05519_ _05512_ vssd1 vssd1 vccd1 vccd1 _05520_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09235__A1 _02497_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_182_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_360 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06491__X _01630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11568_ _01397_ net250 vssd1 vssd1 vccd1 vccd1 _05451_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_188_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13307_ clknet_leaf_120_clk _00899_ net931 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[25\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold708 top.DUT.register\[21\]\[5\] vssd1 vssd1 vccd1 vccd1 net1824 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10519_ net1782 net177 net358 vssd1 vssd1 vccd1 vccd1 _00688_ sky130_fd_sc_hd__mux2_1
Xhold719 top.DUT.register\[16\]\[13\] vssd1 vssd1 vccd1 vccd1 net1835 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_150_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11499_ _05353_ _05381_ vssd1 vssd1 vccd1 vccd1 _05382_ sky130_fd_sc_hd__or2_1
XFILLER_0_0_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_514 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13238_ clknet_leaf_4_clk _00830_ net942 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[23\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_198_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13169_ clknet_leaf_116_clk _00761_ net958 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[21\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06772__A2 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07730_ top.DUT.register\[26\]\[3\] net752 net708 top.DUT.register\[15\]\[3\] vssd1
+ vssd1 vccd1 vccd1 _02869_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_127_2347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06379__A top.a1.instruction\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_2358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_211_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09710__A2 net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07661_ _02773_ _02798_ vssd1 vssd1 vccd1 vccd1 _02800_ sky130_fd_sc_hd__nand2_1
XANTENNA__06524__A2 net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_695 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09400_ net133 _04451_ _04458_ net811 net900 vssd1 vssd1 vccd1 vccd1 _04459_ sky130_fd_sc_hd__o221a_1
X_06612_ top.DUT.register\[6\]\[27\] net569 net457 top.DUT.register\[25\]\[27\] _01750_
+ vssd1 vssd1 vccd1 vccd1 _01751_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_0_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_2547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08594__A net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07592_ top.DUT.register\[12\]\[6\] net738 net714 top.DUT.register\[27\]\[6\] vssd1
+ vssd1 vccd1 vccd1 _02731_ sky130_fd_sc_hd__a22o_1
XFILLER_0_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_153_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09331_ net136 _04379_ _04393_ net897 vssd1 vssd1 vccd1 vccd1 _04394_ sky130_fd_sc_hd__o211ai_1
X_06543_ top.DUT.register\[2\]\[29\] net744 net740 top.DUT.register\[12\]\[29\] vssd1
+ vssd1 vccd1 vccd1 _01682_ sky130_fd_sc_hd__a22o_1
XFILLER_0_177_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_614 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_173_3035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09262_ _04326_ _04327_ vssd1 vssd1 vccd1 vccd1 _04328_ sky130_fd_sc_hd__or2_1
XANTENNA__07485__B1 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_173_3046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06474_ _01601_ _01604_ vssd1 vssd1 vccd1 vccd1 _01613_ sky130_fd_sc_hd__nor2_4
XFILLER_0_117_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_173_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08213_ _03258_ _03350_ vssd1 vssd1 vccd1 vccd1 _03351_ sky130_fd_sc_hd__nor2_1
XANTENNA__09226__A1 net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09193_ _02773_ _02777_ _04245_ vssd1 vssd1 vccd1 vccd1 _04264_ sky130_fd_sc_hd__a21o_1
XFILLER_0_105_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout226_A _04805_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_173_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08144_ _03280_ _03281_ vssd1 vssd1 vccd1 vccd1 _03282_ sky130_fd_sc_hd__nand2_1
XANTENNA__09777__A2 _04403_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07788__B2 top.DUT.register\[19\]\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08075_ _02026_ net299 vssd1 vssd1 vccd1 vccd1 _03214_ sky130_fd_sc_hd__nand2_1
XFILLER_0_141_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07026_ top.DUT.register\[10\]\[20\] net773 net704 top.DUT.register\[3\]\[20\] vssd1
+ vssd1 vccd1 vccd1 _02165_ sky130_fd_sc_hd__a22o_1
XFILLER_0_30_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12945__RESET_B net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout595_A _04966_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12352__Q top.edg2.flip1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13414__CLK clknet_leaf_40_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold13 _00011_ vssd1 vssd1 vccd1 vccd1 net1129 sky130_fd_sc_hd__dlygate4sd3_1
Xhold24 _01177_ vssd1 vssd1 vccd1 vccd1 net1140 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08121__X _03260_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08977_ _03180_ net498 _03336_ _03385_ vssd1 vssd1 vccd1 vccd1 _04052_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout762_A net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold35 top.a1.data\[7\] vssd1 vssd1 vccd1 vccd1 net1151 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout383_X net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold46 top.ramstore\[25\] vssd1 vssd1 vccd1 vccd1 net1162 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07960__A1 _01679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06763__A2 net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold57 top.ramstore\[22\] vssd1 vssd1 vccd1 vccd1 net1173 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10303__S net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07928_ _02286_ _02305_ _02310_ _03066_ vssd1 vssd1 vccd1 vccd1 _03067_ sky130_fd_sc_hd__o22a_1
Xhold68 net98 vssd1 vssd1 vccd1 vccd1 net1184 sky130_fd_sc_hd__dlygate4sd3_1
Xhold79 top.lcd.cnt_20ms\[15\] vssd1 vssd1 vccd1 vccd1 net1195 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09162__B1 net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout550_X net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07859_ _02359_ _02901_ _02997_ net805 vssd1 vssd1 vccd1 vccd1 _02998_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout648_X net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_195_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_168_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_67_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_203_3492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10870_ net197 net2073 net596 vssd1 vssd1 vccd1 vccd1 _01031_ sky130_fd_sc_hd__mux2_1
XFILLER_0_195_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_27_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_27_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09529_ _04578_ _04579_ vssd1 vssd1 vccd1 vccd1 _04580_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_158_2819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09465__A1 net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout815_X net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_195_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_210_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12540_ clknet_leaf_0_clk _00132_ net915 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[1\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07476__B1 net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12527__Q top.a1.halfData\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12471_ clknet_leaf_47_clk _00066_ net1067 vssd1 vssd1 vccd1 vccd1 top.ramstore\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_483 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_193_Right_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11422_ _05303_ _05304_ vssd1 vssd1 vccd1 vccd1 _05305_ sky130_fd_sc_hd__nand2_1
XANTENNA__07228__B1 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12221__B1 net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09768__A2 _04386_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11353_ _05227_ _05235_ vssd1 vssd1 vccd1 vccd1 _05236_ sky130_fd_sc_hd__nor2_1
XANTENNA__08440__A2 net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_111_2104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10304_ net237 net2010 net384 vssd1 vssd1 vccd1 vccd1 _00481_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_111_2115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_1870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11089__B net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11284_ top.a1.row2\[11\] _05139_ _05145_ top.a1.row2\[19\] vssd1 vssd1 vccd1 vccd1
+ _05174_ sky130_fd_sc_hd__a22o_1
XFILLER_0_30_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13094__CLK clknet_leaf_40_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13023_ clknet_leaf_19_clk _00615_ net1026 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[16\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_10235_ net252 net1826 net392 vssd1 vssd1 vccd1 vccd1 _00414_ sky130_fd_sc_hd__mux2_1
Xfanout1000 net1007 vssd1 vssd1 vccd1 vccd1 net1000 sky130_fd_sc_hd__clkbuf_4
Xfanout1011 net1016 vssd1 vssd1 vccd1 vccd1 net1011 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07400__B1 net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06203__B2 net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1022 net1025 vssd1 vssd1 vccd1 vccd1 net1022 sky130_fd_sc_hd__clkbuf_2
X_10166_ net1628 net201 net604 vssd1 vssd1 vccd1 vccd1 _00365_ sky130_fd_sc_hd__mux2_1
Xfanout1033 net1036 vssd1 vssd1 vccd1 vccd1 net1033 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06754__A2 net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1044 net1048 vssd1 vssd1 vccd1 vccd1 net1044 sky130_fd_sc_hd__clkbuf_4
Xfanout1055 net1071 vssd1 vssd1 vccd1 vccd1 net1055 sky130_fd_sc_hd__clkbuf_4
Xfanout1066 net1067 vssd1 vssd1 vccd1 vccd1 net1066 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10213__S net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1077 net1079 vssd1 vssd1 vccd1 vccd1 net1077 sky130_fd_sc_hd__clkbuf_4
Xfanout1088 net1096 vssd1 vssd1 vccd1 vccd1 net1088 sky130_fd_sc_hd__clkbuf_4
X_10097_ net1589 net215 net611 vssd1 vssd1 vccd1 vccd1 _00298_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_109_2077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_2088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06506__A2 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload4_A clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_694 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12807_ clknet_leaf_7_clk _00399_ net944 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[9\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_122_2277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13787_ clknet_leaf_68_clk _01356_ vssd1 vssd1 vccd1 vccd1 top.pad.button_control.r_counter\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_10999_ top.a1.dataInTemp\[9\] net785 vssd1 vssd1 vccd1 vccd1 _05033_ sky130_fd_sc_hd__or2_1
XFILLER_0_186_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09797__X _04815_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12738_ clknet_leaf_10_clk _00330_ net949 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[7\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07467__B1 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_155_742 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10883__S net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_228 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12669_ clknet_leaf_13_clk _00261_ net941 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[5\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_72_559 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06190_ top.a1.hexop\[2\] top.a1.hexop\[1\] top.a1.hexop\[3\] top.a1.hexop\[4\] vssd1
+ vssd1 vccd1 vccd1 _01426_ sky130_fd_sc_hd__or4_1
XFILLER_0_108_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_160_Right_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_464 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold505 top.DUT.register\[27\]\[4\] vssd1 vssd1 vccd1 vccd1 net1621 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_648 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold516 top.DUT.register\[15\]\[20\] vssd1 vssd1 vccd1 vccd1 net1632 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_812 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold527 top.DUT.register\[28\]\[22\] vssd1 vssd1 vccd1 vccd1 net1643 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold538 top.DUT.register\[5\]\[9\] vssd1 vssd1 vccd1 vccd1 net1654 sky130_fd_sc_hd__dlygate4sd3_1
Xhold549 top.DUT.register\[9\]\[26\] vssd1 vssd1 vccd1 vccd1 net1665 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11318__A2 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06993__A2 _02131_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08900_ _03988_ _04008_ vssd1 vssd1 vccd1 vccd1 _04010_ sky130_fd_sc_hd__or2_1
X_09880_ _04879_ _04881_ _04880_ vssd1 vssd1 vccd1 vccd1 _04890_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_51_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08831_ _01834_ net495 _03942_ _03943_ vssd1 vssd1 vccd1 vccd1 _03944_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_5_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06745__A2 net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08762_ net282 _03877_ vssd1 vssd1 vccd1 vccd1 _03878_ sky130_fd_sc_hd__or2_1
XANTENNA__10123__S net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08876__X _03987_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07713_ _02850_ _02851_ vssd1 vssd1 vccd1 vccd1 _02852_ sky130_fd_sc_hd__nand2b_2
X_08693_ _02179_ _03810_ vssd1 vssd1 vccd1 vccd1 _03812_ sky130_fd_sc_hd__xor2_1
XANTENNA__09695__A1 _03391_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07644_ top.DUT.register\[13\]\[5\] net777 net714 top.DUT.register\[27\]\[5\] vssd1
+ vssd1 vccd1 vccd1 _02783_ sky130_fd_sc_hd__a22o_1
XANTENNA__06396__X _01535_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07575_ top.DUT.register\[15\]\[6\] net679 net675 top.DUT.register\[31\]\[6\] vssd1
+ vssd1 vccd1 vccd1 _02714_ sky130_fd_sc_hd__a22o_1
XFILLER_0_165_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout343_A _04992_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09314_ top.pc\[14\] _04360_ vssd1 vssd1 vccd1 vccd1 _04377_ sky130_fd_sc_hd__and2_1
X_06526_ top.DUT.register\[9\]\[29\] net469 net441 top.DUT.register\[5\]\[29\] _01664_
+ vssd1 vssd1 vccd1 vccd1 _01665_ sky130_fd_sc_hd__a221o_1
XANTENNA__07458__B1 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_146_720 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11254__B2 top.a1.row2\[40\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_180_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold1193_A top.ramload\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09245_ _04310_ _04311_ vssd1 vssd1 vccd1 vccd1 _04312_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_62_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06457_ top.a1.instruction\[20\] top.a1.instruction\[21\] net792 vssd1 vssd1 vccd1
+ vccd1 _01596_ sky130_fd_sc_hd__and3_2
XANTENNA_fanout510_A _01565_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10793__S net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout229_X net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout608_A _04956_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_153_2738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09176_ _04246_ _04247_ vssd1 vssd1 vccd1 vccd1 _04248_ sky130_fd_sc_hd__nand2_1
X_06388_ top.a1.instruction\[15\] top.a1.instruction\[16\] net782 vssd1 vssd1 vccd1
+ vccd1 _01527_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_161_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08127_ top.ru.next_write_i _00006_ vssd1 vssd1 vccd1 vccd1 _03266_ sky130_fd_sc_hd__or2_1
XFILLER_0_43_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08058_ _01764_ net328 vssd1 vssd1 vccd1 vccd1 _03197_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_186_3237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07630__B1 net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout977_A net1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout598_X net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06984__A2 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11309__A2 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07009_ top.DUT.register\[28\]\[20\] net557 net544 top.DUT.register\[16\]\[20\] _02147_
+ vssd1 vssd1 vccd1 vccd1 _02148_ sky130_fd_sc_hd__a221o_1
Xoutput47 net47 vssd1 vssd1 vccd1 vccd1 ADR_O[16] sky130_fd_sc_hd__buf_2
Xoutput58 net58 vssd1 vssd1 vccd1 vccd1 ADR_O[26] sky130_fd_sc_hd__buf_2
Xoutput69 net69 vssd1 vssd1 vccd1 vccd1 ADR_O[7] sky130_fd_sc_hd__buf_2
XFILLER_0_11_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10020_ top.DUT.register\[4\]\[6\] net241 net619 vssd1 vssd1 vccd1 vccd1 _00223_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_168_2970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout765_X net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_205_3521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10033__S net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12954__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11971_ _05847_ _05853_ vssd1 vssd1 vccd1 vccd1 _05854_ sky130_fd_sc_hd__and2_1
XFILLER_0_169_823 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13710_ clknet_leaf_92_clk _01281_ net995 vssd1 vssd1 vccd1 vccd1 top.a1.row2\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_10922_ net1328 net266 _04960_ vssd1 vssd1 vccd1 vccd1 _01083_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07697__B1 net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07161__A2 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13641_ clknet_leaf_94_clk _00005_ net982 vssd1 vssd1 vccd1 vccd1 top.ru.state\[0\]
+ sky130_fd_sc_hd__dfstp_1
X_10853_ net1748 net153 net476 vssd1 vssd1 vccd1 vccd1 _01014_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_197_3399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_183_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07449__B1 net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13572_ clknet_leaf_91_clk _01159_ net996 vssd1 vssd1 vccd1 vccd1 net72 sky130_fd_sc_hd__dfrtp_2
X_10784_ net1759 net172 net484 vssd1 vssd1 vccd1 vccd1 _00945_ sky130_fd_sc_hd__mux2_1
X_12523_ clknet_leaf_71_clk _00115_ vssd1 vssd1 vccd1 vccd1 top.a1.halfData\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_164_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_239 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12454_ clknet_leaf_108_clk net34 net975 vssd1 vssd1 vccd1 vccd1 top.testpc.en_latched
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12867__RESET_B net1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08949__B1 _02796_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11405_ _05255_ _05256_ _05285_ vssd1 vssd1 vccd1 vccd1 _05288_ sky130_fd_sc_hd__a21boi_1
XANTENNA__10208__S net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12385_ clknet_leaf_110_clk top.ru.next_FetchedData\[29\] net989 vssd1 vssd1 vccd1
+ vccd1 top.a1.dataIn\[29\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_78_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11336_ _05214_ _05215_ _05217_ _05210_ vssd1 vssd1 vccd1 vccd1 _05219_ sky130_fd_sc_hd__a31o_1
XANTENNA__07621__B1 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06975__A2 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07584__Y _02723_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11267_ top.a1.row1\[121\] _05149_ _05150_ top.a1.row1\[105\] vssd1 vssd1 vccd1 vccd1
+ _05159_ sky130_fd_sc_hd__a22o_1
X_13006_ clknet_leaf_43_clk _00598_ net1062 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[15\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_10218_ net193 net1997 net395 vssd1 vssd1 vccd1 vccd1 _00398_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_105_Left_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11198_ _05105_ net1213 net472 vssd1 vssd1 vccd1 vccd1 _01249_ sky130_fd_sc_hd__mux2_1
XANTENNA__11181__B1 net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06727__A2 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10149_ net1366 net261 net604 vssd1 vssd1 vccd1 vccd1 _00348_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_124_2306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_206_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10878__S net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07152__A2 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_186_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_76 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07360_ top.a1.instruction\[29\] net789 net410 vssd1 vssd1 vccd1 vccd1 _02499_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_114_Left_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_102_1969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06311_ _01449_ _01461_ _01466_ _01448_ vssd1 vssd1 vccd1 vccd1 _00001_ sky130_fd_sc_hd__a22o_1
XFILLER_0_155_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07291_ _02429_ vssd1 vssd1 vccd1 vccd1 _02430_ sky130_fd_sc_hd__inv_2
XFILLER_0_45_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09030_ _03809_ _03850_ _03934_ _03972_ vssd1 vssd1 vccd1 vccd1 _04105_ sky130_fd_sc_hd__nand4_1
X_06242_ net1284 net854 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedData\[3\] sky130_fd_sc_hd__and2_1
XFILLER_0_60_507 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12827__CLK clknet_leaf_120_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_135_2468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10118__S net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06173_ top.a1.halfData\[1\] top.a1.halfData\[2\] top.a1.halfData\[3\] vssd1 vssd1
+ vccd1 vccd1 _01415_ sky130_fd_sc_hd__nand3b_1
Xhold302 top.DUT.register\[3\]\[18\] vssd1 vssd1 vccd1 vccd1 net1418 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold313 top.DUT.register\[1\]\[14\] vssd1 vssd1 vccd1 vccd1 net1429 sky130_fd_sc_hd__dlygate4sd3_1
Xhold324 top.DUT.register\[28\]\[11\] vssd1 vssd1 vccd1 vccd1 net1440 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold335 top.DUT.register\[6\]\[31\] vssd1 vssd1 vccd1 vccd1 net1451 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_159_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold346 top.ramaddr\[5\] vssd1 vssd1 vccd1 vccd1 net1462 sky130_fd_sc_hd__dlygate4sd3_1
Xhold357 top.DUT.register\[23\]\[17\] vssd1 vssd1 vccd1 vccd1 net1473 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06966__A2 net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold368 top.DUT.register\[25\]\[22\] vssd1 vssd1 vccd1 vccd1 net1484 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09932_ _04027_ net405 net490 _04937_ vssd1 vssd1 vccd1 vccd1 _04938_ sky130_fd_sc_hd__o211a_2
XANTENNA__07494__Y _02633_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold379 top.DUT.register\[17\]\[22\] vssd1 vssd1 vccd1 vccd1 net1495 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_123_Left_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout804 _01577_ vssd1 vssd1 vccd1 vccd1 net804 sky130_fd_sc_hd__clkbuf_4
Xfanout815 _01442_ vssd1 vssd1 vccd1 vccd1 net815 sky130_fd_sc_hd__clkbuf_8
Xfanout826 net829 vssd1 vssd1 vccd1 vccd1 net826 sky130_fd_sc_hd__buf_2
XFILLER_0_110_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08707__A3 _03441_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout837 _05045_ vssd1 vssd1 vccd1 vccd1 net837 sky130_fd_sc_hd__buf_8
X_09863_ net798 _04872_ _04873_ _04874_ vssd1 vssd1 vccd1 vccd1 _04875_ sky130_fd_sc_hd__a211o_1
XANTENNA__08112__A _02498_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout848 _04663_ vssd1 vssd1 vccd1 vccd1 net848 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout293_A net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06718__A2 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07915__A1 _02773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout859 top.ru.next_iready vssd1 vssd1 vccd1 vccd1 net859 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_181_3156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08814_ _03091_ _03927_ vssd1 vssd1 vccd1 vccd1 _03928_ sky130_fd_sc_hd__nor2_1
Xhold1002 top.DUT.register\[9\]\[2\] vssd1 vssd1 vccd1 vccd1 net2118 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_181_3167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1013 top.DUT.register\[18\]\[20\] vssd1 vssd1 vccd1 vccd1 net2129 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1000_A net1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1024 top.DUT.register\[24\]\[22\] vssd1 vssd1 vccd1 vccd1 net2140 sky130_fd_sc_hd__dlygate4sd3_1
X_09794_ net798 _04809_ _04810_ _04812_ vssd1 vssd1 vccd1 vccd1 _04813_ sky130_fd_sc_hd__a31o_1
Xhold1035 top.DUT.register\[24\]\[9\] vssd1 vssd1 vccd1 vccd1 net2151 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07391__A2 net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1046 top.DUT.register\[14\]\[20\] vssd1 vssd1 vccd1 vccd1 net2162 sky130_fd_sc_hd__dlygate4sd3_1
X_08745_ _02222_ net492 vssd1 vssd1 vccd1 vccd1 _03862_ sky130_fd_sc_hd__nor2_1
Xhold1057 top.DUT.register\[29\]\[8\] vssd1 vssd1 vccd1 vccd1 net2173 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1068 top.DUT.register\[30\]\[19\] vssd1 vssd1 vccd1 vccd1 net2184 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10788__S net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout460_A _01552_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1079 top.DUT.register\[1\]\[6\] vssd1 vssd1 vccd1 vccd1 net2195 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08766__B net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07679__B1 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08676_ _03755_ _03795_ net287 vssd1 vssd1 vccd1 vccd1 _03796_ sky130_fd_sc_hd__mux2_1
XFILLER_0_178_631 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_200_3440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07143__A2 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_200_3451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07627_ top.DUT.register\[9\]\[5\] net470 net515 top.DUT.register\[7\]\[5\] _02765_
+ vssd1 vssd1 vccd1 vccd1 _02766_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_132_Left_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout725_A _01630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08891__A2 net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout346_X net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1088_X net1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09878__A top.pc\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07558_ top.DUT.register\[24\]\[7\] net643 net639 top.DUT.register\[8\]\[7\] _02696_
+ vssd1 vssd1 vccd1 vccd1 _02697_ sky130_fd_sc_hd__a221o_1
XANTENNA__08782__A net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_2_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06509_ top.DUT.register\[24\]\[30\] net645 net704 top.DUT.register\[3\]\[30\] _01647_
+ vssd1 vssd1 vccd1 vccd1 _01648_ sky130_fd_sc_hd__a221o_1
XANTENNA__07669__Y _02808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07489_ top.DUT.register\[26\]\[14\] net528 net517 top.DUT.register\[7\]\[14\] vssd1
+ vssd1 vccd1 vccd1 _02628_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout513_X net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_146_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09228_ net898 top.pc\[8\] _04296_ net889 vssd1 vssd1 vccd1 vccd1 _00088_ sky130_fd_sc_hd__o211a_1
XFILLER_0_106_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07851__B1 net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12960__RESET_B net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12454__D net34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09159_ _04216_ _04219_ _04230_ vssd1 vssd1 vccd1 vccd1 _04232_ sky130_fd_sc_hd__a21o_1
XANTENNA__10028__S net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12170_ net1308 net846 net796 _06034_ vssd1 vssd1 vccd1 vccd1 _01278_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_141_Left_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout882_X net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06957__A2 net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11121_ net52 net867 vssd1 vssd1 vccd1 vccd1 _05066_ sky130_fd_sc_hd__and2_1
XFILLER_0_7_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold880 top.DUT.register\[7\]\[0\] vssd1 vssd1 vccd1 vccd1 net1996 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_686 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold891 top.DUT.register\[22\]\[12\] vssd1 vssd1 vccd1 vccd1 net2007 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_166_2929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11052_ net1184 net872 net836 top.ramstore\[3\] vssd1 vssd1 vccd1 vccd1 _01163_ sky130_fd_sc_hd__a22o_1
XANTENNA__06709__A2 net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10003_ net176 net1894 net626 vssd1 vssd1 vccd1 vccd1 _00208_ sky130_fd_sc_hd__mux2_1
XANTENNA_input21_A DAT_I[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07861__A _02999_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_199_3428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10698__S net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_204_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06590__B1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_2036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11954_ _05810_ _05774_ vssd1 vssd1 vccd1 vccd1 _05837_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_98_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_150_Left_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08867__C1 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07134__A2 net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10905_ net1307 net217 net479 vssd1 vssd1 vccd1 vccd1 _01066_ sky130_fd_sc_hd__mux2_1
X_11885_ _05730_ _05731_ _05751_ vssd1 vssd1 vccd1 vccd1 _05768_ sky130_fd_sc_hd__a21o_1
XFILLER_0_58_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13624_ clknet_leaf_75_clk _01211_ net1081 vssd1 vssd1 vccd1 vccd1 net50 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_184_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10836_ net1558 net212 net477 vssd1 vssd1 vccd1 vccd1 _00997_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_15_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13555_ clknet_leaf_105_clk _01142_ net969 vssd1 vssd1 vccd1 vccd1 top.ramload\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10767_ net2158 net245 net482 vssd1 vssd1 vccd1 vccd1 _00928_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12506_ clknet_leaf_79_clk _00098_ net1072 vssd1 vssd1 vccd1 vccd1 top.pc\[18\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__07842__B1 net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13486_ clknet_leaf_39_clk _01078_ net1055 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[30\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10698_ net1785 net265 net334 vssd1 vssd1 vccd1 vccd1 _00859_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12437_ clknet_leaf_87_clk _00033_ net1001 vssd1 vssd1 vccd1 vccd1 top.ramaddr\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_124_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08398__A1 net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_117_2198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12368_ clknet_leaf_103_clk top.ru.next_FetchedData\[12\] net974 vssd1 vssd1 vccd1
+ vccd1 top.a1.dataIn\[12\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_196_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11319_ top.a1.row2\[0\] net848 vssd1 vssd1 vccd1 vccd1 _05203_ sky130_fd_sc_hd__and2_1
XANTENNA__10462__A _04712_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12299_ top.pad.button_control.debounce top.pad.button_control.noisy vssd1 vssd1
+ vccd1 vccd1 _06110_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_130_2398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13546__Q top.ramload\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_180_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06860_ top.DUT.register\[10\]\[19\] net773 net729 top.DUT.register\[18\]\[19\] vssd1
+ vssd1 vccd1 vccd1 _01999_ sky130_fd_sc_hd__a22o_1
XANTENNA__07373__A2 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06791_ _01923_ _01925_ _01927_ _01929_ vssd1 vssd1 vccd1 vccd1 _01930_ sky130_fd_sc_hd__or4_4
XFILLER_0_179_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_42 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08530_ _02309_ _02386_ vssd1 vssd1 vccd1 vccd1 _03657_ sky130_fd_sc_hd__or2_1
XANTENNA__10401__S net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08461_ _02523_ _03566_ vssd1 vssd1 vccd1 vccd1 _03591_ sky130_fd_sc_hd__nor2_1
XANTENNA__08873__A2 net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07412_ top.DUT.register\[2\]\[9\] net742 net702 top.DUT.register\[3\]\[9\] _02550_
+ vssd1 vssd1 vccd1 vccd1 _02551_ sky130_fd_sc_hd__a221o_1
XFILLER_0_9_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08392_ _03393_ _03404_ net304 vssd1 vssd1 vccd1 vccd1 _03524_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_34_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_247 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_2508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07343_ top.DUT.register\[19\]\[8\] net536 net455 top.DUT.register\[25\]\[8\] _02481_
+ vssd1 vssd1 vccd1 vccd1 _02482_ sky130_fd_sc_hd__a221o_1
XFILLER_0_175_689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_174_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07274_ top.DUT.register\[1\]\[13\] net757 net720 top.DUT.register\[19\]\[13\] vssd1
+ vssd1 vccd1 vccd1 _02413_ sky130_fd_sc_hd__a22o_1
X_09013_ _03597_ _03620_ _03730_ _04087_ vssd1 vssd1 vccd1 vccd1 _04088_ sky130_fd_sc_hd__or4_1
X_06225_ net2314 net857 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedInstr\[19\] sky130_fd_sc_hd__and2_1
XFILLER_0_72_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1048_A net1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12185__A2 net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold110 top.a1.row1\[122\] vssd1 vssd1 vccd1 vccd1 net1226 sky130_fd_sc_hd__dlygate4sd3_1
X_06156_ top.a1.dataIn\[9\] vssd1 vssd1 vccd1 vccd1 _01399_ sky130_fd_sc_hd__inv_2
Xhold121 top.ramstore\[10\] vssd1 vssd1 vccd1 vccd1 net1237 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09050__A2 _03530_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold132 top.a1.row1\[8\] vssd1 vssd1 vccd1 vccd1 net1248 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_1_clk_A clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06939__A2 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold143 top.pad.button_control.noisy vssd1 vssd1 vccd1 vccd1 net1259 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_595 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold154 top.a1.row1\[1\] vssd1 vssd1 vccd1 vccd1 net1270 sky130_fd_sc_hd__dlygate4sd3_1
Xhold165 top.a1.row2\[32\] vssd1 vssd1 vccd1 vccd1 net1281 sky130_fd_sc_hd__dlygate4sd3_1
Xhold176 top.ramstore\[8\] vssd1 vssd1 vccd1 vccd1 net1292 sky130_fd_sc_hd__dlygate4sd3_1
Xhold187 top.a1.row2\[16\] vssd1 vssd1 vccd1 vccd1 net1303 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout601 _04965_ vssd1 vssd1 vccd1 vccd1 net601 sky130_fd_sc_hd__clkbuf_8
Xfanout612 _04955_ vssd1 vssd1 vccd1 vccd1 net612 sky130_fd_sc_hd__buf_6
Xhold198 top.DUT.register\[15\]\[13\] vssd1 vssd1 vccd1 vccd1 net1314 sky130_fd_sc_hd__dlygate4sd3_1
X_09915_ _04907_ _04920_ vssd1 vssd1 vccd1 vccd1 _04922_ sky130_fd_sc_hd__nor2_1
Xfanout623 net626 vssd1 vssd1 vccd1 vccd1 net623 sky130_fd_sc_hd__clkbuf_8
Xfanout634 _04714_ vssd1 vssd1 vccd1 vccd1 net634 sky130_fd_sc_hd__buf_4
XANTENNA_fanout296_X net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12360__Q top.a1.dataIn\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout675_A _01548_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout645 _01613_ vssd1 vssd1 vccd1 vccd1 net645 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_148_2659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout656 _01609_ vssd1 vssd1 vccd1 vccd1 net656 sky130_fd_sc_hd__clkbuf_4
Xfanout667 _01599_ vssd1 vssd1 vccd1 vccd1 net667 sky130_fd_sc_hd__buf_6
X_09846_ _01584_ net487 net401 top.a1.dataIn\[23\] net397 vssd1 vssd1 vccd1 vccd1
+ _04859_ sky130_fd_sc_hd__a221o_1
Xfanout678 _01548_ vssd1 vssd1 vccd1 vccd1 net678 sky130_fd_sc_hd__buf_4
Xfanout689 net690 vssd1 vssd1 vccd1 vccd1 net689 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_70_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07364__A2 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09777_ top.pc\[15\] _04403_ _04791_ vssd1 vssd1 vccd1 vccd1 _04797_ sky130_fd_sc_hd__a21o_1
XFILLER_0_197_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout463_X net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06989_ top.DUT.register\[13\]\[23\] net775 net755 top.DUT.register\[1\]\[23\] vssd1
+ vssd1 vccd1 vccd1 _02128_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_161_2859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08728_ net320 _03482_ vssd1 vssd1 vccd1 vccd1 _03846_ sky130_fd_sc_hd__nor2_1
XANTENNA__10311__S net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07116__A2 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_450 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08659_ _02048_ _03185_ _03264_ _03587_ _03779_ vssd1 vssd1 vccd1 vccd1 _03780_ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout630_X net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout728_X net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_205_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_194_3358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11670_ _05542_ _05548_ _05552_ _05547_ vssd1 vssd1 vccd1 vccd1 _05553_ sky130_fd_sc_hd__a22o_2
XFILLER_0_49_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10621_ net169 net1909 net346 vssd1 vssd1 vccd1 vccd1 _00786_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09813__A1 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_654 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_188 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13340_ clknet_leaf_130_clk _00932_ net910 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[26\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09895__X _04904_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10552_ net1485 net180 net354 vssd1 vssd1 vccd1 vccd1 _00719_ sky130_fd_sc_hd__mux2_1
XANTENNA__09120__B _02944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13271_ clknet_leaf_129_clk _00863_ net910 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[24\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_715 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10483_ net1678 net200 net363 vssd1 vssd1 vccd1 vccd1 _00653_ sky130_fd_sc_hd__mux2_1
X_12222_ top.lcd.cnt_20ms\[3\] _06051_ top.lcd.cnt_20ms\[4\] vssd1 vssd1 vccd1 vccd1
+ _06064_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09577__B1 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_595 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12153_ _06007_ _06034_ vssd1 vssd1 vccd1 vccd1 _06036_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_20_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08023__Y _03162_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11104_ _01405_ net1379 _01428_ _05057_ vssd1 vssd1 vccd1 vccd1 _01203_ sky130_fd_sc_hd__a31o_1
X_12084_ _05951_ _05964_ _05966_ vssd1 vssd1 vccd1 vccd1 _05967_ sky130_fd_sc_hd__or3_1
X_11035_ net15 net841 net818 top.ramload\[21\] vssd1 vssd1 vccd1 vccd1 _01147_ sky130_fd_sc_hd__a22o_1
XANTENNA__08552__A1 net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07355__A2 net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_704 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10221__S net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12986_ clknet_leaf_2_clk _00578_ net919 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[15\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07107__A2 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11937_ _05798_ _05813_ _05805_ vssd1 vssd1 vccd1 vccd1 _05820_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_129_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_156_111 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11868_ _05740_ _05748_ _05750_ vssd1 vssd1 vccd1 vccd1 _05751_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_129_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10819_ net161 net1535 net600 vssd1 vssd1 vccd1 vccd1 _00980_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_31_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13607_ clknet_leaf_89_clk _01194_ net1003 vssd1 vssd1 vccd1 vccd1 net62 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_156_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11799_ _05681_ vssd1 vssd1 vccd1 vccd1 _05682_ sky130_fd_sc_hd__inv_2
XANTENNA__09804__A1 _04151_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_2227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_119_2238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07815__B1 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13538_ clknet_leaf_92_clk _01125_ net995 vssd1 vssd1 vccd1 vccd1 top.a1.data\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_41_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13469_ clknet_leaf_13_clk _01061_ net953 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[30\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10891__S net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_2427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_140_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08791__A1 _03258_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07594__A2 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07961_ _03099_ vssd1 vssd1 vccd1 vccd1 _03100_ sky130_fd_sc_hd__inv_2
XFILLER_0_49_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09700_ _03430_ net404 net490 _04732_ vssd1 vssd1 vccd1 vccd1 _04733_ sky130_fd_sc_hd__o211a_1
XFILLER_0_208_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06912_ top.DUT.register\[18\]\[21\] net549 net537 top.DUT.register\[19\]\[21\] vssd1
+ vssd1 vccd1 vccd1 _02051_ sky130_fd_sc_hd__a22o_1
X_07892_ top.DUT.register\[15\]\[1\] net681 net677 top.DUT.register\[31\]\[1\] vssd1
+ vssd1 vccd1 vccd1 _03031_ sky130_fd_sc_hd__a22o_1
XANTENNA__07346__A2 net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09631_ _04164_ _04661_ _04671_ top.a1.state\[2\] vssd1 vssd1 vccd1 vccd1 _00114_
+ sky130_fd_sc_hd__a22o_1
X_06843_ _01975_ _01977_ _01979_ _01981_ vssd1 vssd1 vccd1 vccd1 _01982_ sky130_fd_sc_hd__or4_1
XANTENNA__06554__B1 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_179_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10131__S net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09562_ _04609_ _04610_ vssd1 vssd1 vccd1 vccd1 _04611_ sky130_fd_sc_hd__nand2_1
X_06774_ top.DUT.register\[28\]\[24\] net767 net720 top.DUT.register\[19\]\[24\] vssd1
+ vssd1 vccd1 vccd1 _01913_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_143_2589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08513_ _03060_ _03573_ _02390_ vssd1 vssd1 vccd1 vccd1 _03640_ sky130_fd_sc_hd__a21o_1
XFILLER_0_195_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09493_ _04544_ _04545_ vssd1 vssd1 vccd1 vccd1 _04546_ sky130_fd_sc_hd__nand2_1
XFILLER_0_148_612 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout256_A _04737_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_172_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_407 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08444_ _03572_ _03573_ vssd1 vssd1 vccd1 vccd1 _03574_ sky130_fd_sc_hd__and2_1
XFILLER_0_147_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_163_604 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_176_3088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08375_ net321 _03507_ _03495_ vssd1 vssd1 vccd1 vccd1 _03508_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout423_A net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07326_ top.DUT.register\[24\]\[12\] net643 net738 top.DUT.register\[12\]\[12\] _02464_
+ vssd1 vssd1 vccd1 vccd1 _02465_ sky130_fd_sc_hd__a221o_1
XFILLER_0_61_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_190_456 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07257_ top.DUT.register\[14\]\[13\] net585 net446 top.DUT.register\[1\]\[13\] _02395_
+ vssd1 vssd1 vccd1 vccd1 _02396_ sky130_fd_sc_hd__a221o_1
XFILLER_0_5_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06208_ top.ramload\[2\] net857 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedInstr\[2\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_103_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07188_ top.DUT.register\[9\]\[10\] net467 net523 top.DUT.register\[11\]\[10\] _02326_
+ vssd1 vssd1 vccd1 vccd1 _02327_ sky130_fd_sc_hd__a221o_1
XFILLER_0_60_178 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_197_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06139_ top.lcd.nextState\[0\] vssd1 vssd1 vccd1 vccd1 _01382_ sky130_fd_sc_hd__inv_2
XANTENNA__12545__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10306__S net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08642__A1_N net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout580_X net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout420 net421 vssd1 vssd1 vccd1 vccd1 net420 sky130_fd_sc_hd__buf_4
XANTENNA_fanout678_X net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout431 net433 vssd1 vssd1 vccd1 vccd1 net431 sky130_fd_sc_hd__clkbuf_4
Xfanout442 _01566_ vssd1 vssd1 vccd1 vccd1 net442 sky130_fd_sc_hd__clkbuf_4
Xfanout453 _01561_ vssd1 vssd1 vccd1 vccd1 net453 sky130_fd_sc_hd__buf_6
Xfanout464 net465 vssd1 vssd1 vccd1 vccd1 net464 sky130_fd_sc_hd__clkbuf_8
Xfanout475 net477 vssd1 vssd1 vccd1 vccd1 net475 sky130_fd_sc_hd__clkbuf_8
Xfanout486 net487 vssd1 vssd1 vccd1 vccd1 net486 sky130_fd_sc_hd__buf_2
XANTENNA__09731__B1 _04752_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout497 net498 vssd1 vssd1 vccd1 vccd1 net497 sky130_fd_sc_hd__clkbuf_4
X_09829_ top.pc\[21\] _04499_ vssd1 vssd1 vccd1 vccd1 _04844_ sky130_fd_sc_hd__or2_1
XANTENNA__06545__B1 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10041__S net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12840_ clknet_leaf_26_clk _00432_ net1011 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[10\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09115__B _03040_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08794__X _03909_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_567 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12771_ clknet_leaf_49_clk _00363_ net1061 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[8\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_96_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11722_ _05553_ _05581_ _05569_ _05566_ vssd1 vssd1 vccd1 vccd1 _05605_ sky130_fd_sc_hd__a211o_1
XFILLER_0_56_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_267 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12182__A2_N _05083_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11653_ _05509_ _05531_ _05508_ vssd1 vssd1 vccd1 vccd1 _05536_ sky130_fd_sc_hd__o21a_1
XFILLER_0_138_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_193_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10604_ net237 net2062 net347 vssd1 vssd1 vccd1 vccd1 _00769_ sky130_fd_sc_hd__mux2_1
X_11584_ _05441_ _05466_ vssd1 vssd1 vccd1 vccd1 _05467_ sky130_fd_sc_hd__nor2_2
XFILLER_0_119_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13323_ clknet_leaf_48_clk _00915_ net1069 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[25\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_91_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10535_ net1359 net254 net354 vssd1 vssd1 vccd1 vccd1 _00702_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13254_ clknet_leaf_38_clk _00846_ net1053 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[23\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_10466_ net1403 net261 net363 vssd1 vssd1 vccd1 vccd1 _00636_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_114_2157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12205_ top.lcd.cnt_20ms\[2\] top.lcd.cnt_20ms\[1\] top.lcd.cnt_20ms\[0\] vssd1 vssd1
+ vccd1 vccd1 _06051_ sky130_fd_sc_hd__and3_1
XFILLER_0_60_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10216__S net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13185_ clknet_leaf_16_clk _00777_ net960 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[21\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13428__RESET_B net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10397_ net1309 net144 _04982_ vssd1 vssd1 vccd1 vccd1 _00569_ sky130_fd_sc_hd__mux2_1
XANTENNA__07576__A2 net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12136_ _06014_ _06016_ _06018_ vssd1 vssd1 vccd1 vccd1 _06019_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_20_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06784__B1 net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12067_ _05940_ _05943_ _05948_ vssd1 vssd1 vccd1 vccd1 _05950_ sky130_fd_sc_hd__nor3_1
XANTENNA__06489__X _01628_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07328__A2 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11018_ net28 net840 _05044_ net1224 vssd1 vssd1 vccd1 vccd1 _01130_ sky130_fd_sc_hd__o22a_1
XANTENNA__11124__A3 net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_205_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06536__B1 net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_204_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_177_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10886__S net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12969_ clknet_leaf_51_clk _00561_ net1056 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[14\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_143_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06490_ net787 _01594_ _01611_ vssd1 vssd1 vccd1 vccd1 _01629_ sky130_fd_sc_hd__and3_4
XANTENNA__07500__A2 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_200_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09041__A _01790_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10187__A top.a1.instruction\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08160_ _03290_ _03291_ _03296_ net312 vssd1 vssd1 vccd1 vccd1 _03298_ sky130_fd_sc_hd__o22a_1
XFILLER_0_83_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_172_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_175 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07111_ top.DUT.register\[12\]\[16\] net739 _02246_ _02247_ _02249_ vssd1 vssd1 vccd1
+ vccd1 _02250_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_132_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_172_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08091_ _02724_ net332 vssd1 vssd1 vccd1 vccd1 _03230_ sky130_fd_sc_hd__or2_1
XFILLER_0_153_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12568__CLK clknet_leaf_128_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11060__A2 net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06671__Y _01810_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkload30 clknet_leaf_117_clk vssd1 vssd1 vccd1 vccd1 clkload30/Y sky130_fd_sc_hd__clkinv_8
Xclkload41 clknet_leaf_98_clk vssd1 vssd1 vccd1 vccd1 clkload41/Y sky130_fd_sc_hd__inv_16
X_07042_ top.DUT.register\[19\]\[22\] net536 net448 top.DUT.register\[21\]\[22\] _02180_
+ vssd1 vssd1 vccd1 vccd1 _02181_ sky130_fd_sc_hd__a221o_1
Xclkload52 clknet_leaf_87_clk vssd1 vssd1 vccd1 vccd1 clkload52/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload63 clknet_leaf_27_clk vssd1 vssd1 vccd1 vccd1 clkload63/Y sky130_fd_sc_hd__clkinv_2
Xclkload74 clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 clkload74/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_11_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload85 clknet_leaf_51_clk vssd1 vssd1 vccd1 vccd1 clkload85/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_113_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10126__S net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload96 clknet_leaf_73_clk vssd1 vssd1 vccd1 vccd1 clkload96/Y sky130_fd_sc_hd__inv_16
XANTENNA__07567__A2 net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07783__X _02922_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08993_ _04067_ _03799_ _04065_ vssd1 vssd1 vccd1 vccd1 _04068_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_54_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06775__B1 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07944_ _02070_ _02089_ vssd1 vssd1 vccd1 vccd1 _03083_ sky130_fd_sc_hd__and2_1
XFILLER_0_48_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_145_2618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07319__A2 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09713__B1 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07875_ top.DUT.register\[22\]\[1\] net649 net749 top.DUT.register\[17\]\[1\] vssd1
+ vssd1 vccd1 vccd1 _03014_ sky130_fd_sc_hd__a22o_1
XANTENNA__08120__A _03151_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06527__B1 net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_207_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout373_A _04981_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06826_ top.DUT.register\[16\]\[19\] net544 net537 top.DUT.register\[19\]\[19\] vssd1
+ vssd1 vccd1 vccd1 _01965_ sky130_fd_sc_hd__a22o_1
X_09614_ _01410_ _04657_ vssd1 vssd1 vccd1 vccd1 _04659_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_178_3117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_211_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09545_ net134 _04588_ _04593_ _04594_ vssd1 vssd1 vccd1 vccd1 _04595_ sky130_fd_sc_hd__o22ai_1
X_06757_ _01889_ _01891_ _01893_ _01895_ vssd1 vssd1 vccd1 vccd1 _01896_ sky130_fd_sc_hd__or4_4
XANTENNA__10796__S net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_129_clk clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_129_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_69_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout540_A _01540_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08819__A2 top.pc\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout638_A _01629_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_195_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_174_Right_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09476_ _01585_ _02111_ vssd1 vssd1 vccd1 vccd1 _04530_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_191_3306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06688_ top.DUT.register\[21\]\[26\] net658 net646 top.DUT.register\[24\]\[26\] _01826_
+ vssd1 vssd1 vccd1 vccd1 _01827_ sky130_fd_sc_hd__a221o_1
XANTENNA__08119__X _03258_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12296__B net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_191_3317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_535 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08427_ _03222_ net280 _03255_ net283 vssd1 vssd1 vccd1 vccd1 _03558_ sky130_fd_sc_hd__o22a_1
XFILLER_0_163_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1070_X net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout426_X net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_202_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_451 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10528__C net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08358_ _03342_ _03490_ vssd1 vssd1 vccd1 vccd1 _03491_ sky130_fd_sc_hd__nor2_1
Xclkload2 clknet_4_6__leaf_clk vssd1 vssd1 vccd1 vccd1 clkload2/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_18_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_190_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07309_ top.DUT.register\[19\]\[12\] net535 net519 top.DUT.register\[10\]\[12\] vssd1
+ vssd1 vccd1 vccd1 _02448_ sky130_fd_sc_hd__a22o_1
XANTENNA__11051__A2 net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08452__B1 _03580_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08289_ _03416_ _03421_ _03424_ vssd1 vssd1 vccd1 vccd1 _03425_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_210_3601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_190_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_150_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10320_ net172 net2252 net383 vssd1 vssd1 vccd1 vccd1 _00497_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout795_X net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_189_3279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10251_ net192 net1919 net391 vssd1 vssd1 vccd1 vccd1 _00430_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_375 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10036__S net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07558__A2 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10182_ _04709_ _04947_ _04958_ vssd1 vssd1 vccd1 vccd1 _04962_ sky130_fd_sc_hd__and3_4
XANTENNA__06766__B1 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout250 _05439_ vssd1 vssd1 vccd1 vccd1 net250 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_TAPCELL_ROW_208_3563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08507__A1 _03263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11106__A3 net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout261 net262 vssd1 vssd1 vccd1 vccd1 net261 sky130_fd_sc_hd__buf_2
XFILLER_0_205_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout283 _03171_ vssd1 vssd1 vccd1 vccd1 net283 sky130_fd_sc_hd__clkbuf_4
Xfanout294 net295 vssd1 vssd1 vccd1 vccd1 net294 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09180__A1 net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09413__X _04471_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07730__A2 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12823_ clknet_leaf_2_clk _00415_ net914 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[10\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_2_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_141_Right_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12754_ clknet_leaf_26_clk _00346_ net1014 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[8\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_535 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_395 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11705_ _05550_ _05586_ vssd1 vssd1 vccd1 vccd1 _05588_ sky130_fd_sc_hd__or2_1
XFILLER_0_127_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12685_ clknet_leaf_44_clk _00277_ net1062 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[5\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11290__A2 _05128_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11636_ _05487_ _05511_ _05516_ vssd1 vssd1 vccd1 vccd1 _05519_ sky130_fd_sc_hd__or3_1
XFILLER_0_37_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09235__A2 _02502_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11567_ _05448_ _05449_ vssd1 vssd1 vccd1 vccd1 _05450_ sky130_fd_sc_hd__nor2_1
XFILLER_0_21_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07797__A2 net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13306_ clknet_leaf_4_clk _00898_ net939 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[25\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_10518_ net1627 net182 net360 vssd1 vssd1 vccd1 vccd1 _00687_ sky130_fd_sc_hd__mux2_1
Xhold709 top.DUT.register\[31\]\[0\] vssd1 vssd1 vccd1 vccd1 net1825 sky130_fd_sc_hd__dlygate4sd3_1
X_11498_ _05349_ net273 vssd1 vssd1 vccd1 vccd1 _05381_ sky130_fd_sc_hd__nand2_1
X_13237_ clknet_leaf_32_clk _00829_ net1044 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[23\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10449_ net184 net1685 net366 vssd1 vssd1 vccd1 vccd1 _00620_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07549__A2 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13168_ clknet_leaf_28_clk _00760_ net1011 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[20\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_41_clk_A clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12119_ top.a1.dataIn\[2\] _05982_ _06000_ _05997_ _05996_ vssd1 vssd1 vccd1 vccd1
+ _06002_ sky130_fd_sc_hd__o311a_1
X_13099_ clknet_leaf_50_clk _00691_ net1059 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[18\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_127_2348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06509__B1 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_205_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06379__B top.a1.instruction\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07660_ _02798_ vssd1 vssd1 vccd1 vccd1 _02799_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_0_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_56_clk_A clknet_4_12__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06611_ top.DUT.register\[22\]\[27\] net577 net562 top.DUT.register\[2\]\[27\] vssd1
+ vssd1 vccd1 vccd1 _01750_ sky130_fd_sc_hd__a22o_1
XANTENNA__09323__X _04386_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07721__A2 net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_204_173 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07591_ top.DUT.register\[15\]\[6\] net706 net698 top.DUT.register\[31\]\[6\] vssd1
+ vssd1 vccd1 vccd1 _02730_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_140_2548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09330_ net132 _04384_ _04392_ net810 vssd1 vssd1 vccd1 vccd1 _04393_ sky130_fd_sc_hd__o22a_1
X_06542_ top.DUT.register\[21\]\[29\] net657 net724 top.DUT.register\[29\]\[29\] vssd1
+ vssd1 vccd1 vccd1 _01681_ sky130_fd_sc_hd__a22o_1
XFILLER_0_87_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09474__A2 _04514_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09261_ top.pc\[11\] _04310_ vssd1 vssd1 vccd1 vccd1 _04327_ sky130_fd_sc_hd__nor2_1
X_06473_ net788 _01594_ _01611_ vssd1 vssd1 vccd1 vccd1 _01612_ sky130_fd_sc_hd__and3_4
XFILLER_0_118_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_173_3036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_173_3047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_440 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08212_ net322 _03349_ _03299_ vssd1 vssd1 vccd1 vccd1 _03350_ sky130_fd_sc_hd__o21a_1
XFILLER_0_145_434 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09754__A2_N _04752_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09192_ _04261_ _04262_ vssd1 vssd1 vccd1 vccd1 _04263_ sky130_fd_sc_hd__nand2_1
XFILLER_0_173_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_114_clk_A clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08143_ _02329_ net328 vssd1 vssd1 vccd1 vccd1 _03281_ sky130_fd_sc_hd__nand2_1
XFILLER_0_31_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07788__A2 net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08074_ _03212_ vssd1 vssd1 vccd1 vccd1 _03213_ sky130_fd_sc_hd__inv_2
XFILLER_0_113_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07025_ top.DUT.register\[4\]\[20\] net670 net764 top.DUT.register\[9\]\[20\] _02163_
+ vssd1 vssd1 vccd1 vccd1 _02164_ sky130_fd_sc_hd__a221o_1
XFILLER_0_113_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_141_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_129_clk_A clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08402__X _03534_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout490_A net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold14 top.ramstore\[24\] vssd1 vssd1 vccd1 vccd1 net1130 sky130_fd_sc_hd__dlygate4sd3_1
X_08976_ net890 _01393_ vssd1 vssd1 vccd1 vccd1 _04051_ sky130_fd_sc_hd__nand2_2
Xhold25 top.a1.data\[3\] vssd1 vssd1 vccd1 vccd1 net1141 sky130_fd_sc_hd__dlygate4sd3_1
Xhold36 top.ramstore\[21\] vssd1 vssd1 vccd1 vccd1 net1152 sky130_fd_sc_hd__dlygate4sd3_1
Xhold47 _01185_ vssd1 vssd1 vccd1 vccd1 net1163 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11195__B net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold58 _01182_ vssd1 vssd1 vccd1 vccd1 net1174 sky130_fd_sc_hd__dlygate4sd3_1
X_07927_ _02329_ _02385_ vssd1 vssd1 vccd1 vccd1 _03066_ sky130_fd_sc_hd__nand2b_1
Xhold69 _01163_ vssd1 vssd1 vccd1 vccd1 net1185 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout376_X net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout755_A _01620_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09162__A1 net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07960__Y _03099_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07858_ net820 net410 _02949_ vssd1 vssd1 vccd1 vccd1 _02997_ sky130_fd_sc_hd__and3_1
XFILLER_0_98_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07173__B1 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06809_ top.DUT.register\[7\]\[17\] net659 net747 top.DUT.register\[17\]\[17\] _01947_
+ vssd1 vssd1 vccd1 vccd1 _01948_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout922_A net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout543_X net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07789_ top.DUT.register\[14\]\[2\] net583 net567 top.DUT.register\[6\]\[2\] vssd1
+ vssd1 vccd1 vccd1 _02928_ sky130_fd_sc_hd__a22o_1
XFILLER_0_210_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_203_3493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09528_ _01810_ _04577_ vssd1 vssd1 vccd1 vccd1 _04579_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_158_2809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout710_X net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09459_ net822 _02360_ net422 vssd1 vssd1 vccd1 vccd1 _04514_ sky130_fd_sc_hd__a21o_4
XTAP_TAPCELL_ROW_80_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08673__B1 net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_176_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08009__B top.a1.instruction\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12470_ clknet_leaf_82_clk _00065_ net993 vssd1 vssd1 vccd1 vccd1 top.ramstore\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_108_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11421_ _05259_ _05288_ vssd1 vssd1 vccd1 vccd1 _05304_ sky130_fd_sc_hd__or2_2
XFILLER_0_117_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07779__A2 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11352_ _05228_ _05229_ _05232_ _05233_ vssd1 vssd1 vccd1 vccd1 _05235_ sky130_fd_sc_hd__a211o_1
XFILLER_0_34_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08025__A _01589_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06987__B1 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10303_ net245 top.DUT.register\[12\]\[7\] net381 vssd1 vssd1 vccd1 vccd1 _00480_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_111_2105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_684 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_18_Left_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11283_ top.a1.row1\[115\] _05132_ _05146_ top.a1.row2\[43\] _05172_ vssd1 vssd1
+ vccd1 vccd1 _05173_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_95_1871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_2116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13022_ clknet_leaf_18_clk _00614_ net1029 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[16\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_10234_ net255 top.DUT.register\[10\]\[4\] net390 vssd1 vssd1 vccd1 vccd1 _00413_
+ sky130_fd_sc_hd__mux2_1
Xfanout1001 net1005 vssd1 vssd1 vccd1 vccd1 net1001 sky130_fd_sc_hd__clkbuf_4
Xfanout1012 net1016 vssd1 vssd1 vccd1 vccd1 net1012 sky130_fd_sc_hd__clkbuf_4
X_10165_ net1561 net185 net604 vssd1 vssd1 vccd1 vccd1 _00364_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_7_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1023 net1025 vssd1 vssd1 vccd1 vccd1 net1023 sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_210_Right_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08031__Y _03170_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1034 net1036 vssd1 vssd1 vccd1 vccd1 net1034 sky130_fd_sc_hd__clkbuf_2
Xfanout1045 net1048 vssd1 vssd1 vccd1 vccd1 net1045 sky130_fd_sc_hd__clkbuf_4
Xfanout1056 net1058 vssd1 vssd1 vccd1 vccd1 net1056 sky130_fd_sc_hd__clkbuf_4
Xfanout1067 net1068 vssd1 vssd1 vccd1 vccd1 net1067 sky130_fd_sc_hd__buf_2
X_10096_ net2174 net223 net612 vssd1 vssd1 vccd1 vccd1 _00297_ sky130_fd_sc_hd__mux2_1
Xfanout1078 net1079 vssd1 vssd1 vccd1 vccd1 net1078 sky130_fd_sc_hd__clkbuf_4
Xfanout1089 net1096 vssd1 vssd1 vccd1 vccd1 net1089 sky130_fd_sc_hd__buf_2
XFILLER_0_107_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_109_2078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07703__A2 net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12806_ clknet_leaf_33_clk _00398_ net1046 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[9\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_122_2278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13786_ clknet_leaf_68_clk _01355_ vssd1 vssd1 vccd1 vccd1 top.pad.button_control.r_counter\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_186_367 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10998_ net1172 _05032_ net589 vssd1 vssd1 vccd1 vccd1 _01122_ sky130_fd_sc_hd__mux2_1
XFILLER_0_202_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12737_ clknet_leaf_18_clk _00329_ net1026 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[7\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_516 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12668_ clknet_leaf_130_clk _00260_ net909 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[5\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_154_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11619_ net234 _05476_ top.a1.dataIn\[13\] vssd1 vssd1 vccd1 vccd1 _05502_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11015__A2 net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13443__RESET_B net1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12599_ clknet_leaf_2_clk _00191_ net918 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[3\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_13_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_170_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold506 top.DUT.register\[23\]\[21\] vssd1 vssd1 vccd1 vccd1 net1622 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06978__B1 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold517 top.DUT.register\[13\]\[9\] vssd1 vssd1 vccd1 vccd1 net1633 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold528 top.DUT.register\[26\]\[3\] vssd1 vssd1 vccd1 vccd1 net1644 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold539 top.DUT.register\[26\]\[17\] vssd1 vssd1 vccd1 vccd1 net1655 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_51_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08830_ _03370_ _03922_ vssd1 vssd1 vccd1 vccd1 _03943_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_51_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_max_cap606_X net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07942__A2 _02242_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08761_ _03796_ _03875_ net313 vssd1 vssd1 vccd1 vccd1 _03877_ sky130_fd_sc_hd__mux2_1
X_07712_ net326 _02849_ vssd1 vssd1 vccd1 vccd1 _02851_ sky130_fd_sc_hd__nand2_1
X_08692_ _02179_ _03810_ vssd1 vssd1 vccd1 vccd1 _03811_ sky130_fd_sc_hd__nand2b_1
XANTENNA__07155__B1 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09695__A2 net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07643_ top.DUT.register\[20\]\[5\] net663 net655 top.DUT.register\[21\]\[5\] _02781_
+ vssd1 vssd1 vccd1 vccd1 _02782_ sky130_fd_sc_hd__a221o_1
XFILLER_0_79_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_183 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07574_ _02706_ _02708_ _02710_ _02712_ vssd1 vssd1 vccd1 vccd1 _02713_ sky130_fd_sc_hd__or4_4
XTAP_TAPCELL_ROW_24_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09313_ net897 top.pc\[13\] _04376_ net889 vssd1 vssd1 vccd1 vccd1 _00093_ sky130_fd_sc_hd__o211a_1
X_06525_ top.DUT.register\[16\]\[29\] net544 net505 top.DUT.register\[27\]\[29\] vssd1
+ vssd1 vccd1 vccd1 _01664_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_196_Left_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_192_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout336_A net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_192_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_60_clk clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_60_clk
+ sky130_fd_sc_hd__clkbuf_8
X_09244_ top.pc\[9\] _04284_ top.pc\[10\] vssd1 vssd1 vccd1 vccd1 _04311_ sky130_fd_sc_hd__a21oi_1
X_06456_ top.a1.instruction\[23\] _01593_ vssd1 vssd1 vccd1 vccd1 _01595_ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_62_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09175_ _02773_ _02777_ vssd1 vssd1 vccd1 vccd1 _04247_ sky130_fd_sc_hd__nand2_1
XANTENNA__06681__A2 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_153_2739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_hold1186_A top.a1.row2\[35\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06387_ top.DUT.register\[9\]\[30\] net468 net569 top.DUT.register\[6\]\[30\] vssd1
+ vssd1 vccd1 vccd1 _01526_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout503_A _01567_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08126_ _03180_ _03181_ _03183_ _03262_ vssd1 vssd1 vccd1 vccd1 _03265_ sky130_fd_sc_hd__a31o_1
XFILLER_0_160_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06969__B1 net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12363__Q top.a1.dataIn\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_1_Right_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08057_ _03195_ vssd1 vssd1 vccd1 vccd1 _03196_ sky130_fd_sc_hd__inv_2
XFILLER_0_114_684 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_186_3238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07008_ top.DUT.register\[22\]\[20\] net577 net534 top.DUT.register\[12\]\[20\] vssd1
+ vssd1 vccd1 vccd1 _02147_ sky130_fd_sc_hd__a22o_1
Xoutput48 net48 vssd1 vssd1 vccd1 vccd1 ADR_O[17] sky130_fd_sc_hd__buf_2
XANTENNA_fanout872_A _01427_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout493_X net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput59 net59 vssd1 vssd1 vccd1 vccd1 ADR_O[27] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_168_2960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10314__S net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_168_2971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07394__B1 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_205_3522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08959_ top.ramstore\[15\] net877 _02609_ net693 vssd1 vssd1 vccd1 vccd1 _00065_
+ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout660_X net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout758_X net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11970_ _05846_ _05849_ _05825_ vssd1 vssd1 vccd1 vccd1 _05853_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_168_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10921_ net1376 net268 net591 vssd1 vssd1 vccd1 vccd1 _01082_ sky130_fd_sc_hd__mux2_1
XFILLER_0_169_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_196_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10852_ net1837 net156 net476 vssd1 vssd1 vccd1 vccd1 _01013_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13640_ clknet_leaf_93_clk _01226_ net994 vssd1 vssd1 vccd1 vccd1 top.busy_o sky130_fd_sc_hd__dfrtp_1
XFILLER_0_168_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_630 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13571_ clknet_leaf_89_clk _01158_ net1002 vssd1 vssd1 vccd1 vccd1 net110 sky130_fd_sc_hd__dfrtp_1
X_10783_ net1807 net178 net484 vssd1 vssd1 vccd1 vccd1 _00944_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_51_clk clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_51_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_66_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12522_ clknet_leaf_88_clk _00114_ net1004 vssd1 vssd1 vccd1 vccd1 top.a1.state\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_136_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_590 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_1900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06672__A2 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12453_ clknet_leaf_75_clk _00049_ net1083 vssd1 vssd1 vccd1 vccd1 top.ramaddr\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_152_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11404_ _05277_ _05282_ _05286_ _05279_ vssd1 vssd1 vccd1 vccd1 _05287_ sky130_fd_sc_hd__a22o_2
XANTENNA__08949__B2 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12384_ clknet_leaf_110_clk top.ru.next_FetchedData\[28\] net989 vssd1 vssd1 vccd1
+ vccd1 top.a1.dataIn\[28\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_10_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11335_ _05214_ _05215_ _05217_ _05210_ vssd1 vssd1 vccd1 vccd1 _05218_ sky130_fd_sc_hd__a31oi_4
XANTENNA__06424__A2 net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11266_ top.a1.row1\[113\] _05132_ _05146_ top.a1.row2\[41\] _05154_ vssd1 vssd1
+ vccd1 vccd1 _05158_ sky130_fd_sc_hd__a221o_1
X_13005_ clknet_leaf_44_clk _00597_ net1063 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[15\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_10217_ net201 net2165 net395 vssd1 vssd1 vccd1 vccd1 _00397_ sky130_fd_sc_hd__mux2_1
XANTENNA__10224__S net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11197_ _04664_ _05004_ _05018_ vssd1 vssd1 vccd1 vccd1 _05105_ sky130_fd_sc_hd__and3_1
XFILLER_0_94_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09771__A1_N net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10148_ net1492 net264 net602 vssd1 vssd1 vccd1 vccd1 _00347_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_402 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_124_2307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10079_ net689 _04947_ _04952_ vssd1 vssd1 vccd1 vccd1 _04955_ sky130_fd_sc_hd__and3_4
XANTENNA__09314__A top.pc\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_202_441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10894__S net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13769_ clknet_leaf_100_clk _01340_ vssd1 vssd1 vccd1 vccd1 top.lcd.cnt_500hz\[5\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_42_clk clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_42_clk
+ sky130_fd_sc_hd__clkbuf_8
X_06310_ _01462_ _01465_ vssd1 vssd1 vccd1 vccd1 _01466_ sky130_fd_sc_hd__xor2_1
XFILLER_0_155_540 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07290_ net807 _02428_ net437 vssd1 vssd1 vccd1 vccd1 _02429_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_143_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06241_ top.ramload\[2\] net855 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedData\[2\]
+ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_44_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_415 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06663__A2 net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_519 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06172_ top.a1.halfData\[5\] _01413_ vssd1 vssd1 vccd1 vccd1 _01414_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_135_2469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold303 top.DUT.register\[23\]\[31\] vssd1 vssd1 vccd1 vccd1 net1419 sky130_fd_sc_hd__dlygate4sd3_1
Xhold314 top.DUT.register\[15\]\[24\] vssd1 vssd1 vccd1 vccd1 net1430 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold325 top.DUT.register\[15\]\[8\] vssd1 vssd1 vccd1 vccd1 net1441 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold336 top.DUT.register\[1\]\[5\] vssd1 vssd1 vccd1 vccd1 net1452 sky130_fd_sc_hd__dlygate4sd3_1
Xhold347 top.DUT.register\[2\]\[7\] vssd1 vssd1 vccd1 vccd1 net1463 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold358 top.DUT.register\[6\]\[23\] vssd1 vssd1 vccd1 vccd1 net1474 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_4_3__f_clk clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_3__leaf_clk sky130_fd_sc_hd__clkbuf_16
Xhold369 top.DUT.register\[19\]\[22\] vssd1 vssd1 vccd1 vccd1 net1485 sky130_fd_sc_hd__dlygate4sd3_1
X_09931_ net798 _04934_ _04935_ _04936_ vssd1 vssd1 vccd1 vccd1 _04937_ sky130_fd_sc_hd__a211o_1
Xfanout805 net806 vssd1 vssd1 vccd1 vccd1 net805 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_68_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12577__RESET_B net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout816 net817 vssd1 vssd1 vccd1 vccd1 net816 sky130_fd_sc_hd__buf_2
XANTENNA__09365__A1 net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_7__f_clk_A clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09365__B2 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10134__S net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09862_ top.a1.instruction\[24\] net486 net401 top.a1.dataIn\[24\] net398 vssd1 vssd1
+ vccd1 vccd1 _04874_ sky130_fd_sc_hd__a221o_1
Xfanout827 net828 vssd1 vssd1 vccd1 vccd1 net827 sky130_fd_sc_hd__clkbuf_4
Xfanout838 net839 vssd1 vssd1 vccd1 vccd1 net838 sky130_fd_sc_hd__buf_2
XANTENNA__09739__A1_N net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout849 net851 vssd1 vssd1 vccd1 vccd1 net849 sky130_fd_sc_hd__buf_2
XANTENNA__09923__S net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1003 top.DUT.register\[8\]\[27\] vssd1 vssd1 vccd1 vccd1 net2119 sky130_fd_sc_hd__dlygate4sd3_1
X_08813_ _01878_ _03090_ vssd1 vssd1 vccd1 vccd1 _03927_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_181_3157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1014 top.DUT.register\[15\]\[27\] vssd1 vssd1 vccd1 vccd1 net2130 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_181_3168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09793_ net827 _04430_ _04811_ vssd1 vssd1 vccd1 vccd1 _04812_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_30_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1025 top.DUT.register\[15\]\[7\] vssd1 vssd1 vccd1 vccd1 net2141 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout286_A _03170_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1036 top.DUT.register\[1\]\[20\] vssd1 vssd1 vccd1 vccd1 net2152 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1047 top.DUT.register\[1\]\[27\] vssd1 vssd1 vccd1 vccd1 net2163 sky130_fd_sc_hd__dlygate4sd3_1
X_08744_ _03504_ _03534_ _03689_ net279 _03860_ vssd1 vssd1 vccd1 vccd1 _03861_ sky130_fd_sc_hd__o221a_1
Xhold1058 top.DUT.register\[6\]\[16\] vssd1 vssd1 vccd1 vccd1 net2174 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1069 top.DUT.register\[10\]\[11\] vssd1 vssd1 vccd1 vccd1 net2185 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_163_2890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08675_ _03307_ _03311_ vssd1 vssd1 vccd1 vccd1 _03795_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout453_A _01561_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_200_3441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_200_3452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07626_ top.DUT.register\[12\]\[5\] net532 net503 top.DUT.register\[27\]\[5\] vssd1
+ vssd1 vccd1 vccd1 _02765_ sky130_fd_sc_hd__a22o_1
XFILLER_0_177_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_37_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_490 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12358__Q top.a1.dataIn\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_192_101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07557_ top.DUT.register\[10\]\[7\] net770 net730 top.DUT.register\[14\]\[7\] vssd1
+ vssd1 vccd1 vccd1 _02696_ sky130_fd_sc_hd__a22o_1
XANTENNA__09878__B _04577_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout620_A net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_33_clk clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_33_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout718_A _01635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout339_X net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06508_ top.DUT.register\[30\]\[30\] net760 net744 top.DUT.register\[2\]\[30\] vssd1
+ vssd1 vccd1 vccd1 _01647_ sky130_fd_sc_hd__a22o_1
XFILLER_0_91_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06583__A _01721_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07488_ top.DUT.register\[21\]\[14\] net448 net440 top.DUT.register\[5\]\[14\] _02626_
+ vssd1 vssd1 vccd1 vccd1 _02627_ sky130_fd_sc_hd__a221o_1
XANTENNA__07300__B1 net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06654__A2 net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06439_ _01388_ net896 _01390_ _01502_ vssd1 vssd1 vccd1 vccd1 _01578_ sky130_fd_sc_hd__and4_1
X_09227_ net139 _04286_ _04295_ vssd1 vssd1 vccd1 vccd1 _04296_ sky130_fd_sc_hd__o21ai_1
XANTENNA__10309__S net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout506_X net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12188__B1 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_79_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09158_ _04216_ _04219_ _04230_ vssd1 vssd1 vccd1 vccd1 _04231_ sky130_fd_sc_hd__and3_1
XANTENNA__09894__A net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10738__A1 net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08109_ _02329_ net299 vssd1 vssd1 vccd1 vccd1 _03248_ sky130_fd_sc_hd__nand2_1
XFILLER_0_133_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09089_ top.a1.instruction\[3\] _01502_ _04160_ _04163_ vssd1 vssd1 vccd1 vccd1 _04164_
+ sky130_fd_sc_hd__and4_2
XFILLER_0_102_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11120_ net906 net1294 net861 _05065_ vssd1 vssd1 vccd1 vccd1 _01211_ sky130_fd_sc_hd__a31o_1
XANTENNA__08948__A1_N _02827_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_1830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold870 top.DUT.register\[27\]\[20\] vssd1 vssd1 vccd1 vccd1 net1986 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout875_X net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold881 top.DUT.register\[9\]\[21\] vssd1 vssd1 vccd1 vccd1 net1997 sky130_fd_sc_hd__dlygate4sd3_1
X_11051_ net1210 net866 net837 top.ramstore\[2\] vssd1 vssd1 vccd1 vccd1 _01162_ sky130_fd_sc_hd__a22o_1
Xhold892 top.DUT.register\[23\]\[8\] vssd1 vssd1 vccd1 vccd1 net2008 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10044__S net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07367__B1 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10002_ net180 net1610 net623 vssd1 vssd1 vccd1 vccd1 _00207_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_199_3429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08449__S net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07119__B1 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06758__A _01887_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09134__A top.pc\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_2037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input14_A DAT_I[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11953_ _05755_ _05834_ _05795_ _05833_ vssd1 vssd1 vccd1 vccd1 _05836_ sky130_fd_sc_hd__nor4b_1
XFILLER_0_98_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_169_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10904_ net1939 net223 net479 vssd1 vssd1 vccd1 vccd1 _01065_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11884_ _05722_ _05763_ vssd1 vssd1 vccd1 vccd1 _05767_ sky130_fd_sc_hd__xor2_1
XFILLER_0_168_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13623_ clknet_leaf_73_clk _01210_ net1078 vssd1 vssd1 vccd1 vccd1 net49 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_211_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08619__B1 _03736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06893__A2 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10835_ net1440 net221 net474 vssd1 vssd1 vccd1 vccd1 _00996_ sky130_fd_sc_hd__mux2_1
XANTENNA__09788__B _04438_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_24_clk clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_24_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_15_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13554_ clknet_leaf_104_clk _01141_ net969 vssd1 vssd1 vccd1 vccd1 top.ramload\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_183_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_307 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10766_ net1500 net243 net482 vssd1 vssd1 vccd1 vccd1 _00927_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10977__A1 top.a1.dataIn\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12505_ clknet_leaf_81_clk _00097_ net993 vssd1 vssd1 vccd1 vccd1 top.pc\[17\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_164_381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13485_ clknet_leaf_43_clk _01077_ net1062 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[30\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_180_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10219__S net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10697_ net2044 net270 net335 vssd1 vssd1 vccd1 vccd1 _00858_ sky130_fd_sc_hd__mux2_1
XANTENNA__12179__B1 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12436_ clknet_leaf_87_clk _00032_ net1004 vssd1 vssd1 vccd1 vccd1 top.ramaddr\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_112_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_117_2199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09595__A1 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12367_ clknet_leaf_104_clk top.ru.next_FetchedData\[11\] net973 vssd1 vssd1 vccd1
+ vccd1 top.a1.dataIn\[11\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_1_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07070__A2 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11318_ net1084 net813 _05202_ _05201_ vssd1 vssd1 vccd1 vccd1 _01272_ sky130_fd_sc_hd__a31o_1
X_12298_ net904 net118 _06108_ net2268 vssd1 vssd1 vccd1 vccd1 _01351_ sky130_fd_sc_hd__a22o_1
XANTENNA__08213__A _03258_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09347__A1 net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11249_ net878 net880 _01382_ _05118_ vssd1 vssd1 vccd1 vccd1 _05142_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_130_2399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10889__S net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06790_ top.DUT.register\[21\]\[17\] net448 net504 top.DUT.register\[27\]\[17\] _01928_
+ vssd1 vssd1 vccd1 vccd1 _01929_ sky130_fd_sc_hd__a221o_1
XFILLER_0_145_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_179_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_4_11__f_clk clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_11__leaf_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__13805__RESET_B net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13562__Q top.ramload\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08460_ net430 _03585_ _03589_ net426 vssd1 vssd1 vccd1 vccd1 _03590_ sky130_fd_sc_hd__a22o_1
XANTENNA__09979__A net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_203_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07530__B1 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08873__A3 _03440_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_175_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07411_ top.DUT.register\[13\]\[9\] net774 net726 top.DUT.register\[18\]\[9\] vssd1
+ vssd1 vccd1 vccd1 _02550_ sky130_fd_sc_hd__a22o_1
XFILLER_0_175_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_46_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08391_ _03522_ vssd1 vssd1 vccd1 vccd1 _03523_ sky130_fd_sc_hd__inv_2
XFILLER_0_147_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06884__A2 net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_15_clk clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_15_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_9_259 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07342_ top.DUT.register\[14\]\[8\] net584 net466 top.DUT.register\[13\]\[8\] vssd1
+ vssd1 vccd1 vccd1 _02481_ sky130_fd_sc_hd__a22o_1
XFILLER_0_190_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_162_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10968__A1 top.a1.dataIn\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06636__A2 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07273_ top.DUT.register\[15\]\[13\] net708 net700 top.DUT.register\[31\]\[13\] vssd1
+ vssd1 vccd1 vccd1 _02412_ sky130_fd_sc_hd__a22o_1
XANTENNA__10129__S net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_699 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09012_ _03520_ _03550_ _03574_ _04086_ vssd1 vssd1 vccd1 vccd1 _04087_ sky130_fd_sc_hd__or4b_1
X_06224_ net1706 net856 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedInstr\[18\] sky130_fd_sc_hd__and2_1
XANTENNA__07786__X _02925_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold100 top.DUT.register\[26\]\[14\] vssd1 vssd1 vccd1 vccd1 net1216 sky130_fd_sc_hd__dlygate4sd3_1
X_06155_ top.a1.dataIn\[11\] vssd1 vssd1 vccd1 vccd1 _01398_ sky130_fd_sc_hd__inv_2
XFILLER_0_78_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout201_A _04841_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold111 top.lcd.cnt_20ms\[12\] vssd1 vssd1 vccd1 vccd1 net1227 sky130_fd_sc_hd__dlygate4sd3_1
Xhold122 top.a1.row2\[18\] vssd1 vssd1 vccd1 vccd1 net1238 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07597__B1 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold133 top.a1.row1\[2\] vssd1 vssd1 vccd1 vccd1 net1249 sky130_fd_sc_hd__dlygate4sd3_1
Xhold144 top.DUT.register\[8\]\[17\] vssd1 vssd1 vccd1 vccd1 net1260 sky130_fd_sc_hd__dlygate4sd3_1
Xhold155 top.a1.row2\[3\] vssd1 vssd1 vccd1 vccd1 net1271 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07061__A2 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold166 top.ramload\[1\] vssd1 vssd1 vccd1 vccd1 net1282 sky130_fd_sc_hd__dlygate4sd3_1
Xhold177 _01168_ vssd1 vssd1 vccd1 vccd1 net1293 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold188 top.ramaddr\[21\] vssd1 vssd1 vccd1 vccd1 net1304 sky130_fd_sc_hd__dlygate4sd3_1
Xhold199 top.DUT.register\[30\]\[21\] vssd1 vssd1 vccd1 vccd1 net1315 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout602 _04957_ vssd1 vssd1 vccd1 vccd1 net602 sky130_fd_sc_hd__buf_6
X_09914_ _04907_ _04920_ vssd1 vssd1 vccd1 vccd1 _04921_ sky130_fd_sc_hd__nand2_1
Xfanout613 _04955_ vssd1 vssd1 vccd1 vccd1 net613 sky130_fd_sc_hd__buf_8
XFILLER_0_0_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07349__B1 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout624 net626 vssd1 vssd1 vccd1 vccd1 net624 sky130_fd_sc_hd__clkbuf_8
Xfanout635 _01629_ vssd1 vssd1 vccd1 vccd1 net635 sky130_fd_sc_hd__clkbuf_8
Xfanout646 _01613_ vssd1 vssd1 vccd1 vccd1 net646 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07962__A _01659_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input6_A DAT_I[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09845_ net2102 net180 net632 vssd1 vssd1 vccd1 vccd1 _00143_ sky130_fd_sc_hd__mux2_1
Xfanout657 _01609_ vssd1 vssd1 vccd1 vccd1 net657 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout570_A _01525_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10799__S net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout668 _01599_ vssd1 vssd1 vccd1 vccd1 net668 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout191_X net191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout679 _01547_ vssd1 vssd1 vccd1 vccd1 net679 sky130_fd_sc_hd__buf_4
XANTENNA_fanout668_A _01599_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09776_ net1431 net189 net632 vssd1 vssd1 vccd1 vccd1 _00136_ sky130_fd_sc_hd__mux2_1
X_06988_ top.DUT.register\[6\]\[23\] net636 net719 top.DUT.register\[19\]\[23\] _02126_
+ vssd1 vssd1 vccd1 vccd1 _02127_ sky130_fd_sc_hd__a221o_1
XFILLER_0_198_738 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08727_ net318 _03472_ vssd1 vssd1 vccd1 vccd1 _03845_ sky130_fd_sc_hd__nor2_1
XANTENNA__08849__B1 _03185_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout456_X net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_205_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08658_ _02047_ net502 vssd1 vssd1 vccd1 vccd1 _03779_ sky130_fd_sc_hd__nand2_1
XFILLER_0_178_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07521__B1 net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07609_ _02740_ _02747_ vssd1 vssd1 vccd1 vccd1 _02748_ sky130_fd_sc_hd__or2_4
XTAP_TAPCELL_ROW_194_3359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_495 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06875__A2 net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout623_X net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08589_ _02614_ net494 _03711_ net428 _03712_ vssd1 vssd1 vccd1 vccd1 _03713_ sky130_fd_sc_hd__a221o_1
X_10620_ net172 net2215 net348 vssd1 vssd1 vccd1 vccd1 _00785_ sky130_fd_sc_hd__mux2_1
XFILLER_0_165_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_12_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07202__A net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06627__A2 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10551_ net1635 net194 net355 vssd1 vssd1 vccd1 vccd1 _00718_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10039__S net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_180_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10482_ net1497 net185 net363 vssd1 vssd1 vccd1 vccd1 _00652_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_198 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13270_ clknet_leaf_13_clk _00862_ net943 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[24\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12499__RESET_B net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12221_ _06059_ _06063_ net980 vssd1 vssd1 vccd1 vccd1 _01314_ sky130_fd_sc_hd__o21a_1
XANTENNA__07856__B _02994_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07588__A0 _02679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12152_ _06033_ _06029_ _06030_ vssd1 vssd1 vccd1 vccd1 _06035_ sky130_fd_sc_hd__mux2_1
XANTENNA__09129__A net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07052__A2 net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11103_ net42 net864 vssd1 vssd1 vccd1 vccd1 _05057_ sky130_fd_sc_hd__and2_1
X_12083_ _05953_ _05955_ vssd1 vssd1 vccd1 vccd1 _05966_ sky130_fd_sc_hd__xnor2_1
X_11034_ net14 net838 net816 net2309 vssd1 vssd1 vccd1 vccd1 _01146_ sky130_fd_sc_hd__o22a_1
XPHY_EDGE_ROW_188_Right_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10502__S net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_189_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_204_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12985_ clknet_leaf_15_clk _00577_ net959 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[15\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_115_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11936_ _05817_ _05818_ vssd1 vssd1 vccd1 vccd1 _05819_ sky130_fd_sc_hd__nand2_1
XFILLER_0_197_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_156_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11867_ _05716_ _05749_ vssd1 vssd1 vccd1 vccd1 _05750_ sky130_fd_sc_hd__and2_1
XFILLER_0_86_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_31_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13606_ clknet_leaf_73_clk _01193_ net1078 vssd1 vssd1 vccd1 vccd1 net51 sky130_fd_sc_hd__dfrtp_1
X_10818_ net164 net1554 net600 vssd1 vssd1 vccd1 vccd1 _00979_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_31_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11798_ _05653_ _05679_ vssd1 vssd1 vccd1 vccd1 _05681_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_55_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_2228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06618__A2 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13537_ clknet_leaf_93_clk _01124_ net995 vssd1 vssd1 vccd1 vccd1 top.a1.data\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_10749_ net1570 net192 net420 vssd1 vssd1 vccd1 vccd1 _00910_ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_41_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09738__S net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06951__A _02069_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13468_ clknet_leaf_129_clk _01060_ net910 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[30\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_180_671 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_658 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_132_2428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12419_ clknet_leaf_110_clk top.ru.next_FetchedInstr\[31\] net989 vssd1 vssd1 vccd1
+ vccd1 top.a1.instruction\[31\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__07579__B1 net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13399_ clknet_leaf_129_clk _00991_ net911 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[28\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_140_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07043__A2 net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08791__A2 _03260_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07960_ _01679_ _01698_ _03098_ vssd1 vssd1 vccd1 vccd1 _03099_ sky130_fd_sc_hd__a21oi_2
Xclkbuf_leaf_4_clk clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_4_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_56_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06911_ _01964_ _02007_ _02049_ vssd1 vssd1 vccd1 vccd1 _02050_ sky130_fd_sc_hd__nand3_1
XANTENNA__08230__X _03367_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07891_ _03023_ _03025_ _03027_ _03029_ vssd1 vssd1 vccd1 vccd1 _03030_ sky130_fd_sc_hd__or4_4
XPHY_EDGE_ROW_155_Right_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09630_ _04659_ _04672_ _04670_ top.a1.state\[1\] vssd1 vssd1 vccd1 vccd1 _00113_
+ sky130_fd_sc_hd__o2bb2a_1
X_06842_ top.DUT.register\[20\]\[19\] net565 net441 top.DUT.register\[5\]\[19\] _01980_
+ vssd1 vssd1 vccd1 vccd1 _01981_ sky130_fd_sc_hd__a221o_1
XANTENNA__10412__S net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07751__B1 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_99 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09561_ _04591_ _04593_ _04608_ _01505_ vssd1 vssd1 vccd1 vccd1 _04610_ sky130_fd_sc_hd__o31a_1
X_06773_ top.DUT.register\[21\]\[24\] net657 net649 top.DUT.register\[22\]\[24\] _01911_
+ vssd1 vssd1 vccd1 vccd1 _01912_ sky130_fd_sc_hd__a221o_1
X_08512_ net1379 net833 net803 _03639_ vssd1 vssd1 vccd1 vccd1 _00029_ sky130_fd_sc_hd__a22o_1
X_09492_ _01887_ _01896_ _04543_ vssd1 vssd1 vccd1 vccd1 _04545_ sky130_fd_sc_hd__or3_1
XANTENNA__07503__B1 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_624 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06857__A2 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08443_ _02571_ _03571_ vssd1 vssd1 vccd1 vccd1 _03573_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout151_A _04938_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_419 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08374_ net316 _03498_ _03497_ vssd1 vssd1 vccd1 vccd1 _03507_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_176_3089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07325_ top.DUT.register\[30\]\[12\] net758 net710 top.DUT.register\[11\]\[12\] vssd1
+ vssd1 vccd1 vccd1 _02464_ sky130_fd_sc_hd__a22o_1
XANTENNA__06609__A2 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1060_A net1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07256_ top.DUT.register\[8\]\[13\] net541 net510 top.DUT.register\[4\]\[13\] vssd1
+ vssd1 vccd1 vccd1 _02395_ sky130_fd_sc_hd__a22o_1
XFILLER_0_171_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06207_ net1282 net859 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedInstr\[1\] sky130_fd_sc_hd__and2_1
XFILLER_0_116_598 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_170_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07187_ top.DUT.register\[22\]\[10\] net575 net571 top.DUT.register\[23\]\[10\] vssd1
+ vssd1 vccd1 vccd1 _02326_ sky130_fd_sc_hd__a22o_1
XANTENNA__08124__Y _03263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06138_ net881 vssd1 vssd1 vccd1 vccd1 _01381_ sky130_fd_sc_hd__inv_2
XANTENNA__07034__A2 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_73 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12371__Q top.a1.dataIn\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11118__A1 net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout410 net411 vssd1 vssd1 vccd1 vccd1 net410 sky130_fd_sc_hd__buf_2
Xfanout421 _04961_ vssd1 vssd1 vccd1 vccd1 net421 sky130_fd_sc_hd__clkbuf_8
XANTENNA__07990__B1 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout432 net433 vssd1 vssd1 vccd1 vccd1 net432 sky130_fd_sc_hd__clkbuf_2
Xfanout443 _01564_ vssd1 vssd1 vccd1 vccd1 net443 sky130_fd_sc_hd__clkbuf_8
Xfanout454 _01561_ vssd1 vssd1 vccd1 vccd1 net454 sky130_fd_sc_hd__buf_4
XANTENNA_fanout952_A net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout573_X net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout465 net466 vssd1 vssd1 vccd1 vccd1 net465 sky130_fd_sc_hd__clkbuf_8
Xfanout476 net477 vssd1 vssd1 vccd1 vccd1 net476 sky130_fd_sc_hd__buf_4
XANTENNA__10322__S net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout487 _04776_ vssd1 vssd1 vccd1 vccd1 net487 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09731__B2 top.a1.dataIn\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09828_ top.pc\[21\] _04499_ vssd1 vssd1 vccd1 vccd1 _04843_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_122_Right_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout498 _03335_ vssd1 vssd1 vccd1 vccd1 net498 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07742__B1 net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout740_X net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09759_ net826 _04379_ _04752_ top.a1.dataIn\[14\] vssd1 vssd1 vccd1 vccd1 _04781_
+ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_87_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_179_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12770_ clknet_leaf_25_clk _00362_ net1012 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[8\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_139_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_139_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11721_ _05553_ _05581_ _05566_ vssd1 vssd1 vccd1 vccd1 _05604_ sky130_fd_sc_hd__a21oi_1
XANTENNA__06848__A2 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_279 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_599 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_471 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11652_ _05533_ _05534_ vssd1 vssd1 vccd1 vccd1 _05535_ sky130_fd_sc_hd__nand2_1
XFILLER_0_83_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08028__A _03152_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10603_ net248 net2085 net346 vssd1 vssd1 vccd1 vccd1 _00768_ sky130_fd_sc_hd__mux2_1
XANTENNA__11054__B1 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09798__A1 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11583_ _05430_ net249 _05415_ vssd1 vssd1 vccd1 vccd1 _05466_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_135_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13322_ clknet_leaf_115_clk _00914_ net963 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[25\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_134_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10534_ net2114 net257 net355 vssd1 vssd1 vccd1 vccd1 _00701_ sky130_fd_sc_hd__mux2_1
XANTENNA__07273__A2 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08470__B2 net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13253_ clknet_leaf_33_clk _00845_ net1044 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[23\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_10465_ net1533 net266 net361 vssd1 vssd1 vccd1 vccd1 _00635_ sky130_fd_sc_hd__mux2_1
XANTENNA__07586__B net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_114_2158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12204_ _05968_ net688 _06050_ vssd1 vssd1 vccd1 vccd1 _01310_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07025__A2 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10396_ _04153_ _04155_ _04708_ net399 vssd1 vssd1 vccd1 vccd1 _04984_ sky130_fd_sc_hd__nand4_2
XFILLER_0_20_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13184_ clknet_leaf_113_clk _00776_ net991 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[21\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_12135_ _05994_ _06002_ _06012_ _05998_ vssd1 vssd1 vccd1 vccd1 _06018_ sky130_fd_sc_hd__a22o_1
X_12066_ _05943_ _05948_ vssd1 vssd1 vccd1 vccd1 _05949_ sky130_fd_sc_hd__nor2_1
X_11017_ net27 net842 net819 net1284 vssd1 vssd1 vccd1 vccd1 _01129_ sky130_fd_sc_hd__a22o_1
XANTENNA__10232__S net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13818__1103 vssd1 vssd1 vccd1 vccd1 _13818__1103/HI net1103 sky130_fd_sc_hd__conb_1
XFILLER_0_189_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07733__B1 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_204_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_579 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12968_ clknet_leaf_27_clk _00560_ net1008 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[14\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_176_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_0_clk_A clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06839__A2 net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11919_ _05758_ _05778_ _05787_ _05767_ vssd1 vssd1 vccd1 vccd1 _05802_ sky130_fd_sc_hd__a31o_1
XFILLER_0_59_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12899_ clknet_leaf_53_clk _00491_ net1038 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[12\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10187__B top.a1.instruction\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07110_ top.DUT.register\[22\]\[16\] net648 net640 top.DUT.register\[8\]\[16\] _02248_
+ vssd1 vssd1 vccd1 vccd1 _02249_ sky130_fd_sc_hd__a221o_1
XFILLER_0_27_187 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08090_ net291 _03177_ _03228_ net304 vssd1 vssd1 vccd1 vccd1 _03229_ sky130_fd_sc_hd__a31o_1
XFILLER_0_43_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07264__A2 net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload20 clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 clkload20/Y sky130_fd_sc_hd__bufinv_16
X_07041_ top.DUT.register\[14\]\[22\] net583 net543 top.DUT.register\[16\]\[22\] vssd1
+ vssd1 vccd1 vccd1 _02180_ sky130_fd_sc_hd__a22o_1
Xclkload31 clknet_leaf_103_clk vssd1 vssd1 vccd1 vccd1 clkload31/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_2_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload42 clknet_leaf_99_clk vssd1 vssd1 vccd1 vccd1 clkload42/Y sky130_fd_sc_hd__clkinv_2
XFILLER_0_70_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13295__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload53 clknet_leaf_88_clk vssd1 vssd1 vccd1 vccd1 clkload53/Y sky130_fd_sc_hd__inv_6
Xclkload64 clknet_leaf_28_clk vssd1 vssd1 vccd1 vccd1 clkload64/Y sky130_fd_sc_hd__clkinv_4
Xclkload75 clknet_leaf_36_clk vssd1 vssd1 vccd1 vccd1 clkload75/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_140_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkload86 clknet_leaf_17_clk vssd1 vssd1 vccd1 vccd1 clkload86/Y sky130_fd_sc_hd__clkinv_2
Xclkload97 clknet_leaf_74_clk vssd1 vssd1 vccd1 vccd1 clkload97/Y sky130_fd_sc_hd__inv_12
XFILLER_0_140_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08992_ _03736_ _03759_ _03777_ vssd1 vssd1 vccd1 vccd1 _04067_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_54_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_76 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07943_ _02199_ _02219_ vssd1 vssd1 vccd1 vccd1 _03082_ sky130_fd_sc_hd__and2_1
XANTENNA__08401__A net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_145_2619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09713__A1 top.a1.dataIn\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout199_A _04788_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10142__S net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07874_ top.DUT.register\[4\]\[1\] net669 _03001_ _03012_ vssd1 vssd1 vccd1 vccd1
+ _03013_ sky130_fd_sc_hd__a211o_1
X_09613_ top.a1.halfData\[3\] _01385_ _01411_ top.a1.halfData\[5\] vssd1 vssd1 vccd1
+ vccd1 _04658_ sky130_fd_sc_hd__or4bb_4
XANTENNA__07017__A _02155_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_207_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06825_ _01962_ _01963_ vssd1 vssd1 vccd1 vccd1 _01964_ sky130_fd_sc_hd__or2_2
XANTENNA_fanout366_A net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_178_3118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_211_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09544_ _04578_ _04582_ _04592_ net812 vssd1 vssd1 vccd1 vccd1 _04594_ sky130_fd_sc_hd__a31o_1
X_06756_ top.DUT.register\[11\]\[24\] net526 net454 top.DUT.register\[29\]\[24\] _01894_
+ vssd1 vssd1 vccd1 vccd1 _01895_ sky130_fd_sc_hd__a221o_1
XFILLER_0_78_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07304__X _02443_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06687_ top.DUT.register\[7\]\[26\] net661 net650 top.DUT.register\[22\]\[26\] vssd1
+ vssd1 vccd1 vccd1 _01826_ sky130_fd_sc_hd__a22o_1
XFILLER_0_93_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09475_ _01585_ _02111_ vssd1 vssd1 vccd1 vccd1 _04529_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout533_A _01542_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_191_3307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_191_3318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08426_ net434 _03556_ vssd1 vssd1 vccd1 vccd1 _03557_ sky130_fd_sc_hd__nor2_1
XFILLER_0_93_547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12366__Q top.a1.dataIn\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_202_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_463 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout700_A _01643_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08357_ _02754_ _03054_ vssd1 vssd1 vccd1 vccd1 _03490_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_117_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout419_X net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload3 clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 clkload3/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_190_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07308_ top.DUT.register\[30\]\[12\] net579 net439 top.DUT.register\[5\]\[12\] _02446_
+ vssd1 vssd1 vccd1 vccd1 _02447_ sky130_fd_sc_hd__a221o_1
XFILLER_0_116_351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07255__A2 net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08452__B2 net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08288_ _03342_ _03414_ _03423_ net496 vssd1 vssd1 vccd1 vccd1 _03424_ sky130_fd_sc_hd__o22a_1
XFILLER_0_144_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_210_3602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10317__S net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07239_ top.DUT.register\[24\]\[10\] net643 net635 top.DUT.register\[6\]\[10\] _02377_
+ vssd1 vssd1 vccd1 vccd1 _02378_ sky130_fd_sc_hd__a221o_1
X_10250_ net202 net1930 net391 vssd1 vssd1 vccd1 vccd1 _00429_ sky130_fd_sc_hd__mux2_1
XANTENNA__07007__A2 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout690_X net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10181_ net689 _04959_ vssd1 vssd1 vccd1 vccd1 _04961_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_208_3564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout251 _04741_ vssd1 vssd1 vccd1 vccd1 net251 sky130_fd_sc_hd__buf_2
Xfanout262 _04733_ vssd1 vssd1 vccd1 vccd1 net262 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08507__A2 _03623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout273 _05357_ vssd1 vssd1 vccd1 vccd1 net273 sky130_fd_sc_hd__buf_2
XANTENNA__10052__S net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout284 _03170_ vssd1 vssd1 vccd1 vccd1 net284 sky130_fd_sc_hd__clkbuf_4
Xfanout295 _03020_ vssd1 vssd1 vccd1 vccd1 net295 sky130_fd_sc_hd__buf_2
XANTENNA__06469__C _01607_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_202_826 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11672__A top.a1.dataIn\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12822_ clknet_leaf_13_clk _00414_ net941 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[10\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_2_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11275__B1 _05149_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12753_ clknet_leaf_111_clk _00345_ net988 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[8\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_96_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06485__B _01607_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08029__Y _03168_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11704_ _05550_ _05583_ vssd1 vssd1 vccd1 vccd1 _05587_ sky130_fd_sc_hd__xor2_2
XFILLER_0_166_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12684_ clknet_leaf_62_clk _00276_ net1093 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[5\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_167_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_194_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11635_ _05511_ _05516_ vssd1 vssd1 vccd1 vccd1 _05518_ sky130_fd_sc_hd__nor2_1
XFILLER_0_112_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12443__RESET_B net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11566_ _05418_ net250 _01397_ vssd1 vssd1 vccd1 vccd1 _05449_ sky130_fd_sc_hd__and3b_1
XFILLER_0_135_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13305_ clknet_leaf_14_clk _00897_ net956 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[25\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_10517_ net2012 net195 net359 vssd1 vssd1 vccd1 vccd1 _00686_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10227__S net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11497_ _05375_ _05379_ vssd1 vssd1 vccd1 vccd1 _05380_ sky130_fd_sc_hd__nand2_1
XFILLER_0_122_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13236_ clknet_leaf_58_clk _00828_ net1076 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[23\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_10448_ net205 net2052 net366 vssd1 vssd1 vccd1 vccd1 _00619_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11847__A top.a1.dataIn\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13167_ clknet_leaf_51_clk _00759_ net1035 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[20\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_209_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10379_ net2283 net215 net374 vssd1 vssd1 vccd1 vccd1 _00554_ sky130_fd_sc_hd__mux2_1
XFILLER_0_209_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12118_ top.a1.dataIn\[2\] _05982_ _06000_ vssd1 vssd1 vccd1 vccd1 _06001_ sky130_fd_sc_hd__nor3_1
X_13098_ clknet_leaf_115_clk _00690_ net963 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[18\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_12049_ _05919_ _05929_ _05913_ vssd1 vssd1 vccd1 vccd1 _05932_ sky130_fd_sc_hd__nor3b_2
XFILLER_0_137_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07706__B1 net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_2349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10897__S net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_204_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06610_ top.DUT.register\[13\]\[27\] net464 net554 top.DUT.register\[3\]\[27\] _01748_
+ vssd1 vssd1 vccd1 vccd1 _01749_ sky130_fd_sc_hd__a221o_1
XFILLER_0_177_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07590_ _02728_ vssd1 vssd1 vccd1 vccd1 _02729_ sky130_fd_sc_hd__inv_2
XFILLER_0_204_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_140_2549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_34 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06541_ top.DUT.register\[14\]\[29\] net732 net728 top.DUT.register\[18\]\[29\] vssd1
+ vssd1 vccd1 vccd1 _01680_ sky130_fd_sc_hd__a22o_1
XANTENNA__09052__A _03645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13570__Q top.ramload\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06472_ top.a1.instruction\[20\] top.a1.instruction\[21\] net792 vssd1 vssd1 vccd1
+ vccd1 _01611_ sky130_fd_sc_hd__and3b_2
XFILLER_0_62_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09260_ top.pc\[11\] _04310_ vssd1 vssd1 vccd1 vccd1 _04326_ sky130_fd_sc_hd__and2_1
XANTENNA__08682__A1 _03263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07485__A2 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_173_3037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08211_ _03314_ _03348_ net316 vssd1 vssd1 vccd1 vccd1 _03349_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_173_3048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11018__B1 _05044_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_452 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09191_ _02723_ _02728_ vssd1 vssd1 vccd1 vccd1 _04262_ sky130_fd_sc_hd__nand2_1
XFILLER_0_145_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11569__B2 top.a1.dataIn\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08142_ _02544_ net301 vssd1 vssd1 vccd1 vccd1 _03280_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_155_2770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08073_ _03208_ _03211_ net291 vssd1 vssd1 vccd1 vccd1 _03212_ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10137__S net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07024_ top.DUT.register\[22\]\[20\] net650 net761 top.DUT.register\[30\]\[20\] vssd1
+ vssd1 vccd1 vccd1 _02163_ sky130_fd_sc_hd__a22o_1
XFILLER_0_101_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_141_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10661__A _04155_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1023_A net1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07945__B1 _02156_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08975_ _03141_ net691 net1149 net874 vssd1 vssd1 vccd1 vccd1 _00081_ sky130_fd_sc_hd__a2bb2o_1
Xhold15 _01184_ vssd1 vssd1 vccd1 vccd1 net1131 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout483_A _04962_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_184_3199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold26 top.a1.data\[0\] vssd1 vssd1 vccd1 vccd1 net1142 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09147__C1 net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold37 _01181_ vssd1 vssd1 vccd1 vccd1 net1153 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_194_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07926_ _03064_ vssd1 vssd1 vccd1 vccd1 _03065_ sky130_fd_sc_hd__inv_2
Xhold48 top.a1.data\[5\] vssd1 vssd1 vccd1 vccd1 net1164 sky130_fd_sc_hd__dlygate4sd3_1
Xhold59 top.a1.row1\[112\] vssd1 vssd1 vccd1 vccd1 net1175 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09698__B1 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09100__C_N _04172_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout650_A _01612_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07857_ _02974_ _02994_ vssd1 vssd1 vccd1 vccd1 _02996_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout748_A net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout369_X net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06808_ top.DUT.register\[10\]\[17\] net771 net738 top.DUT.register\[12\]\[17\] vssd1
+ vssd1 vccd1 vccd1 _01947_ sky130_fd_sc_hd__a22o_1
XANTENNA__10600__S net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07788_ top.DUT.register\[9\]\[2\] net467 net535 top.DUT.register\[19\]\[2\] _02926_
+ vssd1 vssd1 vccd1 vccd1 _02927_ sky130_fd_sc_hd__a221o_1
XFILLER_0_211_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_203_3494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09527_ _01810_ _04577_ vssd1 vssd1 vccd1 vccd1 _04578_ sky130_fd_sc_hd__nand2_1
X_06739_ _01877_ vssd1 vssd1 vccd1 vccd1 _01878_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout915_A net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08122__B1 _03256_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout536_X net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07476__A2 net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09458_ _04509_ _04512_ vssd1 vssd1 vccd1 vccd1 _04513_ sky130_fd_sc_hd__xnor2_1
X_08409_ _03474_ _03540_ net288 vssd1 vssd1 vccd1 vccd1 _03541_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07688__Y _02827_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10395__X _04983_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout703_X net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09389_ top.pc\[18\] _04438_ vssd1 vssd1 vccd1 vccd1 _04448_ sky130_fd_sc_hd__and2_1
XFILLER_0_163_254 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11420_ _05259_ _05288_ vssd1 vssd1 vccd1 vccd1 _05303_ sky130_fd_sc_hd__nand2_1
XFILLER_0_151_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07228__A2 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13817__1102 vssd1 vssd1 vccd1 vccd1 _13817__1102/HI net1102 sky130_fd_sc_hd__conb_1
XFILLER_0_105_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11351_ _05232_ _05233_ vssd1 vssd1 vccd1 vccd1 _05234_ sky130_fd_sc_hd__or2_1
XANTENNA__10047__S net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08025__B _03152_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09836__S net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10302_ net242 net1813 net381 vssd1 vssd1 vccd1 vccd1 _00479_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_111_2106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11282_ top.a1.row2\[27\] _05142_ _05150_ top.a1.row1\[107\] vssd1 vssd1 vccd1 vccd1
+ _05172_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_111_2117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_1872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13021_ clknet_leaf_3_clk _00613_ net920 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[16\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09386__C1 net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10233_ net261 net1695 net390 vssd1 vssd1 vccd1 vccd1 _00412_ sky130_fd_sc_hd__mux2_1
X_10164_ net1434 net204 net605 vssd1 vssd1 vccd1 vccd1 _00363_ sky130_fd_sc_hd__mux2_1
Xfanout1002 net1005 vssd1 vssd1 vccd1 vccd1 net1002 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_7_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07400__A2 net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1013 net1016 vssd1 vssd1 vccd1 vccd1 net1013 sky130_fd_sc_hd__buf_2
XFILLER_0_100_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1024 net1025 vssd1 vssd1 vccd1 vccd1 net1024 sky130_fd_sc_hd__clkbuf_2
Xfanout1035 net1036 vssd1 vssd1 vccd1 vccd1 net1035 sky130_fd_sc_hd__clkbuf_4
Xfanout1046 net1048 vssd1 vssd1 vccd1 vccd1 net1046 sky130_fd_sc_hd__clkbuf_4
Xfanout1057 net1058 vssd1 vssd1 vccd1 vccd1 net1057 sky130_fd_sc_hd__clkbuf_4
X_10095_ net2214 net189 net611 vssd1 vssd1 vccd1 vccd1 _00296_ sky130_fd_sc_hd__mux2_1
Xfanout1068 net1069 vssd1 vssd1 vccd1 vccd1 net1068 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08976__A net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1079 net1087 vssd1 vssd1 vccd1 vccd1 net1079 sky130_fd_sc_hd__buf_2
XFILLER_0_107_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_109_2079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09143__Y _04217_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10510__S net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12805_ clknet_leaf_35_clk _00397_ net1040 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[9\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13785_ clknet_leaf_68_clk _01354_ vssd1 vssd1 vccd1 vccd1 top.pad.button_control.r_counter\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_10997_ net843 _05030_ _05031_ net849 top.a1.dataIn\[8\] vssd1 vssd1 vccd1 vccd1
+ _05032_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_122_2279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_379 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12736_ clknet_leaf_114_clk _00328_ net992 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[7\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07467__A2 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06675__B1 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12667_ clknet_leaf_119_clk _00259_ net931 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[5\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_72_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_182_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11618_ _05450_ _05477_ _05499_ _05500_ vssd1 vssd1 vccd1 vccd1 _05501_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__08416__A1 net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_182_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_170_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12598_ clknet_leaf_3_clk _00190_ net940 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[3\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11549_ _05425_ _05429_ _05431_ vssd1 vssd1 vccd1 vccd1 _05432_ sky130_fd_sc_hd__a21o_1
Xhold507 top.DUT.register\[17\]\[31\] vssd1 vssd1 vccd1 vccd1 net1623 sky130_fd_sc_hd__dlygate4sd3_1
Xhold518 top.DUT.register\[3\]\[17\] vssd1 vssd1 vccd1 vccd1 net1634 sky130_fd_sc_hd__dlygate4sd3_1
Xhold529 top.DUT.register\[22\]\[1\] vssd1 vssd1 vccd1 vccd1 net1645 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13219_ clknet_leaf_54_clk _00811_ net1037 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[22\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_51_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13565__Q top.ramload\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08760_ _03875_ vssd1 vssd1 vccd1 vccd1 _03876_ sky130_fd_sc_hd__inv_2
X_07711_ net326 _02849_ vssd1 vssd1 vccd1 vccd1 _02850_ sky130_fd_sc_hd__nor2_1
X_08691_ _03770_ _03809_ _02005_ vssd1 vssd1 vccd1 vccd1 _03810_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_73_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07642_ top.DUT.register\[28\]\[5\] net766 net750 top.DUT.register\[26\]\[5\] vssd1
+ vssd1 vccd1 vccd1 _02781_ sky130_fd_sc_hd__a22o_1
XANTENNA__10420__S net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_177_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07573_ top.DUT.register\[13\]\[6\] net463 net515 top.DUT.register\[7\]\[6\] _02711_
+ vssd1 vssd1 vccd1 vccd1 _02712_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_66_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12365__RESET_B net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09312_ net136 _04362_ _04375_ vssd1 vssd1 vccd1 vccd1 _04376_ sky130_fd_sc_hd__o21ai_1
X_06524_ top.DUT.register\[19\]\[29\] net537 net449 top.DUT.register\[21\]\[29\] _01662_
+ vssd1 vssd1 vccd1 vccd1 _01663_ sky130_fd_sc_hd__a221o_1
XFILLER_0_48_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08655__A1 net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07458__A2 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08655__B2 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09510__A _01854_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06666__B1 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09243_ top.pc\[9\] top.pc\[10\] _04284_ vssd1 vssd1 vccd1 vccd1 _04310_ sky130_fd_sc_hd__and3_1
XFILLER_0_63_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06455_ top.a1.instruction\[23\] _01593_ vssd1 vssd1 vccd1 vccd1 _01594_ sky130_fd_sc_hd__nor2_2
XANTENNA_fanout329_A net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_173_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06386_ net683 _01512_ _01516_ vssd1 vssd1 vccd1 vccd1 _01525_ sky130_fd_sc_hd__and3_4
X_09174_ _02773_ _02777_ vssd1 vssd1 vccd1 vccd1 _04246_ sky130_fd_sc_hd__or2_1
XANTENNA__06418__B1 net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08125_ _03160_ _03181_ vssd1 vssd1 vccd1 vccd1 _03264_ sky130_fd_sc_hd__or2_2
XFILLER_0_31_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07091__B1 net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08056_ _03192_ _03194_ net277 vssd1 vssd1 vccd1 vccd1 _03195_ sky130_fd_sc_hd__mux2_1
XANTENNA__07630__A2 net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_186_3239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout698_A _01643_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07007_ top.DUT.register\[15\]\[20\] net682 net678 top.DUT.register\[31\]\[20\] vssd1
+ vssd1 vccd1 vccd1 _02146_ sky130_fd_sc_hd__a22o_1
XFILLER_0_3_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput49 net49 vssd1 vssd1 vccd1 vccd1 ADR_O[18] sky130_fd_sc_hd__buf_2
XFILLER_0_101_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_168_2961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_168_2972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout865_A net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_208_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08958_ _02652_ net691 net1143 net874 vssd1 vssd1 vccd1 vccd1 _00064_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_90_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_205_3523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07909_ net314 _02944_ _03047_ vssd1 vssd1 vccd1 vccd1 _03048_ sky130_fd_sc_hd__a21o_1
X_08889_ net279 _03838_ _03994_ _03998_ vssd1 vssd1 vccd1 vccd1 _03999_ sky130_fd_sc_hd__o211ai_2
XANTENNA_fanout653_X net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10920_ net1825 net144 _04960_ vssd1 vssd1 vccd1 vccd1 _01081_ sky130_fd_sc_hd__mux2_1
XANTENNA__10330__S net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07697__A2 net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08894__B2 net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12850__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10851_ net1530 net159 net476 vssd1 vssd1 vccd1 vccd1 _01012_ sky130_fd_sc_hd__mux2_1
X_13570_ clknet_leaf_104_clk _01157_ net972 vssd1 vssd1 vccd1 vccd1 top.ramload\[31\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__07449__A2 net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10782_ net2037 net183 net483 vssd1 vssd1 vccd1 vccd1 _00943_ sky130_fd_sc_hd__mux2_1
XFILLER_0_149_582 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06657__B1 net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12521_ clknet_leaf_88_clk _00113_ net1005 vssd1 vssd1 vccd1 vccd1 top.a1.state\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_136_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_40_clk_A clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_1901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12452_ clknet_leaf_75_clk _00048_ net1080 vssd1 vssd1 vccd1 vccd1 top.ramaddr\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_152_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11403_ _05277_ _05281_ _05285_ vssd1 vssd1 vccd1 vccd1 _05286_ sky130_fd_sc_hd__nand3_1
XANTENNA__08949__A2 net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12383_ clknet_leaf_109_clk top.ru.next_FetchedData\[27\] net977 vssd1 vssd1 vccd1
+ vccd1 top.a1.dataIn\[27\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_105_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11334_ _05206_ _05216_ vssd1 vssd1 vccd1 vccd1 _05217_ sky130_fd_sc_hd__nand2_1
XANTENNA__07621__A2 net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_55_clk_A clknet_4_12__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11265_ top.a1.row1\[57\] _05136_ _05139_ top.a1.row2\[9\] net815 vssd1 vssd1 vccd1
+ vccd1 _05157_ sky130_fd_sc_hd__a221o_1
XANTENNA__10505__S net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13004_ clknet_leaf_64_clk _00596_ net1095 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[15\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_10216_ net184 net1940 net395 vssd1 vssd1 vccd1 vccd1 _00396_ sky130_fd_sc_hd__mux2_1
X_11196_ top.a1.state\[1\] top.a1.state\[2\] _05084_ vssd1 vssd1 vccd1 vccd1 _05104_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_118_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10147_ net1582 net268 net604 vssd1 vssd1 vccd1 vccd1 _00346_ sky130_fd_sc_hd__mux2_1
XFILLER_0_118_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_113_clk_A clknet_4_6__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_2308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10078_ net1330 net140 net617 vssd1 vssd1 vccd1 vccd1 _00280_ sky130_fd_sc_hd__mux2_1
XANTENNA__10240__S net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_199_482 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_202_453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_128_clk_A clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08098__C1 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_175_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13768_ clknet_leaf_100_clk _01339_ vssd1 vssd1 vccd1 vccd1 top.lcd.cnt_500hz\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_84_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12719_ clknet_leaf_22_clk _00311_ net1024 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[6\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_0_clk clk vssd1 vssd1 vccd1 vccd1 clknet_0_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_155_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13699_ clknet_leaf_71_clk _01270_ vssd1 vssd1 vccd1 vccd1 net115 sky130_fd_sc_hd__dfxtp_1
X_06240_ net1282 net854 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedData\[1\] sky130_fd_sc_hd__and2_1
XANTENNA__07121__Y _02260_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_170_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12464__Q top.ramstore\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06171_ top.a1.halfData\[3\] _01411_ vssd1 vssd1 vccd1 vccd1 _01413_ sky130_fd_sc_hd__nand2_1
XFILLER_0_25_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07073__B1 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold304 top.DUT.register\[20\]\[13\] vssd1 vssd1 vccd1 vccd1 net1420 sky130_fd_sc_hd__dlygate4sd3_1
Xhold315 top.DUT.register\[1\]\[15\] vssd1 vssd1 vccd1 vccd1 net1431 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08233__X _03370_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold326 top.DUT.register\[10\]\[0\] vssd1 vssd1 vccd1 vccd1 net1442 sky130_fd_sc_hd__dlygate4sd3_1
Xhold337 top.DUT.register\[28\]\[13\] vssd1 vssd1 vccd1 vccd1 net1453 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold348 top.a1.hexop\[1\] vssd1 vssd1 vccd1 vccd1 net1464 sky130_fd_sc_hd__dlygate4sd3_1
X_09930_ top.a1.instruction\[30\] net487 net402 top.a1.dataIn\[30\] net398 vssd1 vssd1
+ vccd1 vccd1 _04936_ sky130_fd_sc_hd__a221o_2
XFILLER_0_68_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold359 top.DUT.register\[31\]\[13\] vssd1 vssd1 vccd1 vccd1 net1475 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10415__S net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_15_Right_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout806 _01576_ vssd1 vssd1 vccd1 vccd1 net806 sky130_fd_sc_hd__buf_2
XANTENNA__08962__A2_N net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout817 _05044_ vssd1 vssd1 vccd1 vccd1 net817 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_68_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09861_ net827 _04535_ vssd1 vssd1 vccd1 vccd1 _04873_ sky130_fd_sc_hd__nor2_1
Xfanout828 net829 vssd1 vssd1 vccd1 vccd1 net828 sky130_fd_sc_hd__clkbuf_4
Xfanout839 net840 vssd1 vssd1 vccd1 vccd1 net839 sky130_fd_sc_hd__clkbuf_2
X_08812_ net435 _03920_ _03925_ vssd1 vssd1 vccd1 vccd1 _03926_ sky130_fd_sc_hd__a21bo_1
XPHY_EDGE_ROW_0_Left_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_181_3158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1004 top.DUT.register\[24\]\[29\] vssd1 vssd1 vccd1 vccd1 net2120 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_37_Left_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09792_ _04438_ net486 net401 top.a1.dataIn\[17\] net397 vssd1 vssd1 vccd1 vccd1
+ _04811_ sky130_fd_sc_hd__a221o_1
Xhold1015 top.ramload\[12\] vssd1 vssd1 vccd1 vccd1 net2131 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1026 top.DUT.register\[12\]\[3\] vssd1 vssd1 vccd1 vccd1 net2142 sky130_fd_sc_hd__dlygate4sd3_1
X_08743_ net285 _03859_ vssd1 vssd1 vccd1 vccd1 _03860_ sky130_fd_sc_hd__nand2_1
Xhold1037 top.DUT.register\[8\]\[29\] vssd1 vssd1 vccd1 vccd1 net2153 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12873__CLK clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1048 top.DUT.register\[10\]\[23\] vssd1 vssd1 vccd1 vccd1 net2164 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout181_A _04858_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1059 top.DUT.register\[10\]\[24\] vssd1 vssd1 vccd1 vccd1 net2175 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_197_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13816__1101 vssd1 vssd1 vccd1 vccd1 _13816__1101/HI net1101 sky130_fd_sc_hd__conb_1
XFILLER_0_23_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10150__S net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08674_ net313 _03715_ vssd1 vssd1 vccd1 vccd1 _03794_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_163_2891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07679__A2 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_200_3442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07625_ top.DUT.register\[15\]\[5\] net679 net675 top.DUT.register\[31\]\[5\] vssd1
+ vssd1 vccd1 vccd1 _02764_ sky130_fd_sc_hd__a22o_1
XFILLER_0_191_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_200_3453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_24_Right_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout446_A _01564_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07556_ top.DUT.register\[4\]\[7\] net667 _02687_ _02694_ vssd1 vssd1 vccd1 vccd1
+ _02695_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_196_3390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09825__B1 net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06507_ _01633_ _01634_ _01644_ _01645_ vssd1 vssd1 vccd1 vccd1 _01646_ sky130_fd_sc_hd__or4_1
XFILLER_0_48_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_46_Left_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07487_ top.DUT.register\[23\]\[14\] net573 net556 top.DUT.register\[28\]\[14\] vssd1
+ vssd1 vccd1 vccd1 _02626_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout613_A _04955_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09226_ net132 _04291_ _04293_ _04294_ net897 vssd1 vssd1 vccd1 vccd1 _04295_ sky130_fd_sc_hd__o221a_1
X_06438_ top.a1.instruction\[3\] _01503_ vssd1 vssd1 vccd1 vccd1 _01577_ sky130_fd_sc_hd__nand2_2
XFILLER_0_134_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07851__A2 net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12188__A1 top.a1.row2\[43\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12374__Q top.a1.dataIn\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09157_ _02808_ _02849_ vssd1 vssd1 vccd1 vccd1 _04230_ sky130_fd_sc_hd__xnor2_1
X_06369_ _01474_ _01507_ vssd1 vssd1 vccd1 vccd1 _01508_ sky130_fd_sc_hd__or2_1
XFILLER_0_17_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_380 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08108_ _03243_ _03246_ net291 vssd1 vssd1 vccd1 vccd1 _03247_ sky130_fd_sc_hd__mux2_1
XANTENNA__07064__B1 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09088_ _01546_ _04161_ _04162_ vssd1 vssd1 vccd1 vccd1 _04163_ sky130_fd_sc_hd__and3_1
XANTENNA__07603__A2 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_169_Right_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_33_Right_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_92_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08039_ net332 _02994_ vssd1 vssd1 vccd1 vccd1 _03178_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_92_1831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10325__S net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold860 top.DUT.register\[21\]\[13\] vssd1 vssd1 vccd1 vccd1 net1976 sky130_fd_sc_hd__dlygate4sd3_1
Xhold871 top.DUT.register\[11\]\[15\] vssd1 vssd1 vccd1 vccd1 net1987 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap590 _05003_ vssd1 vssd1 vccd1 vccd1 net590 sky130_fd_sc_hd__buf_1
Xhold882 top.DUT.register\[8\]\[15\] vssd1 vssd1 vccd1 vccd1 net1998 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07982__X _03121_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11050_ net84 net870 net834 net1176 vssd1 vssd1 vccd1 vccd1 _01161_ sky130_fd_sc_hd__a22o_1
Xhold893 top.DUT.register\[28\]\[24\] vssd1 vssd1 vccd1 vccd1 net2009 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout770_X net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_55_Left_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10001_ net192 net1789 net625 vssd1 vssd1 vccd1 vccd1 _00206_ sky130_fd_sc_hd__mux2_1
XANTENNA__09415__A _01983_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06590__A2 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06758__B _01896_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10123__A0 net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_2038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10060__S net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11952_ _05832_ _05834_ vssd1 vssd1 vccd1 vccd1 _05835_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_42_Right_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06878__B1 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10903_ net1600 net188 net479 vssd1 vssd1 vccd1 vccd1 _01064_ sky130_fd_sc_hd__mux2_1
X_11883_ _05762_ _05765_ vssd1 vssd1 vccd1 vccd1 _05766_ sky130_fd_sc_hd__xnor2_1
X_13622_ clknet_leaf_89_clk _01209_ net1003 vssd1 vssd1 vccd1 vccd1 net48 sky130_fd_sc_hd__dfrtp_1
X_10834_ top.DUT.register\[28\]\[10\] net227 net474 vssd1 vssd1 vccd1 vccd1 _00995_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__08619__B2 net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_64_Left_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13553_ clknet_leaf_104_clk _01140_ net974 vssd1 vssd1 vccd1 vccd1 top.ramload\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_10765_ net1396 net253 net482 vssd1 vssd1 vccd1 vccd1 _00926_ sky130_fd_sc_hd__mux2_1
XANTENNA__08037__Y _03176_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_1960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12504_ clknet_leaf_81_clk _00096_ net993 vssd1 vssd1 vccd1 vccd1 top.pc\[16\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_109_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13484_ clknet_leaf_47_clk _01076_ net1091 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[30\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07842__A2 net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10696_ net2004 net145 net334 vssd1 vssd1 vccd1 vccd1 _00857_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_164_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12435_ clknet_leaf_75_clk _00031_ net1079 vssd1 vssd1 vccd1 vccd1 top.ramaddr\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_120_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_51_Right_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07055__B1 net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12366_ clknet_leaf_102_clk top.ru.next_FetchedData\[10\] net980 vssd1 vssd1 vccd1
+ vccd1 top.a1.dataIn\[10\] sky130_fd_sc_hd__dfrtp_4
XPHY_EDGE_ROW_136_Right_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06802__B1 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11317_ _05131_ _05148_ _05194_ vssd1 vssd1 vccd1 vccd1 _05202_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_200_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10235__S net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12297_ _06108_ _06109_ vssd1 vssd1 vccd1 vccd1 _01350_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_73_Left_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10462__C net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_2389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11248_ top.a1.row2\[8\] _05139_ _05140_ top.a1.row2\[32\] vssd1 vssd1 vccd1 vccd1
+ _05141_ sky130_fd_sc_hd__a22o_1
XANTENNA__08555__B1 net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11179_ _05015_ _05027_ net473 net587 net1239 vssd1 vssd1 vccd1 vccd1 _01237_ sky130_fd_sc_hd__a32o_1
XANTENNA__09325__A _02623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_60_Right_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_166_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11293__C _05182_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09612__X _04657_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06869__B1 net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09979__B _04712_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_82_Left_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_46_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07410_ top.DUT.register\[26\]\[9\] net750 net714 top.DUT.register\[27\]\[9\] vssd1
+ vssd1 vccd1 vccd1 _02549_ sky130_fd_sc_hd__a22o_1
XFILLER_0_161_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08390_ _03519_ _03521_ vssd1 vssd1 vccd1 vccd1 _03522_ sky130_fd_sc_hd__xor2_1
XFILLER_0_175_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_147_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10417__A1 _04841_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07341_ top.DUT.register\[28\]\[8\] net558 net448 top.DUT.register\[21\]\[8\] _02479_
+ vssd1 vssd1 vccd1 vccd1 _02480_ sky130_fd_sc_hd__a221o_1
XFILLER_0_174_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_174_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11090__A1 net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07272_ top.DUT.register\[20\]\[13\] net665 net775 top.DUT.register\[13\]\[13\] vssd1
+ vssd1 vccd1 vccd1 _02411_ sky130_fd_sc_hd__a22o_1
XANTENNA__07833__A2 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09011_ _03463_ _03490_ _04085_ vssd1 vssd1 vccd1 vccd1 _04086_ sky130_fd_sc_hd__and3_1
X_06223_ net1278 net856 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedInstr\[17\] sky130_fd_sc_hd__and2_1
XFILLER_0_72_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06690__Y _01829_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06154_ top.a1.dataIn\[14\] vssd1 vssd1 vccd1 vccd1 _01397_ sky130_fd_sc_hd__inv_2
XANTENNA__07046__B1 net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold101 net101 vssd1 vssd1 vccd1 vccd1 net1217 sky130_fd_sc_hd__dlygate4sd3_1
Xhold112 _01323_ vssd1 vssd1 vccd1 vccd1 net1228 sky130_fd_sc_hd__dlygate4sd3_1
Xhold123 top.a1.row1\[107\] vssd1 vssd1 vccd1 vccd1 net1239 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold134 top.a1.row1\[121\] vssd1 vssd1 vccd1 vccd1 net1250 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_103_Right_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold145 top.a1.row1\[9\] vssd1 vssd1 vccd1 vccd1 net1261 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold156 top.a1.row1\[17\] vssd1 vssd1 vccd1 vccd1 net1272 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08898__X _04008_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold167 top.a1.row2\[12\] vssd1 vssd1 vccd1 vccd1 net1283 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09913_ _04918_ _04919_ vssd1 vssd1 vccd1 vccd1 _04920_ sky130_fd_sc_hd__or2_1
Xhold178 top.ramaddr\[19\] vssd1 vssd1 vccd1 vccd1 net1294 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout603 _04957_ vssd1 vssd1 vccd1 vccd1 net603 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_74_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold189 top.ramaddr\[28\] vssd1 vssd1 vccd1 vccd1 net1305 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout614 _04955_ vssd1 vssd1 vccd1 vccd1 net614 sky130_fd_sc_hd__clkbuf_4
Xfanout625 net626 vssd1 vssd1 vccd1 vccd1 net625 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_165_2920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout636 _01629_ vssd1 vssd1 vccd1 vccd1 net636 sky130_fd_sc_hd__clkbuf_4
Xfanout647 _01612_ vssd1 vssd1 vccd1 vccd1 net647 sky130_fd_sc_hd__clkbuf_8
X_09844_ _03869_ net404 net490 _04857_ vssd1 vssd1 vccd1 vccd1 _04858_ sky130_fd_sc_hd__o211a_4
Xfanout658 _01609_ vssd1 vssd1 vccd1 vccd1 net658 sky130_fd_sc_hd__buf_4
Xfanout669 _01599_ vssd1 vssd1 vccd1 vccd1 net669 sky130_fd_sc_hd__buf_6
X_09775_ _03724_ net406 net488 _04795_ vssd1 vssd1 vccd1 vccd1 _04796_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout563_A _01528_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06987_ top.DUT.register\[24\]\[23\] net644 net737 top.DUT.register\[16\]\[23\] vssd1
+ vssd1 vccd1 vccd1 _02126_ sky130_fd_sc_hd__a22o_1
XANTENNA__12380__RESET_B net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08726_ net434 _03840_ _03843_ vssd1 vssd1 vccd1 vccd1 _03844_ sky130_fd_sc_hd__o21ai_1
XANTENNA__12619__CLK clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12369__Q top.a1.dataIn\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_205_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08657_ net321 _03389_ vssd1 vssd1 vccd1 vccd1 _03778_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout730_A _01627_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09889__B _04590_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout351_X net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1093_X net1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout828_A net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout449_X net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07608_ _02742_ _02744_ _02746_ vssd1 vssd1 vccd1 vccd1 _02747_ sky130_fd_sc_hd__or3_1
XFILLER_0_139_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_194_3349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08588_ _02611_ net431 net499 _02613_ vssd1 vssd1 vccd1 vccd1 _03712_ sky130_fd_sc_hd__a22o_1
XFILLER_0_48_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_165_124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_193_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07539_ _02668_ _02677_ vssd1 vssd1 vccd1 vccd1 _02678_ sky130_fd_sc_hd__or2_4
XFILLER_0_48_174 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout616_X net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12769__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10550_ net1974 net200 net355 vssd1 vssd1 vccd1 vccd1 _00717_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_4_10__f_clk_X clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07285__B1 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07824__A2 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09209_ _04261_ _04266_ _04278_ vssd1 vssd1 vccd1 vccd1 _04279_ sky130_fd_sc_hd__and3_1
X_10481_ net1393 net204 net364 vssd1 vssd1 vccd1 vccd1 _00651_ sky130_fd_sc_hd__mux2_1
X_12220_ top.lcd.cnt_20ms\[3\] _06051_ vssd1 vssd1 vccd1 vccd1 _06063_ sky130_fd_sc_hd__xor2_1
X_12151_ _06029_ _06030_ _06032_ vssd1 vssd1 vccd1 vccd1 _06034_ sky130_fd_sc_hd__a21o_1
XANTENNA__10055__S net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09129__B net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08033__B _02994_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11102_ net905 net1895 net860 _05056_ vssd1 vssd1 vccd1 vccd1 _01202_ sky130_fd_sc_hd__a31o_1
XFILLER_0_208_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12082_ _05946_ _05949_ _05963_ vssd1 vssd1 vccd1 vccd1 _05965_ sky130_fd_sc_hd__a21o_1
Xhold690 top.DUT.register\[10\]\[22\] vssd1 vssd1 vccd1 vccd1 net1806 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08537__B1 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11033_ net12 net841 net818 net2181 vssd1 vssd1 vccd1 vccd1 _01145_ sky130_fd_sc_hd__a22o_1
XANTENNA__06488__B _01607_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12984_ clknet_leaf_125_clk _00576_ net924 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[15\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_188_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11844__B1 top.a1.dataIn\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11935_ _05758_ _05786_ vssd1 vssd1 vccd1 vccd1 _05818_ sky130_fd_sc_hd__nand2_2
XANTENNA__09799__B _04453_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_197_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11866_ _05715_ _05741_ _05713_ vssd1 vssd1 vccd1 vccd1 _05749_ sky130_fd_sc_hd__a21o_1
XFILLER_0_28_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08048__X _03187_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_184_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13605_ clknet_leaf_89_clk _01192_ net1002 vssd1 vssd1 vccd1 vccd1 net40 sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_205_Right_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10817_ net170 net1494 net599 vssd1 vssd1 vccd1 vccd1 _00978_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_31_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_483 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11797_ _05655_ _05656_ _05643_ _05651_ vssd1 vssd1 vccd1 vccd1 _05680_ sky130_fd_sc_hd__a211o_1
XFILLER_0_131_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_2229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13536_ clknet_leaf_93_clk _01123_ net995 vssd1 vssd1 vccd1 vccd1 top.a1.data\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07276__B1 net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10748_ net1885 net202 net420 vssd1 vssd1 vccd1 vccd1 _00909_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07815__A2 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06791__X _01930_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13467_ clknet_leaf_125_clk _01059_ net923 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[30\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_10679_ net1473 net218 net338 vssd1 vssd1 vccd1 vccd1 _00842_ sky130_fd_sc_hd__mux2_1
XFILLER_0_180_683 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13815__1100 vssd1 vssd1 vccd1 vccd1 _13815__1100/HI net1100 sky130_fd_sc_hd__conb_1
X_12418_ clknet_leaf_110_clk top.ru.next_FetchedInstr\[30\] net977 vssd1 vssd1 vccd1
+ vccd1 top.a1.instruction\[30\] sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_132_2429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13398_ clknet_leaf_4_clk _00990_ net940 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[28\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_140_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12349_ net2204 net118 _00016_ vssd1 vssd1 vccd1 vccd1 _01374_ sky130_fd_sc_hd__mux2_1
XANTENNA__08528__B1 _03643_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08878__B _03987_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06910_ _02047_ _02048_ vssd1 vssd1 vccd1 vccd1 _02049_ sky130_fd_sc_hd__or2_4
XTAP_TAPCELL_ROW_56_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07890_ top.DUT.register\[24\]\[1\] net513 net453 top.DUT.register\[29\]\[1\] _03028_
+ vssd1 vssd1 vccd1 vccd1 _03029_ sky130_fd_sc_hd__a221o_1
XANTENNA__09055__A _03980_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_147_2650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06841_ top.DUT.register\[13\]\[19\] net464 net525 top.DUT.register\[11\]\[19\] vssd1
+ vssd1 vccd1 vccd1 _01980_ sky130_fd_sc_hd__a22o_1
XANTENNA__09740__A2 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06554__A2 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11820__A1_N top.a1.dataIn\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09560_ _04591_ _04593_ _04608_ vssd1 vssd1 vccd1 vccd1 _04609_ sky130_fd_sc_hd__o21ai_1
XPHY_EDGE_ROW_90_Left_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06772_ top.DUT.register\[25\]\[24\] net780 net760 top.DUT.register\[30\]\[24\] vssd1
+ vssd1 vccd1 vccd1 _01911_ sky130_fd_sc_hd__a22o_1
XFILLER_0_78_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_160_2850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08511_ net886 top.pc\[11\] net697 _03638_ vssd1 vssd1 vccd1 vccd1 _03639_ sky130_fd_sc_hd__a22o_1
XFILLER_0_210_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_wire417_X net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09491_ _01887_ _01896_ _04543_ vssd1 vssd1 vccd1 vccd1 _04544_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_77_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08700__B1 net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08442_ _02571_ _03571_ vssd1 vssd1 vccd1 vccd1 _03572_ sky130_fd_sc_hd__or2_1
XFILLER_0_148_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_176_3079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08373_ _03169_ _03505_ vssd1 vssd1 vccd1 vccd1 _03506_ sky130_fd_sc_hd__nor2_1
XFILLER_0_92_228 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout144_A net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07324_ _02457_ _02459_ _02461_ _02462_ vssd1 vssd1 vccd1 vccd1 _02463_ sky130_fd_sc_hd__or4_1
XANTENNA__07267__B1 net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07255_ top.DUT.register\[30\]\[13\] net581 net506 top.DUT.register\[27\]\[13\] _02393_
+ vssd1 vssd1 vccd1 vccd1 _02394_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout311_A net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08988__A_N _03256_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_363 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07019__B1 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06206_ top.ramload\[0\] net857 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedInstr\[0\]
+ sky130_fd_sc_hd__and2_1
X_07186_ top.DUT.register\[30\]\[10\] net579 net451 top.DUT.register\[29\]\[10\] _02324_
+ vssd1 vssd1 vccd1 vccd1 _02325_ sky130_fd_sc_hd__a221o_1
XFILLER_0_41_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_170_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_197_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout400 _04975_ vssd1 vssd1 vccd1 vccd1 net400 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout680_A _01547_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout411 _02358_ vssd1 vssd1 vccd1 vccd1 net411 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08519__B1 net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout778_A net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout422 _04470_ vssd1 vssd1 vccd1 vccd1 net422 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06793__A2 net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10603__S net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout433 _03184_ vssd1 vssd1 vccd1 vccd1 net433 sky130_fd_sc_hd__clkbuf_4
Xfanout444 _01564_ vssd1 vssd1 vccd1 vccd1 net444 sky130_fd_sc_hd__clkbuf_4
Xfanout455 _01553_ vssd1 vssd1 vccd1 vccd1 net455 sky130_fd_sc_hd__clkbuf_8
Xfanout466 _01529_ vssd1 vssd1 vccd1 vccd1 net466 sky130_fd_sc_hd__buf_4
Xfanout477 _04969_ vssd1 vssd1 vccd1 vccd1 net477 sky130_fd_sc_hd__clkbuf_8
X_09827_ _04833_ _04836_ _04834_ vssd1 vssd1 vccd1 vccd1 _04842_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_129_Left_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout488 net491 vssd1 vssd1 vccd1 vccd1 net488 sky130_fd_sc_hd__buf_4
XANTENNA__06545__A2 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout945_A net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout566_X net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout499 net502 vssd1 vssd1 vccd1 vccd1 net499 sky130_fd_sc_hd__clkbuf_4
X_09758_ net1689 net209 net633 vssd1 vssd1 vccd1 vccd1 _00134_ sky130_fd_sc_hd__mux2_1
X_08709_ net497 _03812_ _03816_ _03342_ _03827_ vssd1 vssd1 vccd1 vccd1 _03828_ sky130_fd_sc_hd__o221a_1
XFILLER_0_69_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_87_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_512 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout733_X net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09689_ net1980 net144 net631 vssd1 vssd1 vccd1 vccd1 _00121_ sky130_fd_sc_hd__mux2_1
XFILLER_0_139_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11720_ _05596_ _05600_ _05602_ _05592_ vssd1 vssd1 vccd1 vccd1 _05603_ sky130_fd_sc_hd__o31ai_2
XFILLER_0_194_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_179_794 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09412__B _01585_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11651_ _05509_ _05531_ vssd1 vssd1 vccd1 vccd1 _05534_ sky130_fd_sc_hd__xor2_2
XANTENNA_fanout900_X net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_181_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10602_ net243 net2020 net346 vssd1 vssd1 vccd1 vccd1 _00767_ sky130_fd_sc_hd__mux2_1
XANTENNA__07258__B1 net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_138_Left_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11582_ _05426_ _05454_ vssd1 vssd1 vccd1 vccd1 _05465_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_64_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_181_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13321_ clknet_leaf_52_clk _00913_ net1037 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[25\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_10533_ net1571 net259 net356 vssd1 vssd1 vccd1 vccd1 _00700_ sky130_fd_sc_hd__mux2_1
XANTENNA__08470__A2 _03534_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_9__f_clk_X clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13252_ clknet_leaf_37_clk _00844_ net1052 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[23\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_10464_ net1544 net267 net363 vssd1 vssd1 vccd1 vccd1 _00634_ sky130_fd_sc_hd__mux2_1
XFILLER_0_161_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12203_ net1171 net688 vssd1 vssd1 vccd1 vccd1 _06050_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_114_2159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12649__RESET_B net1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13183_ clknet_leaf_24_clk _00775_ net1013 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[21\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_10395_ _04153_ _04949_ net400 vssd1 vssd1 vccd1 vccd1 _04983_ sky130_fd_sc_hd__and3_1
X_12134_ _06001_ _06003_ _06008_ _06015_ vssd1 vssd1 vccd1 vccd1 _06017_ sky130_fd_sc_hd__a22o_1
XFILLER_0_130_591 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06784__A2 net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_208_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12065_ _05932_ _05942_ _05946_ _05947_ vssd1 vssd1 vccd1 vccd1 _05948_ sky130_fd_sc_hd__a31oi_4
XANTENNA__10513__S net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11016_ net24 net841 net818 top.ramload\[2\] vssd1 vssd1 vccd1 vccd1 _01128_ sky130_fd_sc_hd__a22o_1
XFILLER_0_189_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06536__A2 net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_129_2380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12967_ clknet_leaf_6_clk _00559_ net944 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[14\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_142_2580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11918_ _05799_ _05800_ vssd1 vssd1 vccd1 vccd1 _05801_ sky130_fd_sc_hd__or2_1
XANTENNA__07497__B1 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12898_ clknet_leaf_10_clk _00490_ net950 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[12\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_75_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_185_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11849_ top.a1.dataIn\[6\] _05664_ _05699_ vssd1 vssd1 vccd1 vccd1 _05732_ sky130_fd_sc_hd__or3_1
XFILLER_0_27_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_818 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13519_ clknet_leaf_22_clk _01111_ net1035 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[31\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_363 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload10 clknet_leaf_127_clk vssd1 vssd1 vccd1 vccd1 clkload10/Y sky130_fd_sc_hd__clkinv_4
X_07040_ _02177_ _02178_ vssd1 vssd1 vccd1 vccd1 _02179_ sky130_fd_sc_hd__nand2b_2
Xclkload21 clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 clkload21/Y sky130_fd_sc_hd__clkinv_2
Xclkload32 clknet_leaf_104_clk vssd1 vssd1 vccd1 vccd1 clkload32/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_30_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13568__Q top.ramload\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload43 clknet_leaf_100_clk vssd1 vssd1 vccd1 vccd1 clkload43/Y sky130_fd_sc_hd__clkinv_4
XTAP_TAPCELL_ROW_58_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08749__B1 net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload54 clknet_leaf_90_clk vssd1 vssd1 vccd1 vccd1 clkload54/X sky130_fd_sc_hd__clkbuf_8
Xclkload65 clknet_leaf_15_clk vssd1 vssd1 vccd1 vccd1 clkload65/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload76 clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 clkload76/Y sky130_fd_sc_hd__clkinv_4
Xclkload87 clknet_leaf_54_clk vssd1 vssd1 vccd1 vccd1 clkload87/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_2_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload98 clknet_leaf_76_clk vssd1 vssd1 vccd1 vccd1 clkload98/Y sky130_fd_sc_hd__clkinv_16
XFILLER_0_167_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08991_ _03653_ _03678_ vssd1 vssd1 vccd1 vccd1 _04066_ sky130_fd_sc_hd__nand2_1
XANTENNA__06775__A2 net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07942_ _02050_ _02242_ _02262_ _03079_ vssd1 vssd1 vccd1 vccd1 _03081_ sky130_fd_sc_hd__o31ai_1
XANTENNA__10423__S net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08401__B net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09713__A2 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07873_ top.DUT.register\[29\]\[1\] net724 net700 top.DUT.register\[31\]\[1\] _03008_
+ vssd1 vssd1 vccd1 vccd1 _03012_ sky130_fd_sc_hd__a221o_1
XFILLER_0_207_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06527__A2 net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09612_ top.a1.halfData\[3\] net888 _01411_ top.a1.halfData\[5\] vssd1 vssd1 vccd1
+ vccd1 _04657_ sky130_fd_sc_hd__and4b_2
X_06824_ _01940_ _01961_ vssd1 vssd1 vccd1 vccd1 _01963_ sky130_fd_sc_hd__nor2_1
XFILLER_0_183_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_178_3119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09543_ _04578_ _04582_ _04592_ vssd1 vssd1 vccd1 vccd1 _04593_ sky130_fd_sc_hd__a21oi_1
X_06755_ top.DUT.register\[17\]\[24\] net461 net445 top.DUT.register\[1\]\[24\] vssd1
+ vssd1 vccd1 vccd1 _01894_ sky130_fd_sc_hd__a22o_1
XFILLER_0_78_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout261_A net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout359_A net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07488__B1 net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09232__B _02502_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09474_ _02199_ _04514_ _04517_ vssd1 vssd1 vccd1 vccd1 _04528_ sky130_fd_sc_hd__a21o_1
X_06686_ top.DUT.register\[5\]\[26\] net654 net768 top.DUT.register\[28\]\[26\] _01824_
+ vssd1 vssd1 vccd1 vccd1 _01825_ sky130_fd_sc_hd__a221o_1
XFILLER_0_176_742 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08425_ net319 _03555_ vssd1 vssd1 vccd1 vccd1 _03556_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_191_3308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout147_X net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout526_A _01554_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11036__B2 top.ramload\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08356_ net1462 net832 net802 _03489_ vssd1 vssd1 vccd1 vccd1 _00023_ sky130_fd_sc_hd__a22o_1
XFILLER_0_191_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08416__X _03548_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload4 clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 clkload4/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_46_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07307_ top.DUT.register\[16\]\[12\] net543 net443 top.DUT.register\[1\]\[12\] vssd1
+ vssd1 vccd1 vccd1 _02446_ sky130_fd_sc_hd__a22o_1
XFILLER_0_73_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_22_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_199 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08287_ _03413_ _03422_ vssd1 vssd1 vccd1 vccd1 _03423_ sky130_fd_sc_hd__xnor2_1
XANTENNA__08452__A2 net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout314_X net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_210_3603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07238_ top.DUT.register\[10\]\[10\] net770 net710 top.DUT.register\[11\]\[10\] vssd1
+ vssd1 vccd1 vccd1 _02377_ sky130_fd_sc_hd__a22o_1
XFILLER_0_33_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09401__A1 net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07169_ _02307_ vssd1 vssd1 vccd1 vccd1 _02308_ sky130_fd_sc_hd__inv_2
XANTENNA__08799__A _01877_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07412__B1 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10180_ top.a1.instruction\[11\] _04153_ _04949_ vssd1 vssd1 vccd1 vccd1 _04960_
+ sky130_fd_sc_hd__and3_1
XANTENNA__06766__A2 net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07963__A1 _01572_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09407__B _04453_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10333__S net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout230 _04763_ vssd1 vssd1 vccd1 vccd1 net230 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout241 net242 vssd1 vssd1 vccd1 vccd1 net241 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_208_3565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout252 _04741_ vssd1 vssd1 vccd1 vccd1 net252 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout263 net264 vssd1 vssd1 vccd1 vccd1 net263 sky130_fd_sc_hd__clkbuf_2
Xfanout274 _03238_ vssd1 vssd1 vccd1 vccd1 net274 sky130_fd_sc_hd__clkbuf_4
Xfanout285 _03170_ vssd1 vssd1 vccd1 vccd1 net285 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07715__A1 top.a1.instruction\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout296 net297 vssd1 vssd1 vccd1 vccd1 net296 sky130_fd_sc_hd__buf_4
XANTENNA__07715__B2 top.a1.instruction\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07191__A2 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12821_ clknet_leaf_29_clk _00413_ net1019 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[10\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_202_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_2_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11275__A1 top.a1.row2\[34\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07479__B1 net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09142__B _02899_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12752_ clknet_leaf_29_clk _00344_ net1017 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[7\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08039__A net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11703_ top.a1.dataIn\[9\] _05583_ _05584_ vssd1 vssd1 vccd1 vccd1 _05586_ sky130_fd_sc_hd__or3_1
XFILLER_0_84_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09710__X _04741_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_194_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12683_ clknet_leaf_45_clk _00275_ net1065 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[5\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_182_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11634_ _05516_ vssd1 vssd1 vccd1 vccd1 _05517_ sky130_fd_sc_hd__inv_2
XANTENNA__12224__B1 net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_181_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11565_ _01397_ net250 _05418_ vssd1 vssd1 vccd1 vccd1 _05448_ sky130_fd_sc_hd__a21boi_1
XANTENNA__10508__S net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08045__Y _03184_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13304_ clknet_leaf_128_clk _00896_ net911 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[25\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_10516_ net2129 net201 net359 vssd1 vssd1 vccd1 vccd1 _00685_ sky130_fd_sc_hd__mux2_1
XANTENNA__07651__B1 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11496_ _05376_ _05378_ _05346_ vssd1 vssd1 vccd1 vccd1 _05379_ sky130_fd_sc_hd__nor3b_1
XFILLER_0_12_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13235_ clknet_leaf_124_clk _00827_ net926 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[23\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_10447_ net217 net1724 net367 vssd1 vssd1 vccd1 vccd1 _00618_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_686 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07403__B1 net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13166_ clknet_leaf_43_clk _00758_ net1062 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[20\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_10378_ net1599 net226 net374 vssd1 vssd1 vccd1 vccd1 _00553_ sky130_fd_sc_hd__mux2_1
X_12117_ _05980_ _05992_ vssd1 vssd1 vccd1 vccd1 _06000_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10243__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13097_ clknet_leaf_52_clk _00689_ net1038 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[18\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_12048_ _05912_ _05919_ vssd1 vssd1 vccd1 vccd1 _05931_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_205_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06509__A2 net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07182__A2 net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13112__CLK clknet_leaf_128_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_177_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_140_2539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_204_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06540_ _01678_ vssd1 vssd1 vccd1 vccd1 _01679_ sky130_fd_sc_hd__inv_2
XANTENNA__09052__B _03673_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06471_ net787 _01594_ _01602_ vssd1 vssd1 vccd1 vccd1 _01610_ sky130_fd_sc_hd__and3_4
XFILLER_0_173_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08210_ _03347_ vssd1 vssd1 vccd1 vccd1 _03348_ sky130_fd_sc_hd__inv_2
XFILLER_0_173_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_173_3038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11018__A1 net28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09190_ _02723_ _02728_ vssd1 vssd1 vccd1 vccd1 _04261_ sky130_fd_sc_hd__or2_1
XANTENNA__07890__B1 net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06692__A _01809_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_464 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08141_ _03277_ _03278_ vssd1 vssd1 vccd1 vccd1 _03279_ sky130_fd_sc_hd__nand2_1
XFILLER_0_43_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10418__S net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09631__A1 _04164_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_155_2771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkload110 clknet_leaf_66_clk vssd1 vssd1 vccd1 vccd1 clkload110/Y sky130_fd_sc_hd__inv_12
X_08072_ _03209_ _03210_ vssd1 vssd1 vccd1 vccd1 _03211_ sky130_fd_sc_hd__nand2_1
XFILLER_0_43_467 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07642__B1 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07023_ top.DUT.register\[12\]\[20\] net740 net638 top.DUT.register\[6\]\[20\] _02161_
+ vssd1 vssd1 vccd1 vccd1 _02162_ sky130_fd_sc_hd__a221o_1
XFILLER_0_140_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_188_3270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09395__B1 _04453_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10153__S net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08974_ _01655_ net692 net1136 net875 vssd1 vssd1 vccd1 vccd1 _00080_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA_fanout1016_A net1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold16 top.a1.dataInTemp\[7\] vssd1 vssd1 vccd1 vccd1 net1132 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_89_Right_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09942__S net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold27 top.ramstore\[14\] vssd1 vssd1 vccd1 vccd1 net1143 sky130_fd_sc_hd__dlygate4sd3_1
X_07925_ _02453_ _02473_ vssd1 vssd1 vccd1 vccd1 _03064_ sky130_fd_sc_hd__nor2_1
Xhold38 top.ramstore\[19\] vssd1 vssd1 vccd1 vccd1 net1154 sky130_fd_sc_hd__dlygate4sd3_1
Xhold49 top.a1.data\[2\] vssd1 vssd1 vccd1 vccd1 net1165 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09698__A1 top.a1.dataIn\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout476_A net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07856_ net301 _02994_ vssd1 vssd1 vccd1 vccd1 _02995_ sky130_fd_sc_hd__nor2_1
XANTENNA__06867__A _01983_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07173__A2 net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06807_ top.DUT.register\[5\]\[17\] net652 net648 top.DUT.register\[22\]\[17\] vssd1
+ vssd1 vccd1 vccd1 _01946_ sky130_fd_sc_hd__a22o_1
XFILLER_0_211_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07787_ top.DUT.register\[18\]\[2\] net547 net527 top.DUT.register\[26\]\[2\] vssd1
+ vssd1 vccd1 vccd1 _02926_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_84_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06381__B1 net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout643_A _01613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_203_3484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_203_3495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09526_ top.a1.instruction\[26\] net821 net422 vssd1 vssd1 vccd1 vccd1 _04577_ sky130_fd_sc_hd__a21o_2
XFILLER_0_211_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06738_ _01874_ _01876_ vssd1 vssd1 vccd1 vccd1 _01877_ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_27_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08122__A1 net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09457_ _04510_ _04511_ vssd1 vssd1 vccd1 vccd1 _04512_ sky130_fd_sc_hd__and2b_1
XFILLER_0_210_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06669_ _01801_ _01803_ _01805_ _01807_ vssd1 vssd1 vccd1 vccd1 _01808_ sky130_fd_sc_hd__or4_1
XFILLER_0_164_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout810_A net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout431_X net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_420 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout908_A _01405_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout529_X net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08408_ _02678_ net330 _03294_ vssd1 vssd1 vccd1 vccd1 _03540_ sky130_fd_sc_hd__o21ai_1
XPHY_EDGE_ROW_98_Right_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_639 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07881__A0 _03000_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09388_ _04433_ _04434_ _04431_ vssd1 vssd1 vccd1 vccd1 _04447_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_164_767 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08339_ net322 _03472_ _03466_ vssd1 vssd1 vccd1 vccd1 _03473_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_163_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_434 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11350_ _05214_ _05219_ top.a1.dataIn\[24\] vssd1 vssd1 vccd1 vccd1 _05233_ sky130_fd_sc_hd__a21oi_1
X_10301_ net254 net1933 net381 vssd1 vssd1 vccd1 vccd1 _00478_ sky130_fd_sc_hd__mux2_1
XANTENNA__06987__A2 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08025__C _03157_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11281_ top.a1.row1\[3\] _05124_ _05125_ top.a1.row1\[19\] vssd1 vssd1 vccd1 vccd1
+ _05171_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_111_2107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_95_1873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_2118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13020_ clknet_leaf_130_clk _00612_ net910 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[16\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_10232_ net264 net2154 net389 vssd1 vssd1 vccd1 vccd1 _00411_ sky130_fd_sc_hd__mux2_1
XANTENNA__11193__B1 net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1003 net1004 vssd1 vssd1 vccd1 vccd1 net1003 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10063__S net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10163_ net1260 net217 net604 vssd1 vssd1 vccd1 vccd1 _00362_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08041__B _03172_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1014 net1016 vssd1 vssd1 vccd1 vccd1 net1014 sky130_fd_sc_hd__clkbuf_4
Xfanout1025 net1071 vssd1 vssd1 vccd1 vccd1 net1025 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09705__X _04737_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1036 net1039 vssd1 vssd1 vccd1 vccd1 net1036 sky130_fd_sc_hd__clkbuf_2
XANTENNA__13135__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1047 net1048 vssd1 vssd1 vccd1 vccd1 net1047 sky130_fd_sc_hd__clkbuf_2
XANTENNA_input37_A gpio_in[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10094_ net1368 net196 net611 vssd1 vssd1 vccd1 vccd1 _00295_ sky130_fd_sc_hd__mux2_1
Xfanout1058 net1070 vssd1 vssd1 vccd1 vccd1 net1058 sky130_fd_sc_hd__clkbuf_4
Xfanout1069 net1070 vssd1 vssd1 vccd1 vccd1 net1069 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08976__B _01393_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07164__A2 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12804_ clknet_leaf_36_clk _00396_ net1049 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[9\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_13784_ clknet_leaf_68_clk net1266 vssd1 vssd1 vccd1 vccd1 top.pad.button_control.r_counter\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__08992__A _03736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10996_ top.a1.dataInTemp\[8\] _04999_ vssd1 vssd1 vccd1 vccd1 _05031_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_122_2269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_695 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12735_ clknet_leaf_19_clk _00327_ net1026 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[7\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_123_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_201_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12666_ clknet_leaf_1_clk _00258_ net916 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[5\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11617_ top.a1.dataIn\[13\] _05418_ _05451_ vssd1 vssd1 vccd1 vccd1 _05500_ sky130_fd_sc_hd__or3_1
XANTENNA__10238__S net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12597_ clknet_leaf_29_clk _00189_ net1019 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[3\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_154_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11548_ _05378_ _05406_ _05410_ _05415_ vssd1 vssd1 vccd1 vccd1 _05431_ sky130_fd_sc_hd__or4b_1
XFILLER_0_123_631 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06978__A2 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold508 top.DUT.register\[22\]\[3\] vssd1 vssd1 vccd1 vccd1 net1624 sky130_fd_sc_hd__dlygate4sd3_1
Xhold519 top.DUT.register\[19\]\[21\] vssd1 vssd1 vccd1 vccd1 net1635 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_38_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11479_ _01396_ net273 _05328_ vssd1 vssd1 vccd1 vccd1 _05362_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_12_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13218_ clknet_leaf_25_clk _00810_ net1012 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[22\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_150_2690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11184__B1 net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_196_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13149_ clknet_leaf_13_clk _00741_ net953 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[20\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_148_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_51_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07710_ _02839_ _02848_ vssd1 vssd1 vccd1 vccd1 _02849_ sky130_fd_sc_hd__nor2_8
X_08690_ _01983_ _02004_ _02047_ vssd1 vssd1 vccd1 vccd1 _03809_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10701__S net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07155__A2 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07641_ top.DUT.register\[25\]\[5\] net778 net754 top.DUT.register\[1\]\[5\] vssd1
+ vssd1 vccd1 vccd1 _02780_ sky130_fd_sc_hd__a22o_1
XFILLER_0_178_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06902__A2 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07572_ top.DUT.register\[3\]\[6\] net551 net455 top.DUT.register\[25\]\[6\] vssd1
+ vssd1 vccd1 vccd1 _02711_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_66_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09311_ net132 _04367_ _04374_ net810 net897 vssd1 vssd1 vccd1 vccd1 _04375_ sky130_fd_sc_hd__o221a_1
X_06523_ top.DUT.register\[6\]\[29\] net570 net525 top.DUT.register\[11\]\[29\] vssd1
+ vssd1 vccd1 vccd1 _01662_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_157_2800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08655__A2 _03387_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09242_ net898 top.pc\[9\] _04309_ net889 vssd1 vssd1 vccd1 vccd1 _00089_ sky130_fd_sc_hd__o211a_1
XFILLER_0_7_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06454_ top.a1.instruction\[22\] net792 vssd1 vssd1 vccd1 vccd1 _01593_ sky130_fd_sc_hd__nand2_1
XANTENNA__09510__B _04560_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07863__B1 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09173_ _02808_ _02849_ _04232_ vssd1 vssd1 vccd1 vccd1 _04245_ sky130_fd_sc_hd__o21a_1
X_06385_ _01511_ _01521_ _01523_ vssd1 vssd1 vccd1 vccd1 _01524_ sky130_fd_sc_hd__and3_1
XANTENNA__10148__S net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout224_A _04805_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08124_ _03160_ _03181_ vssd1 vssd1 vccd1 vccd1 _03263_ sky130_fd_sc_hd__nor2_2
XFILLER_0_43_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_415 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_584 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06969__A2 net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08055_ net330 _03122_ _03193_ vssd1 vssd1 vccd1 vccd1 _03194_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_3_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_186_3229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07006_ _02138_ _02140_ _02142_ _02144_ vssd1 vssd1 vccd1 vccd1 _02145_ sky130_fd_sc_hd__or4_1
XANTENNA__08142__A _02544_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout593_A _04971_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07918__A1 _02678_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_168_2962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_168_2973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07394__A2 net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_208_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08957_ _02428_ net692 net1199 net875 vssd1 vssd1 vccd1 vccd1 _00063_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA_fanout381_X net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout760_A _01617_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_205_3524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06868__Y _02007_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout858_A net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout479_X net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10611__S net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07908_ _02947_ _03046_ vssd1 vssd1 vccd1 vccd1 _03047_ sky130_fd_sc_hd__nor2_1
X_08888_ net306 _03917_ _03997_ net282 vssd1 vssd1 vccd1 vccd1 _03998_ sky130_fd_sc_hd__a211o_1
X_07839_ top.DUT.register\[30\]\[0\] net579 net439 top.DUT.register\[5\]\[0\] vssd1
+ vssd1 vccd1 vccd1 _02978_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout646_X net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10850_ net1867 net164 net476 vssd1 vssd1 vccd1 vccd1 _01011_ sky130_fd_sc_hd__mux2_1
XFILLER_0_211_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09509_ _01854_ _04560_ vssd1 vssd1 vccd1 vccd1 _04561_ sky130_fd_sc_hd__nand2_1
X_10781_ net1246 net193 net485 vssd1 vssd1 vccd1 vccd1 _00942_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout813_X net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12520_ clknet_leaf_88_clk _00112_ net1001 vssd1 vssd1 vccd1 vccd1 top.a1.state\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_149_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_164_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_117_Right_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12451_ clknet_leaf_72_clk _00047_ net1080 vssd1 vssd1 vccd1 vccd1 top.ramaddr\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10058__S net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_1902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11402_ _05277_ _05282_ _05284_ vssd1 vssd1 vccd1 vccd1 _05285_ sky130_fd_sc_hd__a21o_2
XANTENNA__07606__B1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12382_ clknet_leaf_110_clk top.ru.next_FetchedData\[26\] net976 vssd1 vssd1 vccd1
+ vccd1 top.a1.dataIn\[26\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_62_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11333_ top.a1.dataIn\[22\] top.a1.dataIn\[21\] top.a1.dataIn\[23\] vssd1 vssd1 vccd1
+ vccd1 _05216_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_105_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09148__A top.pc\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11264_ top.a1.row2\[1\] _05143_ _05153_ _01382_ _05155_ vssd1 vssd1 vccd1 vccd1
+ _05156_ sky130_fd_sc_hd__a221o_1
XFILLER_0_120_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11166__A0 top.a1.row1\[59\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07909__A1 net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13003_ clknet_leaf_45_clk _00595_ net1069 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[15\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_10215_ net204 net1697 net395 vssd1 vssd1 vccd1 vccd1 _00395_ sky130_fd_sc_hd__mux2_1
X_11195_ net1350 net588 vssd1 vssd1 vccd1 vccd1 _01248_ sky130_fd_sc_hd__nand2b_1
XANTENNA__11181__A3 net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_207_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10146_ net1934 net146 net603 vssd1 vssd1 vccd1 vccd1 _00345_ sky130_fd_sc_hd__mux2_1
XFILLER_0_118_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06593__B1 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10521__S net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10077_ net1797 net150 net617 vssd1 vssd1 vccd1 vccd1 _00279_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_124_2309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkload2_A clknet_4_6__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13767_ clknet_leaf_100_clk _01338_ vssd1 vssd1 vccd1 vccd1 top.lcd.cnt_500hz\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_48_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09295__C1 net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10979_ top.a1.data\[0\] net784 vssd1 vssd1 vccd1 vccd1 _05018_ sky130_fd_sc_hd__or2_1
XFILLER_0_57_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12718_ clknet_leaf_39_clk _00310_ net1054 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[6\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_139_2530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12180__A2_N _05083_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13698_ clknet_leaf_73_clk _01269_ vssd1 vssd1 vccd1 vccd1 net114 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_143_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_61_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_182_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12649_ clknet_leaf_53_clk _00241_ net1038 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[4\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_150_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10195__C net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06170_ top.a1.halfData\[3\] _01411_ vssd1 vssd1 vccd1 vccd1 _01412_ sky130_fd_sc_hd__and2_1
XFILLER_0_142_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_152_2730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold305 top.DUT.register\[19\]\[13\] vssd1 vssd1 vccd1 vccd1 net1421 sky130_fd_sc_hd__dlygate4sd3_1
Xhold316 top.DUT.register\[20\]\[12\] vssd1 vssd1 vccd1 vccd1 net1432 sky130_fd_sc_hd__dlygate4sd3_1
Xhold327 top.DUT.register\[9\]\[9\] vssd1 vssd1 vccd1 vccd1 net1443 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold338 top.DUT.register\[25\]\[26\] vssd1 vssd1 vccd1 vccd1 net1454 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_159_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold349 top.DUT.register\[2\]\[15\] vssd1 vssd1 vccd1 vccd1 net1465 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout807 net809 vssd1 vssd1 vccd1 vccd1 net807 sky130_fd_sc_hd__clkbuf_4
X_09860_ _04869_ _04870_ vssd1 vssd1 vccd1 vccd1 _04872_ sky130_fd_sc_hd__xnor2_1
XANTENNA__08022__B1 _03151_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout818 net819 vssd1 vssd1 vccd1 vccd1 net818 sky130_fd_sc_hd__buf_2
Xfanout829 _01504_ vssd1 vssd1 vccd1 vccd1 net829 sky130_fd_sc_hd__buf_4
XANTENNA__07376__A2 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08573__A1 net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08811_ _03260_ _03921_ _03922_ _03348_ _03924_ vssd1 vssd1 vccd1 vccd1 _03925_ sky130_fd_sc_hd__o221a_1
XANTENNA__08573__B2 net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09791_ _04807_ _04808_ _04806_ vssd1 vssd1 vccd1 vccd1 _04810_ sky130_fd_sc_hd__o21ai_1
XANTENNA__06584__B1 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1005 top.DUT.register\[2\]\[19\] vssd1 vssd1 vccd1 vccd1 net2121 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_181_3159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1016 top.pad.button_control.r_counter\[5\] vssd1 vssd1 vccd1 vccd1 net2132 sky130_fd_sc_hd__dlygate4sd3_1
X_08742_ _03774_ _03858_ net308 vssd1 vssd1 vccd1 vccd1 _03859_ sky130_fd_sc_hd__mux2_1
Xhold1027 top.DUT.register\[26\]\[27\] vssd1 vssd1 vccd1 vccd1 net2143 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1038 top.DUT.register\[10\]\[2\] vssd1 vssd1 vccd1 vccd1 net2154 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10431__S net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1049 top.DUT.register\[9\]\[20\] vssd1 vssd1 vccd1 vccd1 net2165 sky130_fd_sc_hd__dlygate4sd3_1
X_08673_ _03333_ _03419_ net320 vssd1 vssd1 vccd1 vccd1 _03793_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_178_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08876__A2 net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_163_2892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout174_A _04876_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_205_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07624_ _02756_ _02758_ _02760_ _02762_ vssd1 vssd1 vccd1 vccd1 _02763_ sky130_fd_sc_hd__or4_2
XFILLER_0_178_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_200_3443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09080__X _04155_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07740__S net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09521__A top.pc\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07555_ top.DUT.register\[5\]\[7\] net651 net635 top.DUT.register\[6\]\[7\] _02690_
+ vssd1 vssd1 vccd1 vccd1 _02694_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout341_A _04993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09825__A1 _03829_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_196_3380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_196_3391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout439_A _01566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12515__RESET_B net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1083_A net1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_192_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06506_ top.DUT.register\[12\]\[30\] net740 net708 top.DUT.register\[15\]\[30\] _01636_
+ vssd1 vssd1 vccd1 vccd1 _01645_ sky130_fd_sc_hd__a221o_1
XANTENNA__07836__A0 _02952_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07486_ top.DUT.register\[29\]\[14\] net453 _02624_ vssd1 vssd1 vccd1 vccd1 _02625_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_48_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07300__A2 net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_180_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09225_ _04276_ _04280_ _04292_ net810 vssd1 vssd1 vccd1 vccd1 _04294_ sky130_fd_sc_hd__a31o_1
XPHY_EDGE_ROW_101_Left_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06437_ _01388_ net826 vssd1 vssd1 vccd1 vccd1 _01576_ sky130_fd_sc_hd__nor2_1
XFILLER_0_16_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12188__A2 net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09156_ _04225_ _04228_ vssd1 vssd1 vccd1 vccd1 _04229_ sky130_fd_sc_hd__xnor2_1
X_06368_ _01484_ net810 vssd1 vssd1 vccd1 vccd1 _01507_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_79_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08107_ _03244_ _03245_ vssd1 vssd1 vccd1 vccd1 _03246_ sky130_fd_sc_hd__and2_1
XFILLER_0_31_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09087_ net895 top.a1.instruction\[20\] _01485_ _01607_ vssd1 vssd1 vccd1 vccd1 _04162_
+ sky130_fd_sc_hd__and4_1
XANTENNA__10606__S net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_110_clk clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_110_clk
+ sky130_fd_sc_hd__clkbuf_8
X_06299_ _01452_ _01454_ _01456_ vssd1 vssd1 vccd1 vccd1 _01457_ sky130_fd_sc_hd__or3_1
XFILLER_0_31_245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08038_ net332 _02994_ vssd1 vssd1 vccd1 vccd1 _03177_ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_92_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold850 top.lcd.cnt_500hz\[9\] vssd1 vssd1 vccd1 vccd1 net1966 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_1832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold861 top.DUT.register\[8\]\[26\] vssd1 vssd1 vccd1 vccd1 net1977 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout975_A net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout596_X net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11010__B net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold872 top.DUT.register\[18\]\[14\] vssd1 vssd1 vccd1 vccd1 net1988 sky130_fd_sc_hd__dlygate4sd3_1
Xhold883 top.DUT.register\[24\]\[24\] vssd1 vssd1 vccd1 vccd1 net1999 sky130_fd_sc_hd__dlygate4sd3_1
Xhold894 top.DUT.register\[12\]\[8\] vssd1 vssd1 vccd1 vccd1 net2010 sky130_fd_sc_hd__dlygate4sd3_1
X_10000_ net202 net2022 net625 vssd1 vssd1 vccd1 vccd1 _00205_ sky130_fd_sc_hd__mux2_1
XANTENNA__07367__A2 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_110_Left_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06373__A_N top.a1.instruction\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06575__B1 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09989_ net231 net1854 net623 vssd1 vssd1 vccd1 vccd1 _00194_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout763_X net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10341__S net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09415__B _04471_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07119__A2 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09513__B1 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_203_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11951_ _05797_ net128 _05818_ vssd1 vssd1 vccd1 vccd1 _05834_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_106_2039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_99_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10902_ net1502 net199 net480 vssd1 vssd1 vccd1 vccd1 _01063_ sky130_fd_sc_hd__mux2_1
XFILLER_0_168_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11882_ _05710_ _05737_ _05739_ _05752_ vssd1 vssd1 vccd1 vccd1 _05765_ sky130_fd_sc_hd__and4bb_1
XANTENNA__09431__A _02155_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10833_ net1702 net231 net474 vssd1 vssd1 vccd1 vccd1 _00994_ sky130_fd_sc_hd__mux2_1
X_13621_ clknet_leaf_90_clk _01208_ net1002 vssd1 vssd1 vccd1 vccd1 net47 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_196_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09277__C1 net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08619__A2 net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10764_ net1287 net257 net485 vssd1 vssd1 vccd1 vccd1 _00925_ sky130_fd_sc_hd__mux2_1
X_13552_ clknet_leaf_104_clk _01139_ net972 vssd1 vssd1 vccd1 vccd1 top.ramload\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07827__B1 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12503_ clknet_4_6__leaf_clk _00095_ net993 vssd1 vssd1 vccd1 vccd1 top.pc\[15\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_101_1961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_564 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13483_ clknet_leaf_46_clk _01075_ net1068 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[30\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_180_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10695_ top.a1.instruction\[10\] net690 net399 _04994_ vssd1 vssd1 vccd1 vccd1 _04995_
+ sky130_fd_sc_hd__o211a_1
XANTENNA__12179__A2 net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12434_ clknet_leaf_76_clk _00030_ net1077 vssd1 vssd1 vccd1 vccd1 top.ramaddr\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_152_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_191_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08252__B1 _03367_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12365_ clknet_leaf_103_clk top.ru.next_FetchedData\[9\] net980 vssd1 vssd1 vccd1
+ vccd1 top.a1.dataIn\[9\] sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_134_2460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10516__S net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13473__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_792 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11316_ top.lcd.lcd_rs net1084 _01442_ vssd1 vssd1 vccd1 vccd1 _05201_ sky130_fd_sc_hd__and3_1
X_12296_ top.pad.count\[0\] net904 vssd1 vssd1 vccd1 vccd1 _06109_ sky130_fd_sc_hd__or2_1
XFILLER_0_120_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11247_ net880 _01382_ _05119_ vssd1 vssd1 vccd1 vccd1 _05140_ sky130_fd_sc_hd__and3_1
XANTENNA__09752__B1 _04151_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11178_ _05012_ _05024_ net473 net587 net1169 vssd1 vssd1 vccd1 vccd1 _01236_ sky130_fd_sc_hd__a32o_1
XANTENNA__06566__B1 net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10251__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10129_ net225 net1975 net609 vssd1 vssd1 vccd1 vccd1 _00329_ sky130_fd_sc_hd__mux2_1
XFILLER_0_209_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09325__B _02632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08858__A2 _03968_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11871__A top.a1.dataIn\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_203_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07530__A2 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13819_ top.lcd.lcd_en vssd1 vssd1 vccd1 vccd1 net121 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_34_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07340_ top.DUT.register\[6\]\[8\] net568 net552 top.DUT.register\[3\]\[8\] vssd1
+ vssd1 vccd1 vccd1 _02479_ sky130_fd_sc_hd__a22o_1
XFILLER_0_161_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07818__B1 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_162_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_14_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07271_ top.DUT.register\[28\]\[13\] net767 net728 top.DUT.register\[18\]\[13\] vssd1
+ vssd1 vccd1 vccd1 _02410_ sky130_fd_sc_hd__a22o_1
XFILLER_0_143_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_171_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09010_ _03180_ _03457_ _04084_ _03043_ vssd1 vssd1 vccd1 vccd1 _04085_ sky130_fd_sc_hd__and4b_1
X_06222_ net1178 net856 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedInstr\[16\] sky130_fd_sc_hd__and2_1
XFILLER_0_115_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08243__A0 _03172_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06153_ top.a1.dataIn\[16\] vssd1 vssd1 vccd1 vccd1 _01396_ sky130_fd_sc_hd__inv_2
XANTENNA__10426__S net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold102 _01166_ vssd1 vssd1 vccd1 vccd1 net1218 sky130_fd_sc_hd__dlygate4sd3_1
Xhold113 top.ramstore\[26\] vssd1 vssd1 vccd1 vccd1 net1229 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07597__A2 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold124 top.lcd.cnt_20ms\[9\] vssd1 vssd1 vccd1 vccd1 net1240 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold135 top.a1.row1\[3\] vssd1 vssd1 vccd1 vccd1 net1251 sky130_fd_sc_hd__dlygate4sd3_1
Xhold146 top.DUT.register\[6\]\[29\] vssd1 vssd1 vccd1 vccd1 net1262 sky130_fd_sc_hd__dlygate4sd3_1
Xhold157 top.DUT.register\[6\]\[12\] vssd1 vssd1 vccd1 vccd1 net1273 sky130_fd_sc_hd__dlygate4sd3_1
Xhold168 top.ramload\[3\] vssd1 vssd1 vccd1 vccd1 net1284 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09912_ top.pc\[29\] _04620_ vssd1 vssd1 vccd1 vccd1 _04919_ sky130_fd_sc_hd__nor2_1
Xhold179 top.ramaddr\[31\] vssd1 vssd1 vccd1 vccd1 net1295 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout604 net606 vssd1 vssd1 vccd1 vccd1 net604 sky130_fd_sc_hd__buf_6
XANTENNA__08546__A1 net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout615 _04954_ vssd1 vssd1 vccd1 vccd1 net615 sky130_fd_sc_hd__clkbuf_8
XANTENNA__07349__A2 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout626 _04950_ vssd1 vssd1 vccd1 vccd1 net626 sky130_fd_sc_hd__clkbuf_8
XANTENNA__09516__A top.pc\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_165_2921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09843_ _04853_ _04854_ _04856_ vssd1 vssd1 vccd1 vccd1 _04857_ sky130_fd_sc_hd__o21ai_1
Xfanout637 _01629_ vssd1 vssd1 vccd1 vccd1 net637 sky130_fd_sc_hd__clkbuf_8
Xfanout648 _01612_ vssd1 vssd1 vccd1 vccd1 net648 sky130_fd_sc_hd__clkbuf_4
Xfanout659 net662 vssd1 vssd1 vccd1 vccd1 net659 sky130_fd_sc_hd__buf_6
XANTENNA_fanout389_A net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10161__S net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09774_ _04754_ _04792_ _04794_ vssd1 vssd1 vccd1 vccd1 _04795_ sky130_fd_sc_hd__or3_1
X_06986_ top.DUT.register\[10\]\[23\] net772 _02118_ _02124_ vssd1 vssd1 vccd1 vccd1
+ _02125_ sky130_fd_sc_hd__a211o_1
XANTENNA__09950__S net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08725_ _02090_ _03841_ _03842_ _03740_ vssd1 vssd1 vccd1 vccd1 _03843_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_198_3420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11302__B1 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout556_A net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08656_ net279 _03603_ _03776_ vssd1 vssd1 vccd1 vccd1 _03777_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_205_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07521__A2 net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_54_clk_A clknet_4_12__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07607_ top.DUT.register\[13\]\[6\] net774 net655 top.DUT.register\[21\]\[6\] _02745_
+ vssd1 vssd1 vccd1 vccd1 _02746_ sky130_fd_sc_hd__a221o_1
XFILLER_0_95_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08587_ net320 _03710_ _03709_ vssd1 vssd1 vccd1 vccd1 _03711_ sky130_fd_sc_hd__a21oi_2
XANTENNA__09259__C1 net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout723_A _01630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout344_X net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_136 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07538_ _02670_ _02672_ _02674_ _02676_ vssd1 vssd1 vccd1 vccd1 _02677_ sky130_fd_sc_hd__or4_1
XFILLER_0_48_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_12_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout511_X net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07469_ _02603_ _02605_ _02607_ vssd1 vssd1 vccd1 vccd1 _02608_ sky130_fd_sc_hd__or3_1
XANTENNA_clkbuf_leaf_69_clk_A clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout609_X net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09208_ _04276_ _04277_ vssd1 vssd1 vccd1 vccd1 _04278_ sky130_fd_sc_hd__nand2_1
XFILLER_0_63_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10480_ net1698 net217 net362 vssd1 vssd1 vccd1 vccd1 _00650_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_112_clk_A clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09139_ _04211_ _04212_ vssd1 vssd1 vccd1 vccd1 _04213_ sky130_fd_sc_hd__nor2_1
XFILLER_0_161_375 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10336__S net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12150_ _06029_ _06032_ vssd1 vssd1 vccd1 vccd1 _06033_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_116_2190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06796__B1 net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11101_ net41 net865 vssd1 vssd1 vccd1 vccd1 _05056_ sky130_fd_sc_hd__and2_1
X_12081_ _05945_ _05950_ vssd1 vssd1 vccd1 vccd1 _05964_ sky130_fd_sc_hd__xor2_1
XFILLER_0_102_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold680 top.DUT.register\[5\]\[4\] vssd1 vssd1 vccd1 vccd1 net1796 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_127_clk_A clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08537__A1 net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold691 top.DUT.register\[26\]\[23\] vssd1 vssd1 vccd1 vccd1 net1807 sky130_fd_sc_hd__dlygate4sd3_1
X_11032_ net11 net841 net818 net1706 vssd1 vssd1 vccd1 vccd1 _01144_ sky130_fd_sc_hd__a22o_1
XANTENNA__08537__B2 _03663_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06402__X _01541_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10344__A1 net191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06548__B1 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10071__S net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold935_A top.ramload\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12983_ clknet_leaf_3_clk _00575_ net920 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[15\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08476__S net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11934_ _05807_ _05814_ _05815_ _05798_ _05816_ vssd1 vssd1 vccd1 vccd1 _05817_ sky130_fd_sc_hd__a221oi_4
XFILLER_0_87_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11865_ _05742_ _05747_ vssd1 vssd1 vccd1 vccd1 _05748_ sky130_fd_sc_hd__and2b_1
XANTENNA__06720__B1 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_200_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12713__CLK clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_760 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13604_ clknet_leaf_63_clk net1150 net1090 vssd1 vssd1 vccd1 vccd1 net97 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_200_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10816_ net174 net1737 net601 vssd1 vssd1 vccd1 vccd1 _00977_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11796_ _05650_ _05676_ _05648_ vssd1 vssd1 vccd1 vccd1 _05679_ sky130_fd_sc_hd__nand3b_1
XTAP_TAPCELL_ROW_31_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13535_ clknet_leaf_93_clk _01122_ net998 vssd1 vssd1 vccd1 vccd1 top.a1.data\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_131_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10747_ net1887 net187 net420 vssd1 vssd1 vccd1 vccd1 _00908_ sky130_fd_sc_hd__mux2_1
X_13466_ clknet_leaf_5_clk _01058_ net936 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[30\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_10678_ net1938 net223 net339 vssd1 vssd1 vccd1 vccd1 _00841_ sky130_fd_sc_hd__mux2_1
XANTENNA__08505__A net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_2419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12417_ clknet_leaf_110_clk top.ru.next_FetchedInstr\[29\] net989 vssd1 vssd1 vccd1
+ vccd1 top.a1.instruction\[29\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_180_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10246__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13397_ clknet_leaf_30_clk _00989_ net1019 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[28\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13225__RESET_B net1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07579__A2 net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12348_ net2090 net117 _00016_ vssd1 vssd1 vccd1 vccd1 _01373_ sky130_fd_sc_hd__mux2_1
XANTENNA__06787__B1 net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_206_Left_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12279_ top.lcd.cnt_500hz\[9\] _06097_ net686 vssd1 vssd1 vccd1 vccd1 _06098_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_120_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_208_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09725__B1 net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_310 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06840_ top.DUT.register\[14\]\[19\] net586 net521 top.DUT.register\[10\]\[19\] _01978_
+ vssd1 vssd1 vccd1 vccd1 _01979_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_147_2651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07751__A2 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06771_ top.DUT.register\[29\]\[24\] net725 _01908_ _01909_ vssd1 vssd1 vccd1 vccd1
+ _01910_ sky130_fd_sc_hd__a211o_1
XANTENNA__08914__A2_N net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08510_ net423 _03620_ _03637_ _03334_ _03635_ vssd1 vssd1 vccd1 vccd1 _03638_ sky130_fd_sc_hd__a221o_2
XTAP_TAPCELL_ROW_160_2840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_160_2851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09490_ top.a1.instruction\[24\] net822 _04470_ vssd1 vssd1 vccd1 vccd1 _04543_ sky130_fd_sc_hd__a21o_2
XANTENNA__11296__C1 _05118_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_203_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08700__A1 net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07503__A2 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08441_ _02525_ _03058_ _03061_ vssd1 vssd1 vccd1 vccd1 _03571_ sky130_fd_sc_hd__a21o_1
XFILLER_0_175_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06711__B1 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08372_ net283 _03504_ vssd1 vssd1 vccd1 vccd1 _03505_ sky130_fd_sc_hd__or2_1
XFILLER_0_19_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07323_ top.DUT.register\[9\]\[12\] net762 net726 top.DUT.register\[18\]\[12\] _02455_
+ vssd1 vssd1 vccd1 vccd1 _02462_ sky130_fd_sc_hd__a221o_1
XFILLER_0_116_512 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout137_A net139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07254_ top.DUT.register\[22\]\[13\] net576 net553 top.DUT.register\[3\]\[13\] vssd1
+ vssd1 vccd1 vccd1 _02393_ sky130_fd_sc_hd__a22o_1
XFILLER_0_171_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06205_ net887 top.ru.state\[2\] vssd1 vssd1 vccd1 vccd1 top.ru.next_iready sky130_fd_sc_hd__and2b_1
XFILLER_0_83_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_375 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07185_ top.DUT.register\[3\]\[10\] net551 net531 top.DUT.register\[12\]\[10\] vssd1
+ vssd1 vccd1 vccd1 _02324_ sky130_fd_sc_hd__a22o_1
XANTENNA__10156__S net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout304_A net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1046_A net1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_239 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09945__S net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout401 net402 vssd1 vssd1 vccd1 vccd1 net401 sky130_fd_sc_hd__buf_2
XANTENNA__11118__A3 net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07990__A2 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout423 net425 vssd1 vssd1 vccd1 vccd1 net423 sky130_fd_sc_hd__clkbuf_4
Xfanout434 _03169_ vssd1 vssd1 vccd1 vccd1 net434 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout294_X net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout445 net446 vssd1 vssd1 vccd1 vccd1 net445 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout673_A net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout456 _01553_ vssd1 vssd1 vccd1 vccd1 net456 sky130_fd_sc_hd__buf_4
X_09826_ net2152 net200 net633 vssd1 vssd1 vccd1 vccd1 _00141_ sky130_fd_sc_hd__mux2_1
Xfanout467 net470 vssd1 vssd1 vccd1 vccd1 net467 sky130_fd_sc_hd__clkbuf_8
Xfanout478 _04964_ vssd1 vssd1 vccd1 vccd1 net478 sky130_fd_sc_hd__clkbuf_8
Xfanout489 net490 vssd1 vssd1 vccd1 vccd1 net489 sky130_fd_sc_hd__buf_4
XANTENNA__07742__A2 net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout461_X net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09757_ _03682_ net405 net489 _04779_ vssd1 vssd1 vccd1 vccd1 _04780_ sky130_fd_sc_hd__o211a_1
X_06969_ top.DUT.register\[22\]\[23\] net576 net556 top.DUT.register\[28\]\[23\] vssd1
+ vssd1 vccd1 vccd1 _02108_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout559_X net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08708_ net427 _03817_ _03824_ _03168_ _03826_ vssd1 vssd1 vccd1 vccd1 _03827_ sky130_fd_sc_hd__a221oi_2
XTAP_TAPCELL_ROW_87_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09688_ _03265_ net406 net488 _04723_ vssd1 vssd1 vccd1 vccd1 _04724_ sky130_fd_sc_hd__o211a_1
XFILLER_0_96_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_178_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08639_ _02266_ _03074_ _03080_ vssd1 vssd1 vccd1 vccd1 _03761_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_96_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout726_X net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06702__B1 net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11650_ _05501_ _05512_ _05513_ _05531_ _05532_ vssd1 vssd1 vccd1 vccd1 _05533_ sky130_fd_sc_hd__o32a_1
XFILLER_0_64_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10601_ net252 net1824 net346 vssd1 vssd1 vccd1 vccd1 _00766_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11581_ _05378_ _05463_ vssd1 vssd1 vccd1 vccd1 _05464_ sky130_fd_sc_hd__xor2_1
XANTENNA__11054__A2 net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10532_ top.DUT.register\[19\]\[2\] net263 net354 vssd1 vssd1 vccd1 vccd1 _00699_
+ sky130_fd_sc_hd__mux2_1
X_13320_ clknet_leaf_27_clk _00912_ net1009 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[25\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_134_320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_796 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10066__S net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10463_ top.DUT.register\[17\]\[0\] net145 net362 vssd1 vssd1 vccd1 vccd1 _00633_
+ sky130_fd_sc_hd__mux2_1
X_13251_ clknet_leaf_57_clk _00843_ net1076 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[23\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12202_ net1290 _05978_ net688 vssd1 vssd1 vccd1 vccd1 _01309_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_114_2149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13182_ clknet_leaf_20_clk _00774_ net1029 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[21\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_10394_ _04153_ _04949_ net400 vssd1 vssd1 vccd1 vccd1 _04982_ sky130_fd_sc_hd__and3_1
XFILLER_0_103_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06769__B1 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12133_ _06001_ _06003_ _06008_ _06015_ vssd1 vssd1 vccd1 vccd1 _06016_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_19_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12689__RESET_B net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12064_ _05927_ _05928_ _05936_ vssd1 vssd1 vccd1 vccd1 _05947_ sky130_fd_sc_hd__mux2_1
X_11015_ net13 net842 net819 net1282 vssd1 vssd1 vccd1 vccd1 _01127_ sky130_fd_sc_hd__a22o_1
Xfanout990 net1007 vssd1 vssd1 vccd1 vccd1 net990 sky130_fd_sc_hd__buf_2
XANTENNA__09443__X _04499_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07733__A2 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_2381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06941__B1 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09603__B _04628_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12966_ clknet_leaf_38_clk _00558_ net1054 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[14\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_142_2570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_142_2581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11917_ _05759_ _05770_ _05777_ _05786_ vssd1 vssd1 vccd1 vccd1 _05800_ sky130_fd_sc_hd__nor4_1
XFILLER_0_185_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12897_ clknet_leaf_17_clk _00489_ net964 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[12\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_142_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_185_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11848_ _05699_ _05727_ vssd1 vssd1 vccd1 vccd1 _05731_ sky130_fd_sc_hd__xor2_1
XFILLER_0_184_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11779_ _05655_ _05656_ top.a1.dataIn\[8\] vssd1 vssd1 vccd1 vccd1 _05662_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_55_465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13518_ clknet_leaf_43_clk _01110_ net1062 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[31\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_172_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkload11 clknet_leaf_128_clk vssd1 vssd1 vccd1 vccd1 clkload11/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_125_375 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13449_ clknet_leaf_49_clk _01041_ net1061 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[29\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload22 clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 clkload22/Y sky130_fd_sc_hd__clkinv_4
Xclkload33 clknet_leaf_106_clk vssd1 vssd1 vccd1 vccd1 clkload33/Y sky130_fd_sc_hd__clkinv_8
XFILLER_0_42_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkload44 clknet_leaf_102_clk vssd1 vssd1 vccd1 vccd1 clkload44/Y sky130_fd_sc_hd__inv_12
XFILLER_0_23_351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload55 clknet_leaf_91_clk vssd1 vssd1 vccd1 vccd1 clkload55/Y sky130_fd_sc_hd__clkinv_2
XFILLER_0_2_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkload66 clknet_leaf_19_clk vssd1 vssd1 vccd1 vccd1 clkload66/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload77 clknet_leaf_38_clk vssd1 vssd1 vccd1 vccd1 clkload77/Y sky130_fd_sc_hd__inv_6
Xclkload88 clknet_leaf_56_clk vssd1 vssd1 vccd1 vccd1 clkload88/Y sky130_fd_sc_hd__inv_8
Xclkload99 clknet_leaf_77_clk vssd1 vssd1 vccd1 vccd1 clkload99/Y sky130_fd_sc_hd__clkinv_16
XFILLER_0_140_378 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10704__S net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08990_ _03824_ _03840_ _03861_ _03879_ vssd1 vssd1 vccd1 vccd1 _04065_ sky130_fd_sc_hd__and4b_1
XFILLER_0_167_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_71_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07941_ _02242_ _02262_ vssd1 vssd1 vccd1 vccd1 _03080_ sky130_fd_sc_hd__nor2_1
XANTENNA__12759__CLK clknet_leaf_128_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07872_ _03004_ _03006_ _03009_ _03010_ vssd1 vssd1 vccd1 vccd1 _03011_ sky130_fd_sc_hd__or4_1
XANTENNA__07185__B1 net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07724__A2 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09611_ top.edg2.flip1 _01394_ _04164_ vssd1 vssd1 vccd1 vccd1 _04656_ sky130_fd_sc_hd__a21oi_1
X_06823_ _01940_ _01961_ vssd1 vssd1 vccd1 vccd1 _01962_ sky130_fd_sc_hd__and2_1
XANTENNA__06932__B1 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_183_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_178_3109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06754_ top.DUT.register\[3\]\[24\] net554 net442 top.DUT.register\[5\]\[24\] _01892_
+ vssd1 vssd1 vccd1 vccd1 _01893_ sky130_fd_sc_hd__a221o_1
X_09542_ _01764_ _04590_ vssd1 vssd1 vccd1 vccd1 _04592_ sky130_fd_sc_hd__xor2_1
XANTENNA__07314__A _02443_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06685_ top.DUT.register\[16\]\[26\] net735 net725 top.DUT.register\[29\]\[26\] vssd1
+ vssd1 vccd1 vccd1 _01824_ sky130_fd_sc_hd__a22o_1
X_09473_ _04524_ _04525_ vssd1 vssd1 vccd1 vccd1 _04527_ sky130_fd_sc_hd__nor2_1
XFILLER_0_188_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout254_A _04741_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_90_clk clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_90_clk
+ sky130_fd_sc_hd__clkbuf_8
X_08424_ _03175_ _03554_ net296 vssd1 vssd1 vccd1 vccd1 _03555_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_191_3309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_82_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_191_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_82_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08355_ net885 top.pc\[5\] net696 _03488_ vssd1 vssd1 vccd1 vccd1 _03489_ sky130_fd_sc_hd__a22o_1
Xclkbuf_4_9__f_clk clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_9__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_148_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_426 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout519_A net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07306_ top.DUT.register\[25\]\[12\] net455 _02444_ vssd1 vssd1 vccd1 vccd1 _02445_
+ sky130_fd_sc_hd__a21o_1
Xclkload5 clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 clkload5/X sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_22_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08286_ _02946_ _03384_ _02945_ vssd1 vssd1 vccd1 vccd1 _03422_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_34_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06999__B1 net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07237_ _02370_ _02373_ _02374_ _02375_ vssd1 vssd1 vccd1 vccd1 _02376_ sky130_fd_sc_hd__or4_1
XFILLER_0_15_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07168_ _02286_ _02306_ vssd1 vssd1 vccd1 vccd1 _02307_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout888_A top.a1.halfData\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_570 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10614__S net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07099_ top.DUT.register\[9\]\[16\] net468 net520 top.DUT.register\[10\]\[16\] _02237_
+ vssd1 vssd1 vccd1 vccd1 _02238_ sky130_fd_sc_hd__a221o_1
XFILLER_0_100_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout220 _04766_ vssd1 vssd1 vccd1 vccd1 net220 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout231 net232 vssd1 vssd1 vccd1 vccd1 net231 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout676_X net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout242 _04745_ vssd1 vssd1 vccd1 vccd1 net242 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_208_3566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout253 _04741_ vssd1 vssd1 vccd1 vccd1 net253 sky130_fd_sc_hd__buf_2
Xfanout264 _04729_ vssd1 vssd1 vccd1 vccd1 net264 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07176__B1 net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout275 _03238_ vssd1 vssd1 vccd1 vccd1 net275 sky130_fd_sc_hd__clkbuf_2
Xfanout286 _03170_ vssd1 vssd1 vccd1 vccd1 net286 sky130_fd_sc_hd__buf_2
XANTENNA__08912__A1 _03170_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout297 net298 vssd1 vssd1 vccd1 vccd1 net297 sky130_fd_sc_hd__clkbuf_4
X_09809_ top.pc\[19\] _04471_ vssd1 vssd1 vccd1 vccd1 _04826_ sky130_fd_sc_hd__nor2_1
XANTENNA__09704__A _04716_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06923__B1 net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12820_ clknet_leaf_57_clk _00412_ net1075 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[10\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_2_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12751_ clknet_leaf_22_clk _00343_ net1021 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[7\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08039__B _02994_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_81_clk clknet_4_6__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_81_clk
+ sky130_fd_sc_hd__clkbuf_8
X_11702_ _05583_ _05584_ vssd1 vssd1 vccd1 vccd1 _05585_ sky130_fd_sc_hd__or2_1
X_12682_ clknet_leaf_115_clk _00274_ net957 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[5\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_166_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_182_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11633_ _05514_ _05515_ vssd1 vssd1 vccd1 vccd1 _05516_ sky130_fd_sc_hd__and2_1
XFILLER_0_112_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_182_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11564_ _05421_ net250 _05446_ _05445_ vssd1 vssd1 vccd1 vccd1 _05447_ sky130_fd_sc_hd__a31o_1
XFILLER_0_107_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07100__B1 net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_435 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13303_ clknet_leaf_2_clk _00895_ net919 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[25\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_10515_ net1436 net185 net358 vssd1 vssd1 vccd1 vccd1 _00684_ sky130_fd_sc_hd__mux2_1
XFILLER_0_190_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11495_ _05348_ net273 _05377_ vssd1 vssd1 vccd1 vccd1 _05378_ sky130_fd_sc_hd__a21o_1
XFILLER_0_150_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10446_ net223 net2135 net365 vssd1 vssd1 vccd1 vccd1 _00617_ sky130_fd_sc_hd__mux2_1
X_13234_ clknet_leaf_23_clk _00826_ net1022 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[23\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_150_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13165_ clknet_leaf_44_clk _00757_ net1063 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[20\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10524__S net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10377_ net1322 net188 net373 vssd1 vssd1 vccd1 vccd1 _00552_ sky130_fd_sc_hd__mux2_1
X_12116_ _05980_ _05992_ vssd1 vssd1 vccd1 vccd1 _05999_ sky130_fd_sc_hd__nand2_1
X_13096_ clknet_leaf_27_clk _00688_ net1008 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[18\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_53_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12047_ _05919_ _05929_ vssd1 vssd1 vccd1 vccd1 _05930_ sky130_fd_sc_hd__nor2_1
XANTENNA__12160__B1 top.a1.dataIn\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_144_2610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07706__A2 net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06914__B1 net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13781__D _00016_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10112__X _04956_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07405__Y _02544_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_149_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12949_ clknet_leaf_32_clk _00541_ net1044 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[14\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_29_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11266__A2 _05132_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09864__C1 _04875_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_72_clk clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_72_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_153_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08131__A2 net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06470_ net788 _01594_ _01602_ vssd1 vssd1 vccd1 vccd1 _01609_ sky130_fd_sc_hd__and3_4
XANTENNA__06973__A _02111_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_173_3039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11018__A2 net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10495__A _04712_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_508 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08140_ _02453_ net327 vssd1 vssd1 vccd1 vccd1 _03278_ sky130_fd_sc_hd__nand2_1
XFILLER_0_16_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_155_2772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08071_ _02069_ net327 vssd1 vssd1 vccd1 vccd1 _03210_ sky130_fd_sc_hd__nand2_1
Xclkload100 clknet_leaf_47_clk vssd1 vssd1 vccd1 vccd1 clkload100/Y sky130_fd_sc_hd__clkinv_2
Xclkload111 clknet_leaf_69_clk vssd1 vssd1 vccd1 vccd1 clkload111/Y sky130_fd_sc_hd__clkinv_8
XFILLER_0_43_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07022_ top.DUT.register\[13\]\[20\] net776 net712 top.DUT.register\[11\]\[20\] vssd1
+ vssd1 vccd1 vccd1 _02161_ sky130_fd_sc_hd__a22o_1
XFILLER_0_70_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_157_Left_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_140_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_188_3260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09395__A1 _02016_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_188_3271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09067__Y _04142_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10434__S net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08973_ _01697_ net692 net1147 net875 vssd1 vssd1 vccd1 vccd1 _00079_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__06213__A top.ramload\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09147__A1 net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold17 net110 vssd1 vssd1 vccd1 vccd1 net1133 sky130_fd_sc_hd__dlygate4sd3_1
Xhold28 _01174_ vssd1 vssd1 vccd1 vccd1 net1144 sky130_fd_sc_hd__dlygate4sd3_1
X_07924_ _02409_ _02429_ vssd1 vssd1 vccd1 vccd1 _03063_ sky130_fd_sc_hd__or2_1
Xhold39 _01179_ vssd1 vssd1 vccd1 vccd1 net1155 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07158__B1 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09698__A2 _01489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1009_A net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07855_ _02984_ _02993_ vssd1 vssd1 vccd1 vccd1 _02994_ sky130_fd_sc_hd__or2_4
XANTENNA_fanout371_A net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout469_A net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06806_ top.DUT.register\[27\]\[17\] net715 _01941_ _01944_ vssd1 vssd1 vccd1 vccd1
+ _01945_ sky130_fd_sc_hd__a211o_1
XPHY_EDGE_ROW_166_Left_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_84_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07786_ net823 _02904_ _02923_ vssd1 vssd1 vccd1 vccd1 _02925_ sky130_fd_sc_hd__o21a_2
XTAP_TAPCELL_ROW_203_3485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_84_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_203_3496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09525_ net134 _04575_ vssd1 vssd1 vccd1 vccd1 _04576_ sky130_fd_sc_hd__nor2_1
XFILLER_0_195_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06737_ _01853_ _01873_ vssd1 vssd1 vccd1 vccd1 _01876_ sky130_fd_sc_hd__nor2_1
XFILLER_0_211_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_63_clk clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_63_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout636_A _01629_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08122__A2 net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06668_ top.DUT.register\[4\]\[26\] net509 net442 top.DUT.register\[5\]\[26\] _01806_
+ vssd1 vssd1 vccd1 vccd1 _01807_ sky130_fd_sc_hd__a221o_1
X_09456_ top.pc\[22\] _04499_ vssd1 vssd1 vccd1 vccd1 _04511_ sky130_fd_sc_hd__or2_1
XANTENNA__07330__B1 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_148_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08407_ net275 _03524_ _03528_ _03538_ _03526_ vssd1 vssd1 vccd1 vccd1 _03539_ sky130_fd_sc_hd__a221o_1
XANTENNA__06684__A2 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07881__A1 _03019_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06599_ top.DUT.register\[26\]\[28\] net753 net733 top.DUT.register\[14\]\[28\] vssd1
+ vssd1 vccd1 vccd1 _01738_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout424_X net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout803_A _03269_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09387_ top.pc\[18\] _04428_ vssd1 vssd1 vccd1 vccd1 _04446_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10609__S net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08338_ net297 _03471_ _03469_ vssd1 vssd1 vccd1 vccd1 _03472_ sky130_fd_sc_hd__o21a_1
XFILLER_0_164_779 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_446 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08269_ _03403_ _03404_ net312 vssd1 vssd1 vccd1 vccd1 _03405_ sky130_fd_sc_hd__mux2_1
XANTENNA__11013__B net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_175_Left_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_479 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10300_ net257 net1568 net383 vssd1 vssd1 vccd1 vccd1 _00477_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11280_ net880 top.lcd.nextState\[0\] _05148_ vssd1 vssd1 vccd1 vccd1 _05170_ sky130_fd_sc_hd__and3_1
XFILLER_0_120_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_111_2108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_1874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09386__A1 net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10231_ net269 net1795 net390 vssd1 vssd1 vccd1 vccd1 _00410_ sky130_fd_sc_hd__mux2_1
XANTENNA__10344__S net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12125__A top.a1.dataIn\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07397__B1 net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_674 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10162_ net1822 net225 net602 vssd1 vssd1 vccd1 vccd1 _00361_ sky130_fd_sc_hd__mux2_1
Xfanout1004 net1005 vssd1 vssd1 vccd1 vccd1 net1004 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_7_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1015 net1016 vssd1 vssd1 vccd1 vccd1 net1015 sky130_fd_sc_hd__buf_2
Xfanout1026 net1029 vssd1 vssd1 vccd1 vccd1 net1026 sky130_fd_sc_hd__clkbuf_4
X_10093_ net1771 net207 net613 vssd1 vssd1 vccd1 vccd1 _00294_ sky130_fd_sc_hd__mux2_1
Xfanout1037 net1038 vssd1 vssd1 vccd1 vccd1 net1037 sky130_fd_sc_hd__clkbuf_4
Xfanout1048 net1071 vssd1 vssd1 vccd1 vccd1 net1048 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07149__B1 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1059 net1070 vssd1 vssd1 vccd1 vccd1 net1059 sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_184_Left_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_199_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_126_2340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_199_643 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09153__B _02857_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12803_ clknet_leaf_61_clk _00395_ net1088 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[9\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_201_124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13783_ clknet_leaf_68_clk _01352_ vssd1 vssd1 vccd1 vccd1 top.pad.button_control.r_counter\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_97_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_198_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10995_ top.a1.data\[4\] net784 vssd1 vssd1 vccd1 vccd1 _05030_ sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_54_clk clknet_4_12__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_54_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_186_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12734_ clknet_leaf_18_clk _00326_ net1030 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[7\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_32_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07321__B1 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06675__A2 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12665_ clknet_leaf_14_clk _00257_ net959 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[5\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10519__S net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11616_ net234 _05476_ _05452_ vssd1 vssd1 vccd1 vccd1 _05499_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_4_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12596_ clknet_leaf_79_clk _00188_ net1072 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[3\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11547_ _05425_ _05429_ vssd1 vssd1 vccd1 vccd1 _05430_ sky130_fd_sc_hd__nand2_1
XFILLER_0_123_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold509 top.DUT.register\[15\]\[3\] vssd1 vssd1 vccd1 vccd1 net1625 sky130_fd_sc_hd__dlygate4sd3_1
X_11478_ _01396_ net273 vssd1 vssd1 vccd1 vccd1 _05361_ sky130_fd_sc_hd__xnor2_2
Xmax_cap239 net240 vssd1 vssd1 vccd1 vccd1 net239 sky130_fd_sc_hd__clkbuf_1
X_13217_ clknet_leaf_18_clk _00809_ net1030 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[22\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_10429_ _04720_ net399 vssd1 vssd1 vccd1 vccd1 _04985_ sky130_fd_sc_hd__nand2b_1
XANTENNA__10254__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07388__B1 net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_150_2691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_162 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13148_ clknet_leaf_130_clk _00740_ net910 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[20\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_209_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13079_ clknet_leaf_129_clk _00671_ net935 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[18\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_183_3190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07640_ top.DUT.register\[15\]\[5\] net706 net698 top.DUT.register\[31\]\[5\] vssd1
+ vssd1 vccd1 vccd1 _02779_ sky130_fd_sc_hd__a22o_1
XFILLER_0_73_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07560__B1 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13492__RESET_B net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07571_ top.DUT.register\[29\]\[6\] net451 net507 top.DUT.register\[4\]\[6\] _02709_
+ vssd1 vssd1 vccd1 vccd1 _02710_ sky130_fd_sc_hd__a221o_1
XFILLER_0_177_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_66_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_45_clk clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_45_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_66_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06522_ top.DUT.register\[18\]\[29\] net549 net454 top.DUT.register\[29\]\[29\] _01660_
+ vssd1 vssd1 vccd1 vccd1 _01661_ sky130_fd_sc_hd__a221o_1
X_09310_ _04368_ _04373_ vssd1 vssd1 vccd1 vccd1 _04374_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_24_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07312__B1 net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_157_2801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06453_ top.a1.instruction\[24\] net792 vssd1 vssd1 vccd1 vccd1 _01592_ sky130_fd_sc_hd__nand2_1
X_09241_ net136 _04297_ _04308_ vssd1 vssd1 vccd1 vccd1 _04309_ sky130_fd_sc_hd__o21ai_1
XANTENNA__06666__A2 net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_200_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_146_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09172_ net134 _04243_ vssd1 vssd1 vccd1 vccd1 _04244_ sky130_fd_sc_hd__nor2_1
X_06384_ top.a1.instruction\[16\] _01522_ vssd1 vssd1 vccd1 vccd1 _01523_ sky130_fd_sc_hd__and2b_2
XANTENNA__06208__A top.ramload\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_267 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08123_ net436 _03176_ _03188_ _03261_ _03166_ vssd1 vssd1 vccd1 vccd1 _03262_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_44_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06418__A2 net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10953__A top.a1.halfData\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08054_ _01572_ net330 vssd1 vssd1 vccd1 vccd1 _03193_ sky130_fd_sc_hd__nor2_1
XFILLER_0_31_427 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_596 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09519__A net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07091__A2 net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07005_ top.DUT.register\[19\]\[20\] net537 net461 top.DUT.register\[17\]\[20\] _02143_
+ vssd1 vssd1 vccd1 vccd1 _02144_ sky130_fd_sc_hd__a221o_1
XFILLER_0_3_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_96 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10164__S net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07379__B1 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07039__A _02155_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09953__S net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07918__A2 _02703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08710__X _03829_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout586_A _01513_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_168_2963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08956_ net1202 net874 _02472_ net693 vssd1 vssd1 vccd1 vccd1 _00062_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_4_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_205_3514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_205_3525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07907_ _03021_ _03040_ _03045_ vssd1 vssd1 vccd1 vccd1 _03046_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout753_A _01621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08887_ net306 _03996_ vssd1 vssd1 vccd1 vccd1 _03997_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout374_X net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09540__A1 top.a1.instruction\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07838_ top.DUT.register\[16\]\[0\] net546 net516 top.DUT.register\[7\]\[0\] _02976_
+ vssd1 vssd1 vccd1 vccd1 _02977_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_108_2070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07551__B1 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07769_ top.DUT.register\[13\]\[2\] net774 net770 top.DUT.register\[10\]\[2\] vssd1
+ vssd1 vccd1 vccd1 _02908_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout541_X net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_36_clk clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_36_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout639_X net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13162__RESET_B net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09508_ top.a1.instruction\[25\] net821 net422 vssd1 vssd1 vccd1 vccd1 _04560_ sky130_fd_sc_hd__a21o_2
XFILLER_0_195_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10780_ net1381 net202 net485 vssd1 vssd1 vccd1 vccd1 _00941_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07303__B1 net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10989__B2 top.a1.dataIn\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06657__A2 net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_426 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09439_ _04482_ _04483_ _04484_ vssd1 vssd1 vccd1 vccd1 _04495_ sky130_fd_sc_hd__o21a_1
XANTENNA__10339__S net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_192_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12450_ clknet_leaf_75_clk _00046_ net1081 vssd1 vssd1 vccd1 vccd1 top.ramaddr\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_164_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_1903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11401_ _05249_ _05283_ vssd1 vssd1 vccd1 vccd1 _05284_ sky130_fd_sc_hd__and2_1
XFILLER_0_136_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12381_ clknet_leaf_110_clk top.ru.next_FetchedData\[25\] net989 vssd1 vssd1 vccd1
+ vccd1 top.a1.dataIn\[25\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_7_690 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11332_ _05204_ _05208_ vssd1 vssd1 vccd1 vccd1 _05215_ sky130_fd_sc_hd__and2b_1
XANTENNA__13102__CLK clknet_leaf_40_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06290__B1 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10074__S net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11263_ top.a1.row2\[25\] _05142_ _05145_ top.a1.row2\[17\] vssd1 vssd1 vccd1 vccd1
+ _05155_ sky130_fd_sc_hd__a22o_1
XFILLER_0_104_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13002_ clknet_leaf_116_clk _00594_ net958 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[15\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07909__A2 _02944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10214_ net217 net2222 net396 vssd1 vssd1 vccd1 vccd1 _00394_ sky130_fd_sc_hd__mux2_1
X_11194_ _01407_ net588 _04668_ vssd1 vssd1 vccd1 vccd1 _01247_ sky130_fd_sc_hd__a21oi_1
X_10145_ top.a1.instruction\[11\] _04711_ _04719_ vssd1 vssd1 vccd1 vccd1 _04957_
+ sky130_fd_sc_hd__nor3_4
XANTENNA__08582__A2 net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_192_Left_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10802__S net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07790__B1 net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07383__S net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10076_ net2301 net154 net618 vssd1 vssd1 vccd1 vccd1 _00278_ sky130_fd_sc_hd__mux2_1
XANTENNA__07542__B1 net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06896__A2 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_27_clk clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_27_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_202_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13766_ clknet_leaf_100_clk _01337_ vssd1 vssd1 vccd1 vccd1 top.lcd.cnt_500hz\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_48_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10978_ net1141 _05017_ net589 vssd1 vssd1 vccd1 vccd1 _01117_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_806 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12717_ clknet_leaf_51_clk _00309_ net1035 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[6\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10249__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_183_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13697_ clknet_leaf_73_clk _01268_ vssd1 vssd1 vccd1 vccd1 net113 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_139_2531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12648_ clknet_leaf_7_clk _00240_ net946 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[4\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_61_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_152_2720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12579_ clknet_leaf_61_clk _00171_ net1088 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[2\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_142_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_152_2731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_382 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07073__A2 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold306 top.DUT.register\[30\]\[8\] vssd1 vssd1 vccd1 vccd1 net1422 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_235 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold317 top.DUT.register\[11\]\[8\] vssd1 vssd1 vccd1 vccd1 net1433 sky130_fd_sc_hd__dlygate4sd3_1
Xhold328 top.DUT.register\[18\]\[9\] vssd1 vssd1 vccd1 vccd1 net1444 sky130_fd_sc_hd__dlygate4sd3_1
Xhold339 top.DUT.register\[27\]\[0\] vssd1 vssd1 vccd1 vccd1 net1455 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06820__A2 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08022__A1 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout808 net809 vssd1 vssd1 vccd1 vccd1 net808 sky130_fd_sc_hd__buf_2
XFILLER_0_0_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout819 _05043_ vssd1 vssd1 vccd1 vccd1 net819 sky130_fd_sc_hd__clkbuf_2
X_08810_ _01878_ net495 _03923_ vssd1 vssd1 vccd1 vccd1 _03924_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10712__S net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09790_ _04806_ _04807_ _04808_ vssd1 vssd1 vccd1 vccd1 _04809_ sky130_fd_sc_hd__or3_1
Xhold1006 top.DUT.register\[14\]\[19\] vssd1 vssd1 vccd1 vccd1 net2122 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07781__B1 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1017 top.DUT.register\[20\]\[3\] vssd1 vssd1 vccd1 vccd1 net2133 sky130_fd_sc_hd__dlygate4sd3_1
X_08741_ net277 _03209_ _03215_ _03857_ vssd1 vssd1 vccd1 vccd1 _03858_ sky130_fd_sc_hd__a31o_1
XPHY_EDGE_ROW_183_Right_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1028 top.DUT.register\[28\]\[14\] vssd1 vssd1 vccd1 vccd1 net2144 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1039 top.DUT.register\[6\]\[9\] vssd1 vssd1 vccd1 vccd1 net2155 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13602__RESET_B net1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_206_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_61 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08672_ net318 _03428_ vssd1 vssd1 vccd1 vccd1 _03792_ sky130_fd_sc_hd__or2_1
XANTENNA__06210__B net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_163_2893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07533__B1 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_205_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07623_ top.DUT.register\[6\]\[5\] net567 net463 top.DUT.register\[13\]\[5\] _02761_
+ vssd1 vssd1 vccd1 vccd1 _02762_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_5_Right_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_419 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_200_3444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_18_clk clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_18_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout167_A _04895_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_679 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07554_ _02685_ _02686_ _02691_ _02692_ vssd1 vssd1 vccd1 vccd1 _02693_ sky130_fd_sc_hd__or4_1
XANTENNA__09521__B _04560_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_196_3381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09825__A2 net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_196_3392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06505_ top.DUT.register\[23\]\[30\] net673 net752 top.DUT.register\[26\]\[30\] _01639_
+ vssd1 vssd1 vccd1 vccd1 _01644_ sky130_fd_sc_hd__a221o_1
XANTENNA__06639__A2 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07485_ top.DUT.register\[15\]\[14\] net681 net677 top.DUT.register\[31\]\[14\] vssd1
+ vssd1 vccd1 vccd1 _02624_ sky130_fd_sc_hd__a22o_1
XANTENNA__10159__S net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07836__A1 _02973_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_192_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_174_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout334_A net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1076_A net1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09224_ _04276_ _04280_ _04292_ vssd1 vssd1 vccd1 vccd1 _04293_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09948__S net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06436_ top.a1.instruction\[6\] _01472_ _01573_ vssd1 vssd1 vccd1 vccd1 _01575_ sky130_fd_sc_hd__or3_1
XFILLER_0_173_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06367_ _01388_ _01503_ vssd1 vssd1 vccd1 vccd1 _01506_ sky130_fd_sc_hd__nand2_1
X_09155_ _04226_ _04227_ vssd1 vssd1 vccd1 vccd1 _04228_ sky130_fd_sc_hd__nand2_1
XFILLER_0_134_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout501_A net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_563 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_79_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08106_ _02453_ net299 vssd1 vssd1 vccd1 vccd1 _03245_ sky130_fd_sc_hd__nand2_1
XFILLER_0_140_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07064__A2 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09086_ top.a1.instruction\[28\] top.a1.instruction\[29\] top.a1.instruction\[30\]
+ top.a1.instruction\[31\] vssd1 vssd1 vccd1 vccd1 _04161_ sky130_fd_sc_hd__and4_1
XFILLER_0_71_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06298_ _01332_ _01333_ vssd1 vssd1 vccd1 vccd1 _01456_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_114_462 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08037_ net283 _03175_ vssd1 vssd1 vccd1 vccd1 _03176_ sky130_fd_sc_hd__nor2_1
XFILLER_0_3_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06811__A2 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold840 top.DUT.register\[27\]\[11\] vssd1 vssd1 vccd1 vccd1 net1956 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_1833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold851 top.DUT.register\[7\]\[31\] vssd1 vssd1 vccd1 vccd1 net1967 sky130_fd_sc_hd__dlygate4sd3_1
Xhold862 top.DUT.register\[21\]\[4\] vssd1 vssd1 vccd1 vccd1 net1978 sky130_fd_sc_hd__dlygate4sd3_1
Xhold873 top.DUT.register\[2\]\[11\] vssd1 vssd1 vccd1 vccd1 net1989 sky130_fd_sc_hd__dlygate4sd3_1
Xhold884 top.DUT.register\[25\]\[16\] vssd1 vssd1 vccd1 vccd1 net2000 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout491_X net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold895 top.DUT.register\[24\]\[27\] vssd1 vssd1 vccd1 vccd1 net2011 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09761__A1 top.pc\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10622__S net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09988_ net236 net1868 net626 vssd1 vssd1 vccd1 vccd1 _00193_ sky130_fd_sc_hd__mux2_1
XANTENNA__07772__B1 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08600__B _03720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08939_ _04028_ _04045_ vssd1 vssd1 vccd1 vccd1 _04047_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout756_X net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_150_Right_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11950_ net128 _05818_ _05797_ vssd1 vssd1 vccd1 vccd1 _05833_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_106_2029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07524__B1 net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11320__A1 top.a1.dataIn\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09712__A net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10901_ net2123 net209 net480 vssd1 vssd1 vccd1 vccd1 _01062_ sky130_fd_sc_hd__mux2_1
XFILLER_0_196_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06878__A2 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11881_ _05739_ _05752_ vssd1 vssd1 vccd1 vccd1 _05764_ sky130_fd_sc_hd__nand2_2
XFILLER_0_86_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13620_ clknet_leaf_89_clk _01207_ net1002 vssd1 vssd1 vccd1 vccd1 net46 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_196_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10832_ net1369 net236 net474 vssd1 vssd1 vccd1 vccd1 _00993_ sky130_fd_sc_hd__mux2_1
XANTENNA__09431__B _04487_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_115 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13551_ clknet_leaf_104_clk _01138_ net973 vssd1 vssd1 vccd1 vccd1 top.ramload\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_13_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10069__S net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10763_ net1644 net259 net484 vssd1 vssd1 vccd1 vccd1 _00924_ sky130_fd_sc_hd__mux2_1
XFILLER_0_165_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_183_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12502_ clknet_leaf_111_clk _00094_ net990 vssd1 vssd1 vccd1 vccd1 top.pc\[14\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_81_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_192_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13482_ clknet_leaf_117_clk _01074_ net958 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[30\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_101_1962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_576 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_671 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10694_ top.a1.instruction\[11\] _04711_ _04719_ vssd1 vssd1 vccd1 vccd1 _04994_
+ sky130_fd_sc_hd__or3b_1
XFILLER_0_81_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12433_ clknet_leaf_85_clk _00029_ net1001 vssd1 vssd1 vccd1 vccd1 top.ramaddr\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_43_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07055__A2 net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08252__A1 net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12364_ clknet_leaf_102_clk top.ru.next_FetchedData\[8\] net980 vssd1 vssd1 vccd1
+ vccd1 top.a1.dataIn\[8\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_23_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_134_2450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_134_2461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11315_ net1196 net813 _05200_ net1082 vssd1 vssd1 vccd1 vccd1 _01271_ sky130_fd_sc_hd__o211a_1
XANTENNA__06802__A2 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12295_ top.pad.count\[0\] net904 vssd1 vssd1 vccd1 vccd1 _06108_ sky130_fd_sc_hd__nand2_1
X_11246_ net878 _05118_ _05120_ vssd1 vssd1 vccd1 vccd1 _05139_ sky130_fd_sc_hd__and3_1
XANTENNA__08555__A2 net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10532__S net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11177_ _05007_ _05021_ net473 net587 net1192 vssd1 vssd1 vccd1 vccd1 _01235_ sky130_fd_sc_hd__a32o_1
X_10128_ net188 net1950 net607 vssd1 vssd1 vccd1 vccd1 _00328_ sky130_fd_sc_hd__mux2_1
XANTENNA__09325__C _04386_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10059_ net1585 net212 net615 vssd1 vssd1 vccd1 vccd1 _00261_ sky130_fd_sc_hd__mux2_1
XFILLER_0_199_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06869__A2 net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_187_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_159_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13818_ net1103 vssd1 vssd1 vccd1 vccd1 gpio_out[5] sky130_fd_sc_hd__buf_2
XFILLER_0_203_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_34_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13749_ clknet_leaf_99_clk net1241 vssd1 vssd1 vccd1 vccd1 top.lcd.cnt_20ms\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_161_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07270_ _02399_ _02408_ vssd1 vssd1 vccd1 vccd1 _02409_ sky130_fd_sc_hd__nor2_4
XTAP_TAPCELL_ROW_14_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11090__A3 net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06221_ net1204 net856 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedInstr\[15\] sky130_fd_sc_hd__and2_1
XFILLER_0_155_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10707__S net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_360 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06152_ top.a1.dataIn\[18\] vssd1 vssd1 vccd1 vccd1 _01395_ sky130_fd_sc_hd__inv_2
XANTENNA__07046__A2 net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold103 top.a1.row1\[11\] vssd1 vssd1 vccd1 vccd1 net1219 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10050__A1 net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold114 _01186_ vssd1 vssd1 vccd1 vccd1 net1230 sky130_fd_sc_hd__dlygate4sd3_1
Xhold125 _01320_ vssd1 vssd1 vccd1 vccd1 net1241 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold136 top.a1.row1\[16\] vssd1 vssd1 vccd1 vccd1 net1252 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_98 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_7_clk clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_7_clk
+ sky130_fd_sc_hd__clkbuf_8
Xhold147 top.a1.row1\[114\] vssd1 vssd1 vccd1 vccd1 net1263 sky130_fd_sc_hd__dlygate4sd3_1
Xhold158 top.ramload\[5\] vssd1 vssd1 vccd1 vccd1 net1274 sky130_fd_sc_hd__dlygate4sd3_1
X_09911_ top.pc\[29\] _04620_ vssd1 vssd1 vccd1 vccd1 _04918_ sky130_fd_sc_hd__and2_1
Xhold169 top.a1.data\[6\] vssd1 vssd1 vccd1 vccd1 net1285 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_74_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout605 net606 vssd1 vssd1 vccd1 vccd1 net605 sky130_fd_sc_hd__buf_4
XANTENNA__08529__A2_N _03653_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout616 _04954_ vssd1 vssd1 vccd1 vccd1 net616 sky130_fd_sc_hd__clkbuf_4
Xfanout627 _04948_ vssd1 vssd1 vccd1 vccd1 net627 sky130_fd_sc_hd__clkbuf_8
XANTENNA__09075__Y _04150_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10442__S net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09842_ net828 _04508_ _04855_ vssd1 vssd1 vccd1 vccd1 _04856_ sky130_fd_sc_hd__o21ba_1
Xfanout638 _01629_ vssd1 vssd1 vccd1 vccd1 net638 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_165_2922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout649 _01612_ vssd1 vssd1 vccd1 vccd1 net649 sky130_fd_sc_hd__clkbuf_8
XANTENNA__07754__B1 net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09773_ _04403_ _04776_ _04793_ net799 vssd1 vssd1 vccd1 vccd1 _04794_ sky130_fd_sc_hd__a22o_1
X_06985_ top.DUT.register\[5\]\[23\] net653 net752 top.DUT.register\[26\]\[23\] _02123_
+ vssd1 vssd1 vccd1 vccd1 _02124_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout284_A _03170_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08724_ _02091_ net501 vssd1 vssd1 vccd1 vccd1 _03842_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_198_3410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_198_3421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07506__B1 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08655_ net324 _03387_ _03775_ net283 vssd1 vssd1 vccd1 vccd1 _03776_ sky130_fd_sc_hd__o22a_1
XFILLER_0_178_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout451_A _01561_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout549_A net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11292__B1_N _05121_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07606_ top.DUT.register\[16\]\[6\] net734 net722 top.DUT.register\[29\]\[6\] vssd1
+ vssd1 vccd1 vccd1 _02745_ sky130_fd_sc_hd__a22o_1
X_08586_ _03333_ _03426_ vssd1 vssd1 vccd1 vccd1 _03710_ sky130_fd_sc_hd__or2_1
XANTENNA__08148__A _02849_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07537_ top.DUT.register\[14\]\[7\] net583 net451 top.DUT.register\[29\]\[7\] _02675_
+ vssd1 vssd1 vccd1 vccd1 _02676_ sky130_fd_sc_hd__a221o_1
XFILLER_0_147_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout716_A net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout337_X net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07468_ top.DUT.register\[4\]\[15\] net668 net663 top.DUT.register\[20\]\[15\] _02606_
+ vssd1 vssd1 vccd1 vccd1 _02607_ sky130_fd_sc_hd__a221o_1
XANTENNA__07285__A2 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08482__A1 net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08482__B2 net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06493__B1 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09207_ _02678_ _02682_ vssd1 vssd1 vccd1 vccd1 _04277_ sky130_fd_sc_hd__or2_1
X_06419_ net683 _01516_ _01518_ vssd1 vssd1 vccd1 vccd1 _01558_ sky130_fd_sc_hd__and3_4
XFILLER_0_8_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10617__S net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout504_X net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07399_ top.DUT.register\[24\]\[9\] net511 _02535_ _02537_ vssd1 vssd1 vccd1 vccd1
+ _02538_ sky130_fd_sc_hd__a211o_1
XFILLER_0_161_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07037__A2 _02175_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09138_ top.pc\[3\] _02904_ vssd1 vssd1 vccd1 vccd1 _04212_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_32_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_161_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_116_2180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09069_ _01477_ _01485_ _01588_ _02336_ _04143_ vssd1 vssd1 vccd1 vccd1 _04144_ sky130_fd_sc_hd__o32a_1
XTAP_TAPCELL_ROW_116_2191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11100_ net905 net1874 net860 _05055_ vssd1 vssd1 vccd1 vccd1 _01201_ sky130_fd_sc_hd__a31o_1
XANTENNA__07993__B1 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09707__A net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12080_ _05945_ _05950_ vssd1 vssd1 vccd1 vccd1 _05963_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout873_X net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold670 top.DUT.register\[4\]\[24\] vssd1 vssd1 vccd1 vccd1 net1786 sky130_fd_sc_hd__dlygate4sd3_1
Xhold681 top.DUT.register\[5\]\[30\] vssd1 vssd1 vccd1 vccd1 net1797 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08537__A2 top.pc\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold692 top.DUT.register\[7\]\[24\] vssd1 vssd1 vccd1 vccd1 net1808 sky130_fd_sc_hd__dlygate4sd3_1
X_11031_ net10 net841 net818 net1278 vssd1 vssd1 vccd1 vccd1 _01143_ sky130_fd_sc_hd__a22o_1
XANTENNA__10352__S net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09426__B _04471_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07745__B1 net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12982_ clknet_leaf_3_clk _00574_ net920 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[15\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09498__B1 _04051_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input12_A DAT_I[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11933_ _05805_ _05808_ _05813_ vssd1 vssd1 vccd1 vccd1 _05816_ sky130_fd_sc_hd__and3b_1
XFILLER_0_169_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_196_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_197_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11864_ _05744_ _05746_ vssd1 vssd1 vccd1 vccd1 _05747_ sky130_fd_sc_hd__xnor2_1
XANTENNA__08058__A _01764_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13603_ clknet_leaf_65_clk net1137 net1094 vssd1 vssd1 vccd1 vccd1 net96 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_45_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11057__B1 _05045_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10815_ net177 net1800 net601 vssd1 vssd1 vccd1 vccd1 _00976_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11795_ _05668_ _05672_ _05674_ _05677_ _05650_ vssd1 vssd1 vccd1 vccd1 _05678_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_82_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_200_789 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_31_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13534_ clknet_leaf_92_clk _01121_ net995 vssd1 vssd1 vccd1 vccd1 top.a1.data\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_10746_ net1656 net204 net420 vssd1 vssd1 vccd1 vccd1 _00907_ sky130_fd_sc_hd__mux2_1
XFILLER_0_40_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07276__A2 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09670__B1 top.pc\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13465_ clknet_leaf_16_clk _01057_ net960 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[30\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10527__S net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10677_ net1509 net191 net340 vssd1 vssd1 vccd1 vccd1 _00840_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12416_ clknet_leaf_111_clk top.ru.next_FetchedInstr\[28\] net989 vssd1 vssd1 vccd1
+ vccd1 top.a1.instruction\[28\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_125_579 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13396_ clknet_leaf_55_clk _00988_ net1072 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[28\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12347_ net2295 _01408_ net38 vssd1 vssd1 vccd1 vccd1 _01372_ sky130_fd_sc_hd__a21o_1
XFILLER_0_105_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07984__B1 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12278_ _06097_ net687 _06096_ vssd1 vssd1 vccd1 vccd1 _01343_ sky130_fd_sc_hd__and3b_1
XFILLER_0_120_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13265__RESET_B net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09725__A1 top.a1.dataIn\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11229_ top.lcd.nextState\[5\] top.lcd.nextState\[4\] vssd1 vssd1 vccd1 vccd1 _05122_
+ sky130_fd_sc_hd__and2b_1
XFILLER_0_4_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07736__B1 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_207_322 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_147_2652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09623__Y _04668_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06770_ top.DUT.register\[9\]\[24\] net764 net756 top.DUT.register\[1\]\[24\] _01907_
+ vssd1 vssd1 vccd1 vccd1 _01909_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_160_2841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_160_2852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12538__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08440_ net1631 net833 net803 _03570_ vssd1 vssd1 vccd1 vccd1 _00026_ sky130_fd_sc_hd__a22o_1
XFILLER_0_81_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08371_ _03380_ _03503_ net309 vssd1 vssd1 vccd1 vccd1 _03504_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_193_3340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07322_ top.DUT.register\[22\]\[12\] net647 net742 top.DUT.register\[2\]\[12\] _02460_
+ vssd1 vssd1 vccd1 vccd1 _02461_ sky130_fd_sc_hd__a221o_1
XFILLER_0_45_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07267__A2 net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07253_ top.DUT.register\[24\]\[13\] net513 net453 top.DUT.register\[29\]\[13\] _02391_
+ vssd1 vssd1 vccd1 vccd1 _02392_ sky130_fd_sc_hd__a221o_1
XFILLER_0_171_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10437__S net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06204_ top.Wen wb.curr_state\[0\] _01387_ wb.curr_state\[2\] net905 vssd1 vssd1
+ vccd1 vccd1 _00015_ sky130_fd_sc_hd__a32o_1
XFILLER_0_116_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07019__A2 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07184_ top.DUT.register\[20\]\[10\] net563 net443 top.DUT.register\[1\]\[10\] _02322_
+ vssd1 vssd1 vccd1 vccd1 _02323_ sky130_fd_sc_hd__a221o_1
XFILLER_0_171_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_207 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08216__B2 _03353_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07975__B1 net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1039_A net1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09527__A _01810_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06503__X _01642_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout402 _04802_ vssd1 vssd1 vccd1 vccd1 net402 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08519__A2 net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout499_A net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10172__S net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout424 net425 vssd1 vssd1 vccd1 vccd1 net424 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08150__B _03040_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout435 net436 vssd1 vssd1 vccd1 vccd1 net435 sky130_fd_sc_hd__buf_2
XANTENNA__07727__B1 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09961__S net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout446 _01564_ vssd1 vssd1 vccd1 vccd1 net446 sky130_fd_sc_hd__buf_4
Xfanout457 net458 vssd1 vssd1 vccd1 vccd1 net457 sky130_fd_sc_hd__clkbuf_8
XANTENNA_input4_A DAT_I[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13313__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09825_ _03829_ net405 net489 _04840_ vssd1 vssd1 vccd1 vccd1 _04841_ sky130_fd_sc_hd__o211a_4
Xfanout468 net470 vssd1 vssd1 vccd1 vccd1 net468 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout666_A _01605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout479 _04964_ vssd1 vssd1 vccd1 vccd1 net479 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10900__S net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09756_ _04370_ _04776_ _04778_ _04754_ vssd1 vssd1 vccd1 vccd1 _04779_ sky130_fd_sc_hd__a211o_1
X_06968_ top.DUT.register\[7\]\[23\] net516 net444 top.DUT.register\[1\]\[23\] _02106_
+ vssd1 vssd1 vccd1 vccd1 _02107_ sky130_fd_sc_hd__a221o_1
X_08707_ net323 net429 _03441_ _03825_ vssd1 vssd1 vccd1 vccd1 _03826_ sky130_fd_sc_hd__a31o_1
X_09687_ top.a1.dataIn\[0\] net795 _04722_ top.pc\[0\] net407 vssd1 vssd1 vccd1 vccd1
+ _04723_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_87_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06899_ top.DUT.register\[25\]\[18\] net780 net748 top.DUT.register\[17\]\[18\] vssd1
+ vssd1 vccd1 vccd1 _02038_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout454_X net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout833_A _01499_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13463__CLK clknet_leaf_128_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08638_ _03264_ _03749_ _03759_ net435 vssd1 vssd1 vccd1 vccd1 _03760_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_166_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12396__Q top.a1.instruction\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08569_ _03171_ _03492_ _03496_ net280 vssd1 vssd1 vccd1 vccd1 _03694_ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout621_X net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_0__f_clk_A clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10695__X _04995_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_608 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout719_X net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10600_ net255 net1978 net348 vssd1 vssd1 vccd1 vccd1 _00765_ sky130_fd_sc_hd__mux2_1
XFILLER_0_166_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07258__A2 net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11580_ _05409_ _05415_ _05430_ net249 _05402_ vssd1 vssd1 vccd1 vccd1 _05463_ sky130_fd_sc_hd__a41o_1
XFILLER_0_64_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08606__A net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_2220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10531_ net2028 net269 net355 vssd1 vssd1 vccd1 vccd1 _00698_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10347__S net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_691 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13250_ clknet_leaf_26_clk _00842_ net1009 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[23\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_10462_ _04712_ _04713_ net400 vssd1 vssd1 vccd1 vccd1 _04986_ sky130_fd_sc_hd__and3_1
XFILLER_0_17_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout990_X net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12201_ net1138 _05992_ net688 vssd1 vssd1 vccd1 vccd1 _01308_ sky130_fd_sc_hd__mux2_1
XANTENNA__10014__A1 net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09955__A1 net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13181_ clknet_leaf_119_clk _00773_ net931 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[21\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_10393_ net1780 net142 net375 vssd1 vssd1 vccd1 vccd1 _00568_ sky130_fd_sc_hd__mux2_1
XANTENNA__07966__B1 net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12132_ _05983_ _05992_ _05999_ _05982_ vssd1 vssd1 vccd1 vccd1 _06015_ sky130_fd_sc_hd__a22o_1
XFILLER_0_32_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06413__X _01552_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12063_ _05938_ _05939_ _05945_ vssd1 vssd1 vccd1 vccd1 _05946_ sky130_fd_sc_hd__o21a_1
XANTENNA__10082__S net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11014_ net2 net840 _05044_ net1793 vssd1 vssd1 vccd1 vccd1 _01126_ sky130_fd_sc_hd__o22a_1
XANTENNA__09724__X _04752_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08995__B _04020_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout980 net987 vssd1 vssd1 vccd1 vccd1 net980 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10810__S net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout991 net993 vssd1 vssd1 vccd1 vccd1 net991 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_129_2382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07244__X _02383_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09172__A net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_204_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12965_ clknet_leaf_35_clk _00557_ net1041 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[14\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_99_363 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13690__Q top.lcd.nextState\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11916_ _05759_ _05770_ _05776_ _05786_ _05773_ vssd1 vssd1 vccd1 vccd1 _05799_ sky130_fd_sc_hd__o41a_1
XFILLER_0_87_547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_142_2571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07497__A2 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_142_2582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12896_ clknet_leaf_114_clk _00488_ net963 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[12\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_68_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11847_ top.a1.dataIn\[5\] _05727_ _05728_ vssd1 vssd1 vccd1 vccd1 _05730_ sky130_fd_sc_hd__or3_1
XFILLER_0_142_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_200_575 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_185_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_175_3070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_660 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11778_ _05628_ _05657_ _05658_ _05660_ vssd1 vssd1 vccd1 vccd1 _05661_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_126_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13517_ clknet_leaf_44_clk _01109_ net1063 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[31\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10257__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10729_ net1804 net267 net419 vssd1 vssd1 vccd1 vccd1 _00890_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkload12 clknet_leaf_129_clk vssd1 vssd1 vccd1 vccd1 clkload12/Y sky130_fd_sc_hd__inv_6
X_13448_ clknet_leaf_27_clk _01040_ net1009 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[29\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_180_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkload23 clknet_leaf_11_clk vssd1 vssd1 vccd1 vccd1 clkload23/Y sky130_fd_sc_hd__inv_6
XFILLER_0_153_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkload34 clknet_leaf_107_clk vssd1 vssd1 vccd1 vccd1 clkload34/Y sky130_fd_sc_hd__inv_16
XTAP_TAPCELL_ROW_58_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08749__A2 net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload45 clknet_leaf_80_clk vssd1 vssd1 vccd1 vccd1 clkload45/Y sky130_fd_sc_hd__inv_6
XFILLER_0_23_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_58_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload56 clknet_leaf_92_clk vssd1 vssd1 vccd1 vccd1 clkload56/Y sky130_fd_sc_hd__clkinv_2
X_13379_ clknet_leaf_49_clk _00971_ net1061 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[27\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload67 clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 clkload67/Y sky130_fd_sc_hd__inv_6
Xclkload78 clknet_leaf_39_clk vssd1 vssd1 vccd1 vccd1 clkload78/Y sky130_fd_sc_hd__inv_6
Xclkload89 clknet_leaf_57_clk vssd1 vssd1 vccd1 vccd1 clkload89/Y sky130_fd_sc_hd__clkinv_4
XANTENNA_clkbuf_leaf_53_clk_A clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07421__A2 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_4_11__f_clk_A clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07940_ _02007_ _03078_ _03075_ vssd1 vssd1 vccd1 vccd1 _03079_ sky130_fd_sc_hd__a21oi_1
X_07871_ top.DUT.register\[25\]\[1\] net780 net767 top.DUT.register\[28\]\[1\] _03007_
+ vssd1 vssd1 vccd1 vccd1 _03010_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_79_Left_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08382__B1 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09610_ net902 top.pc\[31\] _04647_ _04655_ net890 vssd1 vssd1 vccd1 vccd1 _00111_
+ sky130_fd_sc_hd__o221a_1
XANTENNA_clkbuf_leaf_68_clk_A clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06822_ net807 _01960_ net437 vssd1 vssd1 vccd1 vccd1 _01961_ sky130_fd_sc_hd__o21a_1
XANTENNA__10720__S net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_111_clk_A clknet_4_6__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09541_ _01754_ _01763_ _04590_ vssd1 vssd1 vccd1 vccd1 _04591_ sky130_fd_sc_hd__o21a_1
X_06753_ top.DUT.register\[6\]\[24\] net570 net566 top.DUT.register\[20\]\[24\] vssd1
+ vssd1 vccd1 vccd1 _01892_ sky130_fd_sc_hd__a22o_1
XFILLER_0_78_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09331__C1 net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_69_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07314__B _02452_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07488__A2 net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09472_ _04524_ _04525_ vssd1 vssd1 vccd1 vccd1 _04526_ sky130_fd_sc_hd__and2_1
X_06684_ top.DUT.register\[25\]\[26\] net781 _01812_ _01822_ vssd1 vssd1 vccd1 vccd1
+ _01823_ sky130_fd_sc_hd__a211o_1
XFILLER_0_78_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08423_ _03452_ _03553_ net308 vssd1 vssd1 vccd1 vccd1 _03554_ sky130_fd_sc_hd__mux2_1
XANTENNA__06696__B1 net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10956__A _04657_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_126_clk_A clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout247_A _04749_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_82_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08354_ _03342_ _03463_ _03487_ net496 _03485_ vssd1 vssd1 vccd1 vccd1 _03488_ sky130_fd_sc_hd__o221ai_4
XFILLER_0_117_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08426__A net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07305_ top.DUT.register\[15\]\[12\] net679 net675 top.DUT.register\[31\]\[12\] vssd1
+ vssd1 vccd1 vccd1 _02444_ sky130_fd_sc_hd__a22o_1
XFILLER_0_132_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_144_630 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload6 clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 clkload6/Y sky130_fd_sc_hd__inv_6
XANTENNA__10167__S net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08285_ net435 net284 _03420_ vssd1 vssd1 vccd1 vccd1 _03421_ sky130_fd_sc_hd__and3_1
XFILLER_0_132_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10394__C net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09956__S net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07236_ top.DUT.register\[23\]\[10\] net671 net718 top.DUT.register\[19\]\[10\] _02371_
+ vssd1 vssd1 vccd1 vccd1 _02375_ sky130_fd_sc_hd__a221o_1
XFILLER_0_116_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_398 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07167_ _02305_ vssd1 vssd1 vccd1 vccd1 _02306_ sky130_fd_sc_hd__inv_2
XFILLER_0_30_823 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07948__B1 _02111_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07412__A2 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07098_ top.DUT.register\[22\]\[16\] net576 net465 top.DUT.register\[13\]\[16\] vssd1
+ vssd1 vccd1 vccd1 _02237_ sky130_fd_sc_hd__a22o_1
XFILLER_0_112_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06620__B1 net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout210 _04780_ vssd1 vssd1 vccd1 vccd1 net210 sky130_fd_sc_hd__clkbuf_2
Xfanout221 _04766_ vssd1 vssd1 vccd1 vccd1 net221 sky130_fd_sc_hd__clkbuf_2
Xfanout232 _04760_ vssd1 vssd1 vccd1 vccd1 net232 sky130_fd_sc_hd__buf_2
XANTENNA__08960__A2_N net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout243 _04745_ vssd1 vssd1 vccd1 vccd1 net243 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_208_3567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout571_X net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout254 _04741_ vssd1 vssd1 vccd1 vccd1 net254 sky130_fd_sc_hd__buf_1
Xfanout265 _04729_ vssd1 vssd1 vccd1 vccd1 net265 sky130_fd_sc_hd__buf_2
XANTENNA__06887__Y _02026_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout276 net277 vssd1 vssd1 vccd1 vccd1 net276 sky130_fd_sc_hd__buf_2
XANTENNA_fanout669_X net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout287 net294 vssd1 vssd1 vccd1 vccd1 net287 sky130_fd_sc_hd__clkbuf_4
X_09808_ top.pc\[19\] _04471_ vssd1 vssd1 vccd1 vccd1 _04825_ sky130_fd_sc_hd__and2_1
XANTENNA__10630__S net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09704__B _04735_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout298 _02879_ vssd1 vssd1 vccd1 vccd1 net298 sky130_fd_sc_hd__buf_4
XANTENNA__06923__B2 top.DUT.register\[11\]\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09739_ net826 _04328_ _04752_ top.a1.dataIn\[11\] vssd1 vssd1 vccd1 vccd1 _04764_
+ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_2_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_3_4_0_clk_X clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12750_ clknet_leaf_41_clk _00342_ net1056 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[7\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07479__A2 net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11701_ top.a1.dataIn\[10\] _05553_ _05581_ vssd1 vssd1 vccd1 vccd1 _05584_ sky130_fd_sc_hd__and3_1
XANTENNA__06687__B1 net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12681_ clknet_leaf_50_clk _00273_ net1061 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[5\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_166_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11632_ _05488_ _05497_ _05513_ vssd1 vssd1 vccd1 vccd1 _05515_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_108_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06408__X _01547_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_182_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11563_ _05361_ _05419_ vssd1 vssd1 vccd1 vccd1 _05446_ sky130_fd_sc_hd__or2_1
XFILLER_0_9_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10077__S net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13302_ clknet_leaf_4_clk _00894_ net940 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[25\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_123_803 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10514_ net1466 net204 net359 vssd1 vssd1 vccd1 vccd1 _00683_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_447 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13359__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11494_ _05342_ net273 _05343_ vssd1 vssd1 vccd1 vccd1 _05377_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07651__A2 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13233_ clknet_leaf_113_clk _00825_ net990 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[23\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_10445_ net190 top.DUT.register\[16\]\[15\] net367 vssd1 vssd1 vccd1 vccd1 _00616_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_160 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10805__S net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13164_ clknet_leaf_48_clk _00756_ net1060 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[20\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07403__A2 net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08071__A _02069_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10376_ net1382 net199 net375 vssd1 vssd1 vccd1 vccd1 _00551_ sky130_fd_sc_hd__mux2_1
XANTENNA__06611__B1 net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12115_ _05996_ _05997_ vssd1 vssd1 vccd1 vccd1 _05998_ sky130_fd_sc_hd__nand2_1
X_13095_ clknet_leaf_6_clk _00687_ net944 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[18\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_53_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12046_ _05908_ _05916_ _05906_ vssd1 vssd1 vccd1 vccd1 _05929_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_144_2600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_2611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10540__S net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09614__B _04657_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12492__RESET_B net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09313__C1 net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12948_ clknet_leaf_54_clk _00540_ net1075 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[14\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_29_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08667__B2 _03787_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09864__B1 net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09052__D _03711_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06678__B1 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09017__D_N _03708_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12879_ clknet_leaf_32_clk _00471_ net1045 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[11\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_134_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07890__A2 net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_145_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09776__S net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08070_ _02156_ net327 vssd1 vssd1 vccd1 vccd1 _03209_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_155_2773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload101 clknet_leaf_48_clk vssd1 vssd1 vccd1 vccd1 clkload101/Y sky130_fd_sc_hd__inv_6
XANTENNA__07642__A2 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07021_ top.DUT.register\[7\]\[20\] net661 net768 top.DUT.register\[28\]\[20\] _02157_
+ vssd1 vssd1 vccd1 vccd1 _02160_ sky130_fd_sc_hd__a221o_1
XFILLER_0_24_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06850__B1 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10715__S net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_655 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_188_3261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09395__A2 _02025_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_188_3272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08972_ _01741_ net692 net1235 net876 vssd1 vssd1 vccd1 vccd1 _00078_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__06213__B net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07923_ _02571_ _03061_ _03060_ vssd1 vssd1 vccd1 vccd1 _03062_ sky130_fd_sc_hd__a21boi_1
Xhold18 top.ramstore\[18\] vssd1 vssd1 vccd1 vccd1 net1134 sky130_fd_sc_hd__dlygate4sd3_1
Xhold29 top.a1.data\[4\] vssd1 vssd1 vccd1 vccd1 net1145 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08355__B1 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout197_A _04788_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12509__RESET_B net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10450__S net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07854_ _02986_ _02988_ _02990_ _02992_ vssd1 vssd1 vccd1 vccd1 _02993_ sky130_fd_sc_hd__or4_2
X_06805_ top.DUT.register\[1\]\[17\] net755 _01942_ _01943_ vssd1 vssd1 vccd1 vccd1
+ _01944_ sky130_fd_sc_hd__a211o_1
X_07785_ net823 _02904_ _02923_ vssd1 vssd1 vccd1 vccd1 _02924_ sky130_fd_sc_hd__o21ai_1
XANTENNA__06381__A2 net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09524_ _04571_ _04574_ vssd1 vssd1 vccd1 vccd1 _04575_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_203_3486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06736_ _01874_ vssd1 vssd1 vccd1 vccd1 _01875_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_203_3497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09855__B1 net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09455_ top.pc\[22\] _04499_ vssd1 vssd1 vccd1 vccd1 _04510_ sky130_fd_sc_hd__and2_1
X_06667_ top.DUT.register\[22\]\[26\] net577 net445 top.DUT.register\[1\]\[26\] vssd1
+ vssd1 vccd1 vccd1 _01806_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout531_A _01542_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_539 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout629_A _04948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08406_ _03537_ vssd1 vssd1 vccd1 vccd1 _03538_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_164_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09386_ net900 top.pc\[17\] _04445_ net890 vssd1 vssd1 vccd1 vccd1 _00097_ sky130_fd_sc_hd__o211a_1
XANTENNA__08156__A _02723_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06598_ top.DUT.register\[23\]\[28\] net673 net705 top.DUT.register\[3\]\[28\] _01736_
+ vssd1 vssd1 vccd1 vccd1 _01737_ sky130_fd_sc_hd__a221o_1
XFILLER_0_164_736 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07060__A _02198_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08337_ net302 _03346_ vssd1 vssd1 vccd1 vccd1 _03471_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout1061_X net1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07094__B1 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08268_ _03305_ _03309_ net287 vssd1 vssd1 vccd1 vccd1 _03404_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_611 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout998_A net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06841__B1 net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07219_ _02331_ _02356_ vssd1 vssd1 vccd1 vccd1 _02358_ sky130_fd_sc_hd__nor2_1
XANTENNA__10625__S net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08199_ _03042_ net432 net500 _03041_ vssd1 vssd1 vccd1 vccd1 _03337_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_111_2109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_197_Right_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10230_ net144 net1442 net392 vssd1 vssd1 vccd1 vccd1 _00409_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_95_1864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_1875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11193__A2 net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_686 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10161_ net1998 net188 net603 vssd1 vssd1 vccd1 vccd1 _00360_ sky130_fd_sc_hd__mux2_1
Xfanout1005 net1006 vssd1 vssd1 vccd1 vccd1 net1005 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_7_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1016 net1071 vssd1 vssd1 vccd1 vccd1 net1016 sky130_fd_sc_hd__buf_2
Xfanout1027 net1029 vssd1 vssd1 vccd1 vccd1 net1027 sky130_fd_sc_hd__buf_2
XFILLER_0_206_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10092_ net1273 net212 net611 vssd1 vssd1 vccd1 vccd1 _00293_ sky130_fd_sc_hd__mux2_1
Xfanout1038 net1039 vssd1 vssd1 vccd1 vccd1 net1038 sky130_fd_sc_hd__clkbuf_4
Xfanout1049 net1052 vssd1 vssd1 vccd1 vccd1 net1049 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10360__S net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08897__A1 net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_199_655 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12802_ clknet_leaf_10_clk _00394_ net949 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[9\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_187_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13782_ clknet_leaf_69_clk net1119 vssd1 vssd1 vccd1 vccd1 top.pad.button_control.debounce_dly
+ sky130_fd_sc_hd__dfxtp_1
X_10994_ net1151 _05029_ net589 vssd1 vssd1 vccd1 vccd1 _01121_ sky130_fd_sc_hd__mux2_1
XFILLER_0_201_136 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12733_ clknet_leaf_118_clk _00325_ net953 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[7\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_26_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12664_ clknet_leaf_125_clk _00256_ net924 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[5\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_32_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_182_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13720__RESET_B net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11615_ _05497_ vssd1 vssd1 vccd1 vccd1 _05498_ sky130_fd_sc_hd__inv_2
XFILLER_0_182_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12595_ clknet_leaf_122_clk _00187_ net932 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[3\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_65_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07085__B1 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11546_ _05426_ _05427_ vssd1 vssd1 vccd1 vccd1 _05429_ sky130_fd_sc_hd__nor2_1
XFILLER_0_80_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06832__B1 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11477_ _05331_ net273 _05358_ _05359_ vssd1 vssd1 vccd1 vccd1 _05360_ sky130_fd_sc_hd__a31o_1
XFILLER_0_40_428 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10535__S net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13216_ clknet_leaf_80_clk _00808_ net992 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[22\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_10428_ net1411 net143 net370 vssd1 vssd1 vccd1 vccd1 _00600_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_164_Right_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_148_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_150_2692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13147_ clknet_leaf_124_clk _00739_ net925 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[20\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_10359_ net2247 net151 net378 vssd1 vssd1 vccd1 vccd1 _00535_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_209_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13078_ clknet_leaf_3_clk _00670_ net919 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[18\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_183_3191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12029_ _05910_ _05911_ vssd1 vssd1 vccd1 vccd1 _05912_ sky130_fd_sc_hd__nand2_1
XANTENNA__10270__S net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08888__A1 net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06899__B1 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10695__A1 top.a1.instruction\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_205_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07570_ top.DUT.register\[19\]\[6\] net535 net519 top.DUT.register\[10\]\[6\] vssd1
+ vssd1 vccd1 vccd1 _02709_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_66_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06521_ top.DUT.register\[2\]\[29\] net561 net553 top.DUT.register\[3\]\[29\] vssd1
+ vssd1 vccd1 vccd1 _01660_ sky130_fd_sc_hd__a22o_1
XFILLER_0_177_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12197__S _06049_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_157_2802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09240_ net135 _04302_ _04307_ net810 net897 vssd1 vssd1 vccd1 vccd1 _04308_ sky130_fd_sc_hd__o221a_1
X_06452_ top.a1.instruction\[24\] _01590_ vssd1 vssd1 vccd1 vccd1 _01591_ sky130_fd_sc_hd__and2_1
XFILLER_0_29_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07863__A2 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_185_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09171_ _04239_ _04242_ vssd1 vssd1 vccd1 vccd1 _04243_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_146_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06383_ top.a1.instruction\[15\] net782 vssd1 vssd1 vccd1 vccd1 _01522_ sky130_fd_sc_hd__and2_1
X_08122_ net429 net426 _03256_ vssd1 vssd1 vccd1 vccd1 _03261_ sky130_fd_sc_hd__o21a_1
XANTENNA__07076__B1 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_458 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_160_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08053_ _03191_ vssd1 vssd1 vccd1 vccd1 _03192_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10445__S net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07004_ top.DUT.register\[14\]\[20\] net586 net582 top.DUT.register\[30\]\[20\] vssd1
+ vssd1 vccd1 vccd1 _02143_ sky130_fd_sc_hd__a22o_1
XFILLER_0_3_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_131_Right_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_77_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1021_A net1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_168_2964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08955_ net1255 net873 _02304_ net693 vssd1 vssd1 vccd1 vccd1 _00061_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_4_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout481_A _04964_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_208_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_205_3515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout579_A _01514_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_205_3526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07906_ _02996_ _03043_ vssd1 vssd1 vccd1 vccd1 _03045_ sky130_fd_sc_hd__nand2_1
X_08886_ _03956_ _03995_ net287 vssd1 vssd1 vccd1 vccd1 _03996_ sky130_fd_sc_hd__mux2_1
XANTENNA__07000__B1 net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07837_ top.DUT.register\[3\]\[0\] net551 net535 top.DUT.register\[19\]\[0\] vssd1
+ vssd1 vccd1 vccd1 _02976_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_108_2060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout746_A _01622_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_2071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout367_X net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_631 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07768_ top.DUT.register\[21\]\[2\] net655 net750 top.DUT.register\[26\]\[2\] _02906_
+ vssd1 vssd1 vccd1 vccd1 _02907_ sky130_fd_sc_hd__a221o_1
XANTENNA__08438__X _03569_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09507_ net138 _04558_ vssd1 vssd1 vccd1 vccd1 _04559_ sky130_fd_sc_hd__nor2_1
XFILLER_0_94_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06719_ top.DUT.register\[23\]\[25\] net671 net774 top.DUT.register\[13\]\[25\] vssd1
+ vssd1 vccd1 vccd1 _01858_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout534_X net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout913_A net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_2260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07699_ top.DUT.register\[9\]\[4\] net469 net454 top.DUT.register\[29\]\[4\] _02837_
+ vssd1 vssd1 vccd1 vccd1 _02838_ sky130_fd_sc_hd__a221o_1
XFILLER_0_94_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09438_ top.pc\[21\] _04487_ vssd1 vssd1 vccd1 vccd1 _04494_ sky130_fd_sc_hd__xor2_1
XFILLER_0_137_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08945__A1_N _03019_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout701_X net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09369_ top.pc\[17\] _04410_ vssd1 vssd1 vccd1 vccd1 _04429_ sky130_fd_sc_hd__nor2_1
X_11400_ _05246_ _05247_ _05251_ _05218_ top.a1.dataIn\[30\] vssd1 vssd1 vccd1 vccd1
+ _05283_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_97_1904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07067__B1 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07606__A2 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12380_ clknet_leaf_109_clk top.ru.next_FetchedData\[24\] net976 vssd1 vssd1 vccd1
+ vccd1 top.a1.dataIn\[24\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__08614__A net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11331_ top.a1.dataIn\[22\] _05211_ top.a1.dataIn\[23\] vssd1 vssd1 vccd1 vccd1 _05214_
+ sky130_fd_sc_hd__a21o_2
XANTENNA__06814__B1 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10355__S net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11262_ top.a1.row1\[1\] _05124_ _05125_ top.a1.row1\[17\] vssd1 vssd1 vccd1 vccd1
+ _05154_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_37_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_450 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13001_ clknet_leaf_51_clk _00593_ net1035 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[15\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08567__B1 net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10213_ net226 net1768 net394 vssd1 vssd1 vccd1 vccd1 _00393_ sky130_fd_sc_hd__mux2_1
X_11193_ net1264 net587 net473 _05103_ vssd1 vssd1 vccd1 vccd1 _01246_ sky130_fd_sc_hd__a22o_1
XANTENNA__09445__A _02070_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_207_707 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10144_ net142 net1967 net609 vssd1 vssd1 vccd1 vccd1 _00344_ sky130_fd_sc_hd__mux2_1
XFILLER_0_207_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_50_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06593__A2 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10090__S net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10075_ net1994 net157 net618 vssd1 vssd1 vccd1 vccd1 _00277_ sky130_fd_sc_hd__mux2_1
XANTENNA__13547__CLK clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10677__A1 net191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13765_ clknet_leaf_100_clk _01336_ vssd1 vssd1 vccd1 vccd1 top.lcd.cnt_500hz\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__09295__A1 net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10977_ top.a1.dataIn\[3\] net849 _04667_ _05016_ vssd1 vssd1 vccd1 vccd1 _05017_
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_97_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_202_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_703 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12716_ clknet_leaf_65_clk _00308_ net1096 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[6\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13696_ clknet_leaf_89_clk _01267_ vssd1 vssd1 vccd1 vccd1 net112 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_128_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_139_2532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12647_ clknet_leaf_7_clk _00239_ net944 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[4\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_150_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09047__B2 net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_61_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12578_ clknet_leaf_9_clk _00170_ net948 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[2\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_152_2721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_152_2732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11529_ _05396_ _05398_ _05366_ vssd1 vssd1 vccd1 vccd1 _05412_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_13_428 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10265__S net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwire271 net272 vssd1 vssd1 vccd1 vccd1 net271 sky130_fd_sc_hd__clkbuf_1
Xhold307 top.DUT.register\[17\]\[28\] vssd1 vssd1 vccd1 vccd1 net1423 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_151_772 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold318 top.DUT.register\[8\]\[18\] vssd1 vssd1 vccd1 vccd1 net1434 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold329 top.a1.row2\[17\] vssd1 vssd1 vccd1 vccd1 net1445 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_185_3220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_647 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08022__A2 _03142_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout809 _01574_ vssd1 vssd1 vccd1 vccd1 net809 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_0_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07230__B1 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06584__A2 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08740_ net289 _03206_ _03210_ vssd1 vssd1 vccd1 vccd1 _03857_ sky130_fd_sc_hd__and3_1
Xhold1007 top.DUT.register\[30\]\[13\] vssd1 vssd1 vccd1 vccd1 net2123 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1018 top.DUT.register\[9\]\[24\] vssd1 vssd1 vccd1 vccd1 net2134 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1029 top.DUT.register\[23\]\[2\] vssd1 vssd1 vccd1 vccd1 net2145 sky130_fd_sc_hd__dlygate4sd3_1
X_08671_ net322 _03409_ _03535_ vssd1 vssd1 vccd1 vccd1 _03791_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11109__B net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_163_2894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07622_ top.DUT.register\[23\]\[5\] net571 net535 top.DUT.register\[19\]\[5\] vssd1
+ vssd1 vccd1 vccd1 _02761_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_200_3445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07553_ top.DUT.register\[7\]\[7\] net659 net714 top.DUT.register\[27\]\[7\] _02688_
+ vssd1 vssd1 vccd1 vccd1 _02692_ sky130_fd_sc_hd__a221o_1
XFILLER_0_76_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_193_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_196_3382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06504_ net788 _01596_ _01607_ vssd1 vssd1 vccd1 vccd1 _01643_ sky130_fd_sc_hd__and3_4
XFILLER_0_76_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_196_3393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07297__B1 net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07484_ _02616_ _02618_ _02620_ _02622_ vssd1 vssd1 vccd1 vccd1 _02623_ sky130_fd_sc_hd__or4_4
XFILLER_0_146_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_200_Right_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09223_ _02497_ _02502_ vssd1 vssd1 vccd1 vccd1 _04292_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_185_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06435_ _01573_ _01473_ vssd1 vssd1 vccd1 vccd1 _01574_ sky130_fd_sc_hd__and2b_1
XFILLER_0_90_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_173_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1069_A net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09089__X _04164_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09154_ top.pc\[4\] _02857_ vssd1 vssd1 vccd1 vccd1 _04227_ sky130_fd_sc_hd__or2_1
X_06366_ top.a1.instruction\[3\] net829 vssd1 vssd1 vccd1 vccd1 _01505_ sky130_fd_sc_hd__nor2_4
XTAP_TAPCELL_ROW_79_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08105_ _02409_ net327 vssd1 vssd1 vccd1 vccd1 _03244_ sky130_fd_sc_hd__nand2_1
XFILLER_0_161_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_575 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10175__S net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09085_ _04157_ _04158_ _04159_ vssd1 vssd1 vccd1 vccd1 _04160_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_15_Left_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06297_ _01453_ _01454_ _01452_ vssd1 vssd1 vccd1 vccd1 _01455_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09964__S net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08036_ net304 _03173_ vssd1 vssd1 vccd1 vccd1 _03175_ sky130_fd_sc_hd__or2_1
XFILLER_0_114_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold830 top.DUT.register\[7\]\[11\] vssd1 vssd1 vccd1 vccd1 net1946 sky130_fd_sc_hd__dlygate4sd3_1
Xhold841 top.DUT.register\[29\]\[9\] vssd1 vssd1 vccd1 vccd1 net1957 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout696_A net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold852 top.DUT.register\[22\]\[23\] vssd1 vssd1 vccd1 vccd1 net1968 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold863 top.a1.row1\[15\] vssd1 vssd1 vccd1 vccd1 net1979 sky130_fd_sc_hd__dlygate4sd3_1
Xhold874 top.DUT.register\[3\]\[11\] vssd1 vssd1 vccd1 vccd1 net1990 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10903__S net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold885 top.DUT.register\[1\]\[8\] vssd1 vssd1 vccd1 vccd1 net2001 sky130_fd_sc_hd__dlygate4sd3_1
Xhold896 top.DUT.register\[18\]\[21\] vssd1 vssd1 vccd1 vccd1 net2012 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09761__A2 _04370_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09987_ net247 net1886 net623 vssd1 vssd1 vccd1 vccd1 _00192_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout863_A _01428_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout484_X net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06575__A2 net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08938_ _04028_ _04045_ vssd1 vssd1 vccd1 vccd1 _04046_ sky130_fd_sc_hd__nand2_1
XANTENNA__10108__A0 top.DUT.register\[6\]\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12399__Q top.a1.instruction\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08869_ net317 _03654_ _03587_ vssd1 vssd1 vccd1 vccd1 _03980_ sky130_fd_sc_hd__o21ai_2
XANTENNA_fanout651_X net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_24_Left_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11320__A2 _04658_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout749_X net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10900_ net1608 net212 net478 vssd1 vssd1 vccd1 vccd1 _01061_ sky130_fd_sc_hd__mux2_1
XFILLER_0_169_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11880_ _05735_ _05751_ vssd1 vssd1 vccd1 vccd1 _05763_ sky130_fd_sc_hd__nor2_1
XFILLER_0_168_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_196_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10831_ net1651 net247 net474 vssd1 vssd1 vccd1 vccd1 _00992_ sky130_fd_sc_hd__mux2_1
XANTENNA__09277__A1 net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_196_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13550_ clknet_leaf_104_clk _01137_ net972 vssd1 vssd1 vccd1 vccd1 top.ramload\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11084__A1 net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10762_ net2285 net265 net482 vssd1 vssd1 vccd1 vccd1 _00923_ sky130_fd_sc_hd__mux2_1
XFILLER_0_183_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_36_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_11_Right_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07827__A2 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12501_ clknet_leaf_111_clk _00093_ net990 vssd1 vssd1 vccd1 vccd1 top.pc\[13\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_54_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13481_ clknet_leaf_52_clk _01073_ net1039 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[30\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_101_1963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10693_ net1419 net142 net340 vssd1 vssd1 vccd1 vccd1 _00856_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_192_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12432_ clknet_leaf_93_clk _00028_ net998 vssd1 vssd1 vccd1 vccd1 top.ramaddr\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07659__S net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_33_Left_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_43_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08788__B1 net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12363_ clknet_leaf_103_clk top.ru.next_FetchedData\[7\] net980 vssd1 vssd1 vccd1
+ vccd1 top.a1.dataIn\[7\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_62_372 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10085__S net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08252__A2 _03370_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_134_2451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_2462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11314_ top.a1.row1\[111\] _05178_ _05190_ _05199_ vssd1 vssd1 vccd1 vccd1 _05200_
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_133_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07460__B1 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12294_ _01404_ _06106_ _06107_ net686 vssd1 vssd1 vccd1 vccd1 _01349_ sky130_fd_sc_hd__o211a_1
X_11245_ top.a1.row1\[0\] _05124_ _05127_ _05137_ vssd1 vssd1 vccd1 vccd1 _05138_
+ sky130_fd_sc_hd__a211o_1
XANTENNA__10813__S net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_20_Right_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09175__A _02773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11176_ _05004_ _05018_ _05098_ net588 net1161 vssd1 vssd1 vccd1 vccd1 _01234_ sky130_fd_sc_hd__a32o_1
XANTENNA__06566__A2 net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10127_ net198 net2179 net609 vssd1 vssd1 vccd1 vccd1 _00327_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_42_Left_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_180_3150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10058_ net2126 net219 net615 vssd1 vssd1 vccd1 vccd1 _00260_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_199_260 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13817_ net1102 vssd1 vssd1 vccd1 vccd1 gpio_out[4] sky130_fd_sc_hd__buf_2
XFILLER_0_161_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07279__B1 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_34_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13748_ clknet_leaf_99_clk _01319_ vssd1 vssd1 vccd1 vccd1 top.lcd.cnt_20ms\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_678 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07818__A2 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_51_Left_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_14_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13679_ clknet_leaf_91_clk _01255_ net997 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_06220_ top.ramload\[14\] net856 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedInstr\[14\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_183_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_372 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06151_ top.edg2.flip2 vssd1 vssd1 vccd1 vccd1 _01394_ sky130_fd_sc_hd__inv_2
XFILLER_0_130_208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold104 top.DUT.register\[4\]\[7\] vssd1 vssd1 vccd1 vccd1 net1220 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold115 top.pad.button_control.r_counter\[12\] vssd1 vssd1 vccd1 vccd1 net1231 sky130_fd_sc_hd__dlygate4sd3_1
Xhold126 net73 vssd1 vssd1 vccd1 vccd1 net1242 sky130_fd_sc_hd__dlygate4sd3_1
Xhold137 top.DUT.register\[23\]\[20\] vssd1 vssd1 vccd1 vccd1 net1253 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold148 top.a1.row1\[123\] vssd1 vssd1 vccd1 vccd1 net1264 sky130_fd_sc_hd__dlygate4sd3_1
Xhold159 top.DUT.register\[3\]\[19\] vssd1 vssd1 vccd1 vccd1 net1275 sky130_fd_sc_hd__dlygate4sd3_1
X_09910_ _04008_ net407 vssd1 vssd1 vccd1 vccd1 _04917_ sky130_fd_sc_hd__nand2_1
XANTENNA__10723__S net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09841_ _04514_ net486 net401 top.a1.dataIn\[22\] net397 vssd1 vssd1 vccd1 vccd1
+ _04855_ sky130_fd_sc_hd__a221o_1
Xfanout617 _04954_ vssd1 vssd1 vccd1 vccd1 net617 sky130_fd_sc_hd__buf_6
XPHY_EDGE_ROW_60_Left_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout628 _04948_ vssd1 vssd1 vccd1 vccd1 net628 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06557__A2 net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_165_2923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout639 _01619_ vssd1 vssd1 vccd1 vccd1 net639 sky130_fd_sc_hd__clkbuf_8
XANTENNA__08951__B1 _02701_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09772_ _04789_ _04790_ vssd1 vssd1 vccd1 vccd1 _04793_ sky130_fd_sc_hd__xnor2_1
X_06984_ top.DUT.register\[9\]\[23\] net763 net713 top.DUT.register\[11\]\[23\] vssd1
+ vssd1 vccd1 vccd1 _02123_ sky130_fd_sc_hd__a22o_1
XANTENNA__06221__B net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08723_ _02091_ net493 _03185_ vssd1 vssd1 vccd1 vccd1 _03841_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_198_3411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_198_3422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08654_ _03687_ _03774_ net308 vssd1 vssd1 vccd1 vccd1 _03775_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07605_ top.DUT.register\[24\]\[6\] net643 net726 top.DUT.register\[18\]\[6\] _02743_
+ vssd1 vssd1 vccd1 vccd1 _02744_ sky130_fd_sc_hd__a221o_1
X_08585_ net286 _03524_ _03527_ net275 vssd1 vssd1 vccd1 vccd1 _03709_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout444_A _01564_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_431 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07536_ top.DUT.register\[8\]\[7\] net539 net519 top.DUT.register\[10\]\[7\] vssd1
+ vssd1 vccd1 vccd1 _02675_ sky130_fd_sc_hd__a22o_1
XFILLER_0_48_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09959__S net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_522 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_544 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07467_ top.DUT.register\[25\]\[15\] net779 net765 top.DUT.register\[9\]\[15\] vssd1
+ vssd1 vccd1 vccd1 _02606_ sky130_fd_sc_hd__a22o_1
XANTENNA__10694__A top.a1.instruction\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout611_A net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout709_A _01640_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09206_ _02678_ _02682_ vssd1 vssd1 vccd1 vccd1 _04276_ sky130_fd_sc_hd__nand2_1
X_06418_ top.DUT.register\[17\]\[30\] net461 net457 top.DUT.register\[25\]\[30\] _01556_
+ vssd1 vssd1 vccd1 vccd1 _01557_ sky130_fd_sc_hd__a221o_1
XFILLER_0_134_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07398_ top.DUT.register\[23\]\[9\] net571 net539 top.DUT.register\[8\]\[9\] _02536_
+ vssd1 vssd1 vccd1 vccd1 _02537_ sky130_fd_sc_hd__a221o_1
XFILLER_0_161_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09137_ top.pc\[1\] _02952_ _04187_ _04185_ vssd1 vssd1 vccd1 vccd1 _04211_ sky130_fd_sc_hd__a31oi_1
X_06349_ top.d_ready _01479_ _01485_ _01488_ top.ru.next_read_i vssd1 vssd1 vccd1
+ vccd1 _00007_ sky130_fd_sc_hd__o41a_1
XFILLER_0_44_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09068_ _01391_ top.a1.instruction\[13\] _02343_ vssd1 vssd1 vccd1 vccd1 _04143_
+ sky130_fd_sc_hd__o21a_1
XANTENNA__07442__B1 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout980_A net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_2181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_2192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06796__A2 net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout699_X net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08019_ _01589_ _03157_ vssd1 vssd1 vccd1 vccd1 _03158_ sky130_fd_sc_hd__nor2_1
XANTENNA__10633__S net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold660 top.DUT.register\[22\]\[8\] vssd1 vssd1 vccd1 vccd1 net1776 sky130_fd_sc_hd__dlygate4sd3_1
Xhold671 top.DUT.register\[4\]\[25\] vssd1 vssd1 vccd1 vccd1 net1787 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11030_ net9 net839 net817 net1178 vssd1 vssd1 vccd1 vccd1 _01142_ sky130_fd_sc_hd__o22a_1
Xhold682 top.DUT.register\[15\]\[1\] vssd1 vssd1 vccd1 vccd1 net1798 sky130_fd_sc_hd__dlygate4sd3_1
Xhold693 top.DUT.register\[3\]\[24\] vssd1 vssd1 vccd1 vccd1 net1809 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06548__A2 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout866_X net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09723__A _04172_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12981_ clknet_leaf_32_clk _00573_ net1023 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[15\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09498__B2 top.pc\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11932_ _05805_ _05809_ _05813_ _05814_ vssd1 vssd1 vccd1 vccd1 _05815_ sky130_fd_sc_hd__nor4_1
XFILLER_0_87_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_197_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11863_ _05679_ _05745_ vssd1 vssd1 vccd1 vccd1 _05746_ sky130_fd_sc_hd__and2_1
XANTENNA__06720__A2 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13602_ clknet_leaf_64_clk net1148 net1093 vssd1 vssd1 vccd1 vccd1 net94 sky130_fd_sc_hd__dfrtp_1
X_10814_ net182 net1877 net599 vssd1 vssd1 vccd1 vccd1 _00975_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_45_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11794_ _05648_ _05676_ vssd1 vssd1 vccd1 vccd1 _05677_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_156_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13533_ clknet_leaf_93_clk _01120_ net995 vssd1 vssd1 vccd1 vccd1 top.a1.data\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_10745_ net1449 net217 net419 vssd1 vssd1 vccd1 vccd1 _00906_ sky130_fd_sc_hd__mux2_1
XANTENNA__09670__A1 net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10808__S net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_11_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07681__B1 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13464_ clknet_leaf_128_clk _01056_ net913 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[30\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10676_ net1470 net196 net340 vssd1 vssd1 vccd1 vccd1 _00839_ sky130_fd_sc_hd__mux2_1
XANTENNA__13688__Q top.lcd.nextState\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12415_ clknet_leaf_109_clk top.ru.next_FetchedInstr\[27\] net977 vssd1 vssd1 vccd1
+ vccd1 top.a1.instruction\[27\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_106_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13395_ clknet_leaf_121_clk _00987_ net932 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[28\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_152_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12346_ net2278 net904 net37 vssd1 vssd1 vccd1 vccd1 _01371_ sky130_fd_sc_hd__a21o_1
XFILLER_0_11_707 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07433__B1 net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06787__A2 net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12277_ top.lcd.cnt_500hz\[7\] top.lcd.cnt_500hz\[8\] _06094_ vssd1 vssd1 vccd1 vccd1
+ _06097_ sky130_fd_sc_hd__and3_1
XANTENNA__10543__S net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11228_ top.a1.row2\[12\] _05119_ _05120_ _01442_ vssd1 vssd1 vccd1 vccd1 _05121_
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_208_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_207_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11159_ top.a1.hexop\[4\] _01417_ _01414_ net888 vssd1 vssd1 vccd1 vccd1 _05088_
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_65_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_147_2653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_160_2842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_160_2853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire412_A _02260_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09920__X _04927_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_203_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06711__A2 net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08370_ _03450_ _03502_ net292 vssd1 vssd1 vccd1 vccd1 _03503_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_193_3341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08536__X _03663_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_175_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07321_ top.DUT.register\[26\]\[12\] net750 net746 top.DUT.register\[17\]\[12\] vssd1
+ vssd1 vccd1 vccd1 _02460_ sky130_fd_sc_hd__a22o_1
XFILLER_0_190_406 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10718__S net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_156_683 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_300 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07252_ top.DUT.register\[19\]\[13\] net538 net528 top.DUT.register\[26\]\[13\] vssd1
+ vssd1 vccd1 vccd1 _02391_ sky130_fd_sc_hd__a22o_1
XFILLER_0_155_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07672__B1 net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06203_ _01386_ wb.curr_state\[0\] top.Ren wb.curr_state\[1\] net905 vssd1 vssd1
+ vccd1 vccd1 _00014_ sky130_fd_sc_hd__a32o_1
XFILLER_0_26_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07183_ top.DUT.register\[6\]\[10\] net567 net463 top.DUT.register\[13\]\[10\] vssd1
+ vssd1 vccd1 vccd1 _02322_ sky130_fd_sc_hd__a22o_1
XANTENNA__08216__A2 top.pc\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06216__B net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_170_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07424__B1 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10961__B net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06778__A2 _01916_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10453__S net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09527__B _04577_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09177__B1 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout403 net406 vssd1 vssd1 vccd1 vccd1 net403 sky130_fd_sc_hd__buf_4
XANTENNA__06232__A top.ramload\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout425 _03341_ vssd1 vssd1 vccd1 vccd1 net425 sky130_fd_sc_hd__clkbuf_2
Xfanout436 _03168_ vssd1 vssd1 vccd1 vccd1 net436 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout394_A net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout447 _01562_ vssd1 vssd1 vccd1 vccd1 net447 sky130_fd_sc_hd__buf_4
X_09824_ net798 _04837_ _04838_ _04839_ vssd1 vssd1 vccd1 vccd1 _04840_ sky130_fd_sc_hd__a211o_1
Xfanout458 _01553_ vssd1 vssd1 vccd1 vccd1 net458 sky130_fd_sc_hd__buf_4
Xfanout469 net470 vssd1 vssd1 vccd1 vccd1 net469 sky130_fd_sc_hd__buf_4
X_09755_ _04774_ _04775_ _04777_ vssd1 vssd1 vccd1 vccd1 _04778_ sky130_fd_sc_hd__o21ai_1
X_06967_ top.DUT.register\[8\]\[23\] net540 net512 top.DUT.register\[24\]\[23\] vssd1
+ vssd1 vccd1 vccd1 _02106_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout561_A _01532_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06950__A2 net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout659_A net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08706_ _02179_ net492 net433 _02178_ vssd1 vssd1 vccd1 vccd1 _03825_ sky130_fd_sc_hd__a2bb2o_1
X_09686_ _04173_ _04715_ vssd1 vssd1 vccd1 vccd1 _04722_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_87_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06898_ top.DUT.register\[20\]\[18\] net665 net735 top.DUT.register\[16\]\[18\] vssd1
+ vssd1 vccd1 vccd1 _02037_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_87_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08637_ _03754_ _03758_ vssd1 vssd1 vccd1 vccd1 _03759_ sky130_fd_sc_hd__nor2_1
XFILLER_0_179_764 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout447_X net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout826_A net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06702__A2 net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09689__S net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08593__S net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08568_ _02656_ net494 _03691_ net436 _03692_ vssd1 vssd1 vccd1 vccd1 _03693_ sky130_fd_sc_hd__a221o_1
X_07519_ _02525_ _02571_ _02657_ vssd1 vssd1 vccd1 vccd1 _02658_ sky130_fd_sc_hd__and3_1
XFILLER_0_92_732 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08499_ _03277_ _03281_ vssd1 vssd1 vccd1 vccd1 _03627_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout614_X net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10530_ net1409 net144 _04988_ vssd1 vssd1 vccd1 vccd1 _00697_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_118_2210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_118_2221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06407__A top.a1.instruction\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_40_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10461_ net140 net2054 net367 vssd1 vssd1 vccd1 vccd1 _00632_ sky130_fd_sc_hd__mux2_1
X_12200_ net1156 _06005_ _06049_ vssd1 vssd1 vccd1 vccd1 _01307_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13180_ clknet_leaf_0_clk _00772_ net915 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[21\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_3_0_0_clk_X clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07415__B1 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_2410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_731 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10392_ net1917 net149 net375 vssd1 vssd1 vccd1 vccd1 _00567_ sky130_fd_sc_hd__mux2_1
XANTENNA__08622__A _03744_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06769__A2 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12131_ _06012_ _06013_ vssd1 vssd1 vccd1 vccd1 _06014_ sky130_fd_sc_hd__nand2_1
XANTENNA__10363__S net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_208_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12062_ _05935_ _05937_ _05944_ vssd1 vssd1 vccd1 vccd1 _05945_ sky130_fd_sc_hd__a21oi_1
XANTENNA__06142__A net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold490 top.DUT.register\[14\]\[3\] vssd1 vssd1 vccd1 vccd1 net1606 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07718__A1 top.a1.instruction\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11013_ net887 net842 wb.prev_BUSY_O vssd1 vssd1 vccd1 vccd1 _05044_ sky130_fd_sc_hd__or3b_4
Xfanout970 net971 vssd1 vssd1 vccd1 vccd1 net970 sky130_fd_sc_hd__clkbuf_2
Xfanout981 net987 vssd1 vssd1 vccd1 vccd1 net981 sky130_fd_sc_hd__clkbuf_4
Xfanout992 net993 vssd1 vssd1 vccd1 vccd1 net992 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_129_2383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06941__A2 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12964_ clknet_leaf_37_clk _00556_ net1051 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[14\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_99_375 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1190 top.lcd.currentState\[2\] vssd1 vssd1 vccd1 vccd1 net2306 sky130_fd_sc_hd__dlygate4sd3_1
X_11915_ _05795_ _05797_ vssd1 vssd1 vccd1 vccd1 _05798_ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_142_2572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_142_2583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_263 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12895_ clknet_leaf_19_clk _00487_ net1026 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[12\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09900__B _04605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11846_ _05727_ _05728_ vssd1 vssd1 vccd1 vccd1 _05729_ sky130_fd_sc_hd__or2_1
XFILLER_0_51_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07260__X _02399_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_200_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_175_3071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11777_ top.a1.dataIn\[8\] _05585_ _05625_ vssd1 vssd1 vccd1 vccd1 _05660_ sky130_fd_sc_hd__or3_1
XANTENNA__10538__S net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_672 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13516_ clknet_leaf_64_clk _01108_ net1092 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[31\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07654__B1 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10728_ net2200 net146 net421 vssd1 vssd1 vccd1 vccd1 _00889_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13447_ clknet_leaf_6_clk _01039_ net937 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[29\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_10659_ net149 net1838 net344 vssd1 vssd1 vccd1 vccd1 _00823_ sky130_fd_sc_hd__mux2_1
Xclkload13 clknet_leaf_130_clk vssd1 vssd1 vccd1 vccd1 clkload13/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload24 clknet_leaf_12_clk vssd1 vssd1 vccd1 vccd1 clkload24/Y sky130_fd_sc_hd__inv_6
Xclkload35 clknet_leaf_108_clk vssd1 vssd1 vccd1 vccd1 clkload35/Y sky130_fd_sc_hd__clkinv_8
XTAP_TAPCELL_ROW_58_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload46 clknet_leaf_81_clk vssd1 vssd1 vccd1 vccd1 clkload46/Y sky130_fd_sc_hd__inv_8
XFILLER_0_140_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08091__X _03230_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13378_ clknet_leaf_9_clk _00970_ net949 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[27\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload57 clknet_leaf_93_clk vssd1 vssd1 vccd1 vccd1 clkload57/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_23_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload68 clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 clkload68/Y sky130_fd_sc_hd__clkinv_4
Xclkload79 clknet_leaf_40_clk vssd1 vssd1 vccd1 vccd1 clkload79/Y sky130_fd_sc_hd__clkinvlp_4
X_12329_ net1672 _06127_ _06129_ vssd1 vssd1 vccd1 vccd1 _01362_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10273__S net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07870_ top.DUT.register\[13\]\[1\] net775 net713 top.DUT.register\[11\]\[1\] _03002_
+ vssd1 vssd1 vccd1 vccd1 _03009_ sky130_fd_sc_hd__a221o_1
XANTENNA__07185__A2 net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08382__A1 net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08382__B2 _03514_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06821_ _01950_ _01959_ vssd1 vssd1 vccd1 vccd1 _01960_ sky130_fd_sc_hd__nor2_4
XFILLER_0_208_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06932__A2 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09540_ top.a1.instruction\[27\] net821 net422 vssd1 vssd1 vccd1 vccd1 _04590_ sky130_fd_sc_hd__a21o_2
X_06752_ top.DUT.register\[13\]\[24\] net466 net562 top.DUT.register\[2\]\[24\] _01890_
+ vssd1 vssd1 vccd1 vccd1 _01891_ sky130_fd_sc_hd__a221o_1
XANTENNA__09082__B top.a1.instruction\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_183_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_183_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12655__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_wire415_X net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11117__B net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09471_ _04509_ _04510_ _04511_ vssd1 vssd1 vccd1 vccd1 _04525_ sky130_fd_sc_hd__o21a_1
X_06683_ top.DUT.register\[23\]\[26\] net673 net712 top.DUT.register\[11\]\[26\] _01811_
+ vssd1 vssd1 vccd1 vccd1 _01822_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_69_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_370 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_69_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08422_ _03502_ _03552_ net292 vssd1 vssd1 vccd1 vccd1 _03553_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10956__B _04998_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07611__A _02723_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08353_ _02803_ _03486_ vssd1 vssd1 vccd1 vccd1 _03487_ sky130_fd_sc_hd__xor2_2
XANTENNA__10448__S net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_82_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08426__B _03556_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07304_ _02436_ _02438_ _02440_ _02442_ vssd1 vssd1 vccd1 vccd1 _02443_ sky130_fd_sc_hd__or4_4
XPHY_EDGE_ROW_178_Right_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_190_236 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08284_ net307 _03419_ vssd1 vssd1 vccd1 vccd1 _03420_ sky130_fd_sc_hd__nor2_1
XANTENNA__07645__B1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload7 clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 clkload7/Y sky130_fd_sc_hd__clkinv_4
XANTENNA__06227__A top.ramload\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06999__A2 net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07235_ top.DUT.register\[14\]\[10\] net730 net698 top.DUT.register\[31\]\[10\] _02372_
+ vssd1 vssd1 vccd1 vccd1 _02374_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout407_A _04716_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09097__X _04172_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07166_ net823 _02304_ _01586_ vssd1 vssd1 vccd1 vccd1 _02305_ sky130_fd_sc_hd__a21o_1
XFILLER_0_30_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_113_2140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07097_ top.DUT.register\[25\]\[16\] net456 net512 top.DUT.register\[24\]\[16\] _02235_
+ vssd1 vssd1 vccd1 vccd1 _02236_ sky130_fd_sc_hd__a221o_1
XFILLER_0_100_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09972__S net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09825__X _04841_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout200 net201 vssd1 vssd1 vccd1 vccd1 net200 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout776_A net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout211 net214 vssd1 vssd1 vccd1 vccd1 net211 sky130_fd_sc_hd__buf_2
Xfanout222 _04766_ vssd1 vssd1 vccd1 vccd1 net222 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_10_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout233 _04760_ vssd1 vssd1 vccd1 vccd1 net233 sky130_fd_sc_hd__clkbuf_2
Xfanout244 _04745_ vssd1 vssd1 vccd1 vccd1 net244 sky130_fd_sc_hd__buf_1
XANTENNA__10911__S net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout255 _04737_ vssd1 vssd1 vccd1 vccd1 net255 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_208_3568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07176__A2 net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout266 _04729_ vssd1 vssd1 vccd1 vccd1 net266 sky130_fd_sc_hd__buf_1
XANTENNA__09273__A _02286_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout277 _03021_ vssd1 vssd1 vccd1 vccd1 net277 sky130_fd_sc_hd__clkbuf_4
X_09807_ _04819_ _04820_ _04817_ vssd1 vssd1 vccd1 vccd1 _04824_ sky130_fd_sc_hd__o21ai_1
Xfanout288 net294 vssd1 vssd1 vccd1 vccd1 net288 sky130_fd_sc_hd__clkbuf_2
Xfanout299 net300 vssd1 vssd1 vccd1 vccd1 net299 sky130_fd_sc_hd__buf_2
XANTENNA_fanout943_A net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout564_X net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07999_ top.DUT.register\[9\]\[31\] net763 net736 top.DUT.register\[16\]\[31\] vssd1
+ vssd1 vccd1 vccd1 _03138_ sky130_fd_sc_hd__a22o_1
XANTENNA__06923__A2 net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09738_ net2139 net228 net631 vssd1 vssd1 vccd1 vccd1 _00131_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_2_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout731_X net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09669_ _04184_ _04703_ _04705_ _01505_ vssd1 vssd1 vccd1 vccd1 _04706_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout829_X net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11700_ _05553_ _05581_ top.a1.dataIn\[10\] vssd1 vssd1 vccd1 vccd1 _05583_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_167_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12680_ clknet_leaf_26_clk _00272_ net1011 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[5\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07884__B1 net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_194_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_166_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11631_ _05489_ _05497_ _05507_ _05510_ vssd1 vssd1 vccd1 vccd1 _05514_ sky130_fd_sc_hd__or4bb_2
XFILLER_0_194_575 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10358__S net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_194_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13829__1113 vssd1 vssd1 vccd1 vccd1 _13829__1113/HI net1113 sky130_fd_sc_hd__conb_1
X_11562_ net249 _05420_ vssd1 vssd1 vccd1 vccd1 _05445_ sky130_fd_sc_hd__and2b_1
XPHY_EDGE_ROW_7_Left_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_145_Right_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07100__A2 net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10513_ net1326 net215 net360 vssd1 vssd1 vccd1 vccd1 _00682_ sky130_fd_sc_hd__mux2_1
X_13301_ clknet_leaf_31_clk _00893_ net1018 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[25\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_123_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_21_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11493_ _05338_ _05367_ vssd1 vssd1 vccd1 vccd1 _05376_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_52_459 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_612 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_hold988_A top.ramload\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13232_ clknet_leaf_26_clk _00824_ net1011 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[22\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_10444_ net196 net1952 net367 vssd1 vssd1 vccd1 vccd1 _00615_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07939__A1 _02049_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12870__Q top.DUT.register\[11\]\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_172 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13163_ clknet_leaf_48_clk _00755_ net1060 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[20\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10093__S net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10375_ net1221 net209 net375 vssd1 vssd1 vccd1 vccd1 _00550_ sky130_fd_sc_hd__mux2_1
X_12114_ _05986_ _05992_ _05991_ vssd1 vssd1 vccd1 vccd1 _05997_ sky130_fd_sc_hd__a21o_1
X_13094_ clknet_leaf_40_clk _00686_ net1053 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[18\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_12045_ _05922_ _05924_ vssd1 vssd1 vccd1 vccd1 _05928_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_53_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10821__S net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09561__B1 _01505_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_144_2601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_2612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06914__A2 net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_177_3100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12947_ clknet_leaf_124_clk _00539_ net926 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[14\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09864__A1 _03909_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_197_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07875__B1 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12878_ clknet_leaf_39_clk _00470_ net1054 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[11\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_185_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_190_3300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11829_ _05678_ _05682_ net131 vssd1 vssd1 vccd1 vccd1 _05712_ sky130_fd_sc_hd__o21a_1
XANTENNA__10268__S net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10495__C net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07627__B1 net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_112_Right_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13303__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_155_2774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload102 clknet_leaf_49_clk vssd1 vssd1 vccd1 vccd1 clkload102/Y sky130_fd_sc_hd__inv_6
XFILLER_0_102_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07020_ top.DUT.register\[24\]\[20\] net646 net642 top.DUT.register\[8\]\[20\] _02158_
+ vssd1 vssd1 vccd1 vccd1 _02159_ sky130_fd_sc_hd__a221o_1
XFILLER_0_153_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_49_Right_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_141_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_188_3262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_188_3273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08971_ _01783_ net692 net1197 net875 vssd1 vssd1 vccd1 vccd1 _00077_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__12517__SET_B net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10731__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07922_ _02498_ _02522_ vssd1 vssd1 vccd1 vccd1 _03061_ sky130_fd_sc_hd__and2_1
Xhold19 _01178_ vssd1 vssd1 vccd1 vccd1 net1135 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07158__A2 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08355__A1 net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07165__X _02304_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08355__B2 _03488_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07853_ top.DUT.register\[13\]\[0\] net466 net452 top.DUT.register\[29\]\[0\] _02991_
+ vssd1 vssd1 vccd1 vccd1 _02992_ sky130_fd_sc_hd__a221o_1
XANTENNA__06905__A2 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06804_ top.DUT.register\[2\]\[17\] net743 net703 top.DUT.register\[3\]\[17\] vssd1
+ vssd1 vccd1 vccd1 _01943_ sky130_fd_sc_hd__a22o_1
X_07784_ net809 _02922_ vssd1 vssd1 vccd1 vccd1 _02923_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_58_Right_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06735_ _01853_ _01873_ vssd1 vssd1 vccd1 vccd1 _01874_ sky130_fd_sc_hd__and2_1
XFILLER_0_78_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_84_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09523_ _04572_ _04573_ vssd1 vssd1 vccd1 vccd1 _04574_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_203_3487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10967__A top.a1.halfData\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09855__A1 _03890_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_203_3498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout357_A net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09454_ top.pc\[21\] _04487_ _04496_ vssd1 vssd1 vccd1 vccd1 _04509_ sky130_fd_sc_hd__a21o_1
X_06666_ top.DUT.register\[25\]\[26\] net457 net505 top.DUT.register\[27\]\[26\] _01804_
+ vssd1 vssd1 vccd1 vccd1 _01805_ sky130_fd_sc_hd__a221o_1
XANTENNA__07866__B1 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_391 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07330__A2 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08405_ _03533_ _03535_ vssd1 vssd1 vccd1 vccd1 _03537_ sky130_fd_sc_hd__nor2_1
XFILLER_0_93_348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09385_ net137 _04430_ _04444_ vssd1 vssd1 vccd1 vccd1 _04445_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_136_406 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06597_ top.DUT.register\[20\]\[28\] net666 net650 top.DUT.register\[22\]\[28\] vssd1
+ vssd1 vccd1 vccd1 _01736_ sky130_fd_sc_hd__a22o_1
XFILLER_0_176_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout524_A _01554_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_176_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08336_ net302 _03346_ vssd1 vssd1 vccd1 vccd1 _03470_ sky130_fd_sc_hd__nor2_1
XFILLER_0_164_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11414__A1 top.a1.dataIn\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07618__B1 net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09967__S net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_236 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08267_ _03319_ _03302_ net288 vssd1 vssd1 vccd1 vccd1 _03403_ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10906__S net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_67_Right_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_623 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07218_ _02356_ vssd1 vssd1 vccd1 vccd1 _02357_ sky130_fd_sc_hd__inv_2
XFILLER_0_116_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08172__A _01940_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08198_ _03043_ _03179_ vssd1 vssd1 vccd1 vccd1 _03336_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_15_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11178__B1 net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07149_ top.DUT.register\[5\]\[11\] net651 net770 top.DUT.register\[10\]\[11\] vssd1
+ vssd1 vccd1 vccd1 _02288_ sky130_fd_sc_hd__a22o_1
XANTENNA__07059__Y _02198_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_1865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09240__C1 net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_1876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07397__A2 net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10160_ net1954 net199 net604 vssd1 vssd1 vccd1 vccd1 _00359_ sky130_fd_sc_hd__mux2_1
XFILLER_0_112_391 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout681_X net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout779_X net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1006 net1007 vssd1 vssd1 vccd1 vccd1 net1006 sky130_fd_sc_hd__clkbuf_4
X_10091_ net1498 net219 net612 vssd1 vssd1 vccd1 vccd1 _00292_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_7_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10641__S net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1017 net1020 vssd1 vssd1 vccd1 vccd1 net1017 sky130_fd_sc_hd__clkbuf_4
Xfanout1028 net1029 vssd1 vssd1 vccd1 vccd1 net1028 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07149__A2 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1039 net1071 vssd1 vssd1 vccd1 vccd1 net1039 sky130_fd_sc_hd__buf_2
XANTENNA__07516__A _02633_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_76_Right_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_126_2331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12970__CLK clknet_leaf_120_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_199_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_202_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12801_ clknet_leaf_17_clk _00393_ net1030 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[9\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_202_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_201_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13781_ clknet_leaf_68_clk _00016_ net1097 vssd1 vssd1 vccd1 vccd1 top.pad.button_control.noisy
+ sky130_fd_sc_hd__dfrtp_1
X_10993_ net843 _05027_ _05028_ net849 top.a1.dataIn\[7\] vssd1 vssd1 vccd1 vccd1
+ _05029_ sky130_fd_sc_hd__a32o_1
XANTENNA__09846__A1 _01584_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_201_148 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12732_ clknet_leaf_130_clk _00324_ net909 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[7\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_378 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06419__X _01558_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07321__A2 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_52_clk_A clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_194_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12663_ clknet_leaf_129_clk _00255_ net912 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[5\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10088__S net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_154_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_172_3030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11614_ _05484_ _05493_ _05495_ _05492_ vssd1 vssd1 vccd1 vccd1 _05497_ sky130_fd_sc_hd__or4b_2
XFILLER_0_65_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12594_ clknet_leaf_23_clk _00186_ net1021 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[3\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_85_Right_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_182_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10816__S net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11545_ _05427_ vssd1 vssd1 vccd1 vccd1 _05428_ sky130_fd_sc_hd__inv_2
XFILLER_0_163_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_576 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11476_ _05357_ _05330_ vssd1 vssd1 vccd1 vccd1 _05359_ sky130_fd_sc_hd__and2b_1
XFILLER_0_12_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_110_clk_A clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10427_ net1277 net151 net370 vssd1 vssd1 vccd1 vccd1 _00599_ sky130_fd_sc_hd__mux2_1
X_13215_ clknet_leaf_19_clk _00807_ net1026 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[22\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_150_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07388__A2 net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11184__A3 net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_150_2693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10358_ net1709 net153 net378 vssd1 vssd1 vccd1 vccd1 _00534_ sky130_fd_sc_hd__mux2_1
X_13146_ clknet_leaf_5_clk _00738_ net936 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[20\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_103_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_209_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10551__S net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13077_ clknet_leaf_29_clk _00669_ net1019 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[18\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_10289_ net1766 net165 net387 vssd1 vssd1 vccd1 vccd1 _00467_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_125_clk_A clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_94_Right_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12028_ _05894_ _05904_ _05898_ vssd1 vssd1 vccd1 vccd1 _05911_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_183_3192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_4_2__f_clk_X clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10695__A2 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_205_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07560__A2 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08528__Y _03655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06520_ _01657_ _01658_ vssd1 vssd1 vccd1 vccd1 _01659_ sky130_fd_sc_hd__nand2b_2
XTAP_TAPCELL_ROW_66_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07848__B1 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07312__A2 net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_201_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_157_2803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06451_ top.a1.instruction\[5\] _01473_ _01589_ vssd1 vssd1 vccd1 vccd1 _01590_ sky130_fd_sc_hd__a21o_1
XFILLER_0_201_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09170_ _04240_ _04241_ vssd1 vssd1 vccd1 vccd1 _04242_ sky130_fd_sc_hd__nor2_1
X_06382_ top.a1.instruction\[17\] top.a1.instruction\[18\] net782 vssd1 vssd1 vccd1
+ vccd1 _01521_ sky130_fd_sc_hd__and3b_2
XFILLER_0_113_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_173_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08121_ _03151_ _03181_ vssd1 vssd1 vccd1 vccd1 _03260_ sky130_fd_sc_hd__or2_2
XFILLER_0_7_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09359__Y _04420_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_122_clk clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_122_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__10726__S net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08052_ _03189_ _03190_ vssd1 vssd1 vccd1 vccd1 _03191_ sky130_fd_sc_hd__nand2_1
XANTENNA__09088__A _01546_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07003_ top.DUT.register\[11\]\[20\] net525 net518 top.DUT.register\[7\]\[20\] _02141_
+ vssd1 vssd1 vccd1 vccd1 _02142_ sky130_fd_sc_hd__a221o_1
XANTENNA__08974__A2_N net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06224__B net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07379__A2 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_77_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06587__B1 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_168_2965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10461__S net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08954_ net1237 net873 _02383_ net693 vssd1 vssd1 vccd1 vccd1 _00060_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_4_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1014_A net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07336__A _02443_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_205_3516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07905_ _03043_ vssd1 vssd1 vccd1 vccd1 _03044_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_90_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_205_3527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13828__1112 vssd1 vssd1 vccd1 vccd1 _13828__1112/HI net1112 sky130_fd_sc_hd__conb_1
X_08885_ _03315_ _03322_ vssd1 vssd1 vccd1 vccd1 _03995_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout474_A net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07836_ _02952_ _02973_ net824 vssd1 vssd1 vccd1 vccd1 _02975_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_108_2061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07551__A2 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12383__RESET_B net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_2072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07767_ top.DUT.register\[15\]\[2\] net706 net698 top.DUT.register\[31\]\[2\] vssd1
+ vssd1 vccd1 vccd1 _02906_ sky130_fd_sc_hd__a22o_1
XFILLER_0_79_643 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout262_X net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout641_A _01619_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout739_A _01624_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09506_ _04556_ _04557_ vssd1 vssd1 vccd1 vccd1 _04558_ sky130_fd_sc_hd__or2_1
XANTENNA__07839__B1 net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06718_ top.DUT.register\[25\]\[25\] net778 net769 top.DUT.register\[28\]\[25\] _01856_
+ vssd1 vssd1 vccd1 vccd1 _01857_ sky130_fd_sc_hd__a221o_1
XFILLER_0_78_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07698_ top.DUT.register\[6\]\[4\] net569 net541 top.DUT.register\[8\]\[4\] vssd1
+ vssd1 vccd1 vccd1 _02837_ sky130_fd_sc_hd__a22o_1
XFILLER_0_79_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07303__A2 net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_2261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06649_ _01764_ _01784_ vssd1 vssd1 vccd1 vccd1 _01788_ sky130_fd_sc_hd__nor2_1
XFILLER_0_164_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09437_ top.pc\[21\] _04478_ vssd1 vssd1 vccd1 vccd1 _04493_ sky130_fd_sc_hd__xnor2_1
XANTENNA__06511__B1 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout527_X net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout906_A net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09368_ top.pc\[17\] _04410_ vssd1 vssd1 vccd1 vccd1 _04428_ sky130_fd_sc_hd__and2_1
XFILLER_0_164_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08319_ net286 _03453_ vssd1 vssd1 vccd1 vccd1 _03454_ sky130_fd_sc_hd__nand2_2
XFILLER_0_164_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_1905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10636__S net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_543 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09299_ top.pc\[13\] _04352_ vssd1 vssd1 vccd1 vccd1 _04363_ sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_113_clk clknet_4_6__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_113_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_117_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_4_13__f_clk_X clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11330_ top.a1.dataIn\[22\] _05211_ top.a1.dataIn\[23\] vssd1 vssd1 vccd1 vccd1 _05213_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_62_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_97_Left_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11261_ net878 net880 _05148_ vssd1 vssd1 vccd1 vccd1 _05153_ sky130_fd_sc_hd__and3_1
XFILLER_0_104_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06290__A2 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13100__RESET_B net1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10212_ net190 net2197 net394 vssd1 vssd1 vccd1 vccd1 _00392_ sky130_fd_sc_hd__mux2_1
X_13000_ clknet_leaf_25_clk _00592_ net1008 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[15\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_30_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11192_ top.a1.data\[11\] net783 _05039_ vssd1 vssd1 vccd1 vccd1 _05103_ sky130_fd_sc_hd__o21a_1
XANTENNA__06578__B1 net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09007__D_N _03532_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10143_ net148 net1972 net609 vssd1 vssd1 vccd1 vccd1 _00343_ sky130_fd_sc_hd__mux2_1
XANTENNA__10371__S net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09445__B _04499_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_207_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_50_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07790__A2 net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10074_ net1636 net160 net617 vssd1 vssd1 vccd1 vccd1 _00276_ sky130_fd_sc_hd__mux2_1
XANTENNA_input35_A gpio_in[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06150__A net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_187_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_626 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13764_ clknet_leaf_100_clk _01335_ vssd1 vssd1 vccd1 vccd1 top.lcd.cnt_500hz\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__09295__A2 top.pc\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10976_ top.a1.halfData\[3\] net783 _05015_ net843 vssd1 vssd1 vccd1 vccd1 _05016_
+ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_48_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12715_ clknet_leaf_45_clk _00307_ net1065 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[6\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_167_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_167_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13695_ clknet_leaf_91_clk _01266_ vssd1 vssd1 vccd1 vccd1 net124 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_85_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06502__B1 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_139_2533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12646_ clknet_leaf_40_clk _00238_ net1053 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[4\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_104_clk clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_104_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__10546__S net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08255__B1 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12577_ clknet_leaf_17_clk _00169_ net964 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[2\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_142_217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11231__A _05120_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_152_2722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_152_2733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11528_ _05378_ _05410_ vssd1 vssd1 vccd1 vccd1 _05411_ sky130_fd_sc_hd__nor2_1
XFILLER_0_41_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwire272 _04121_ vssd1 vssd1 vccd1 vccd1 net272 sky130_fd_sc_hd__clkbuf_1
Xhold308 top.DUT.register\[26\]\[29\] vssd1 vssd1 vccd1 vccd1 net1424 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold319 top.DUT.register\[20\]\[4\] vssd1 vssd1 vccd1 vccd1 net1435 sky130_fd_sc_hd__dlygate4sd3_1
X_11459_ _05335_ _05341_ vssd1 vssd1 vccd1 vccd1 _05342_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_185_3221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_659 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06569__B1 net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_194_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10281__S net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07427__Y _02566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09355__B _04403_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13129_ clknet_leaf_52_clk _00721_ net1036 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[19\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07781__A2 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1008 top.DUT.register\[31\]\[25\] vssd1 vssd1 vccd1 vccd1 net2124 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1019 top.DUT.register\[16\]\[16\] vssd1 vssd1 vccd1 vccd1 net2135 sky130_fd_sc_hd__dlygate4sd3_1
X_08670_ _02007_ _03789_ vssd1 vssd1 vccd1 vccd1 _03790_ sky130_fd_sc_hd__xnor2_2
XANTENNA__08730__A1 _03334_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_163_2884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07533__A2 net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_163_2895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07621_ top.DUT.register\[16\]\[5\] net543 net511 top.DUT.register\[24\]\[5\] _02759_
+ vssd1 vssd1 vccd1 vccd1 _02760_ sky130_fd_sc_hd__a221o_1
XFILLER_0_108_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06741__B1 net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_177_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_200_3446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07552_ top.DUT.register\[21\]\[7\] net655 net738 top.DUT.register\[12\]\[7\] _02689_
+ vssd1 vssd1 vccd1 vccd1 _02691_ sky130_fd_sc_hd__a221o_1
XFILLER_0_76_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06503_ _01592_ _01596_ _01618_ vssd1 vssd1 vccd1 vccd1 _01642_ sky130_fd_sc_hd__and3_4
XTAP_TAPCELL_ROW_196_3383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_158_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07483_ top.DUT.register\[20\]\[14\] net566 net446 top.DUT.register\[1\]\[14\] _02621_
+ vssd1 vssd1 vccd1 vccd1 _02622_ sky130_fd_sc_hd__a221o_1
XANTENNA__11125__B net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_201_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09691__C1 _04725_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06219__B net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06434_ net896 top.a1.instruction\[5\] vssd1 vssd1 vccd1 vccd1 _01573_ sky130_fd_sc_hd__and2_1
X_09222_ _04287_ _04290_ vssd1 vssd1 vccd1 vccd1 _04291_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_173_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_146_556 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09153_ top.pc\[4\] _02857_ vssd1 vssd1 vccd1 vccd1 _04226_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06365_ net896 _01389_ _01390_ _01502_ vssd1 vssd1 vccd1 vccd1 _01504_ sky130_fd_sc_hd__or4b_1
XFILLER_0_99_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08246__B1 net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10456__S net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout222_A _04766_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08104_ _03242_ vssd1 vssd1 vccd1 vccd1 _03243_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_79_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_239 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09084_ top.a1.instruction\[9\] top.a1.instruction\[10\] _01573_ _04155_ vssd1 vssd1
+ vccd1 vccd1 _04159_ sky130_fd_sc_hd__and4_1
XFILLER_0_44_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_291 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06235__A top.ramload\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06296_ _01450_ _01330_ vssd1 vssd1 vccd1 vccd1 _01454_ sky130_fd_sc_hd__nor2_1
XFILLER_0_16_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08035_ _03173_ vssd1 vssd1 vccd1 vccd1 _03174_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10980__A top.a1.dataInTemp\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold820 top.DUT.register\[12\]\[22\] vssd1 vssd1 vccd1 vccd1 net1936 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold831 top.DUT.register\[18\]\[6\] vssd1 vssd1 vccd1 vccd1 net1947 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12345__A2 net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold842 top.DUT.register\[7\]\[13\] vssd1 vssd1 vccd1 vccd1 net1958 sky130_fd_sc_hd__dlygate4sd3_1
Xhold853 top.DUT.register\[29\]\[0\] vssd1 vssd1 vccd1 vccd1 net1969 sky130_fd_sc_hd__dlygate4sd3_1
Xhold864 top.DUT.register\[1\]\[0\] vssd1 vssd1 vccd1 vccd1 net1980 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08450__A net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold875 top.DUT.register\[19\]\[26\] vssd1 vssd1 vccd1 vccd1 net1991 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout591_A _04971_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout689_A net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold886 top.DUT.register\[21\]\[30\] vssd1 vssd1 vccd1 vccd1 net2002 sky130_fd_sc_hd__dlygate4sd3_1
Xhold897 top.DUT.register\[3\]\[1\] vssd1 vssd1 vccd1 vccd1 net2013 sky130_fd_sc_hd__dlygate4sd3_1
X_09986_ net243 net1803 net623 vssd1 vssd1 vccd1 vccd1 _00191_ sky130_fd_sc_hd__mux2_1
XANTENNA__07772__A2 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13171__CLK clknet_leaf_120_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08937_ net429 _04041_ _04044_ vssd1 vssd1 vccd1 vccd1 _04045_ sky130_fd_sc_hd__a21oi_4
XANTENNA__10108__A1 net156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout477_X net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06980__B1 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08868_ net319 _03652_ _03823_ net274 _03978_ vssd1 vssd1 vccd1 vccd1 _03979_ sky130_fd_sc_hd__a221o_1
XANTENNA__07524__A2 net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_91 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07819_ top.DUT.register\[30\]\[0\] net758 net727 top.DUT.register\[18\]\[0\] vssd1
+ vssd1 vccd1 vccd1 _02958_ sky130_fd_sc_hd__a22o_1
XFILLER_0_211_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08799_ _01877_ _03912_ vssd1 vssd1 vccd1 vccd1 _03913_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout644_X net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10830_ top.DUT.register\[28\]\[6\] net241 net474 vssd1 vssd1 vccd1 vccd1 _00991_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_211_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_184_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout811_X net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10761_ net1601 net270 net484 vssd1 vssd1 vccd1 vccd1 _00922_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_36_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12500_ clknet_leaf_111_clk _00092_ net989 vssd1 vssd1 vccd1 vccd1 top.pc\[12\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_109_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13480_ clknet_leaf_27_clk _01072_ net1010 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[30\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_10692_ net1983 net150 net340 vssd1 vssd1 vccd1 vccd1 _00855_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_180_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_101_1964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_180_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08237__B1 _03363_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12431_ clknet_leaf_93_clk _00027_ net994 vssd1 vssd1 vccd1 vccd1 top.ramaddr\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10366__S net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08344__B net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_671 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12362_ clknet_leaf_95_clk top.ru.next_FetchedData\[6\] net981 vssd1 vssd1 vccd1
+ vccd1 top.a1.dataIn\[6\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_23_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_384 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06799__B1 net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_134_2452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_2463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11313_ net879 _05120_ _05148_ _05196_ _05198_ vssd1 vssd1 vccd1 vccd1 _05199_ sky130_fd_sc_hd__a311o_1
XFILLER_0_160_570 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12293_ top.lcd.cnt_500hz\[14\] _06105_ vssd1 vssd1 vccd1 vccd1 _06107_ sky130_fd_sc_hd__or2_1
XFILLER_0_132_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_200_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09737__B1 net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11244_ top.a1.row1\[112\] _05132_ _05136_ top.a1.row1\[56\] _05134_ vssd1 vssd1
+ vccd1 vccd1 _05137_ sky130_fd_sc_hd__a221o_1
XFILLER_0_38_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11175_ top.a1.state\[2\] net587 vssd1 vssd1 vccd1 vccd1 _05098_ sky130_fd_sc_hd__nor2_1
XFILLER_0_100_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10126_ net207 net1958 net609 vssd1 vssd1 vccd1 vccd1 _00326_ sky130_fd_sc_hd__mux2_1
XFILLER_0_209_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_180_3140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_180_3151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10057_ net2186 net229 net615 vssd1 vssd1 vccd1 vccd1 _00259_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09735__A1_N net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09191__A _02723_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08712__B2 _03830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_187_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_259 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkload0_A clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13816_ net1101 vssd1 vssd1 vccd1 vccd1 gpio_out[3] sky130_fd_sc_hd__buf_2
XFILLER_0_85_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_187_478 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13747_ clknet_leaf_99_clk _01318_ vssd1 vssd1 vccd1 vccd1 top.lcd.cnt_20ms\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_10959_ net844 net784 _05001_ _04667_ _04997_ vssd1 vssd1 vccd1 vccd1 _05002_ sky130_fd_sc_hd__a32o_1
XANTENNA__07710__Y _02849_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13678_ clknet_leaf_91_clk _01254_ net996 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_14_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12629_ clknet_leaf_34_clk _00221_ net1040 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[4\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10276__S net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13827__1111 vssd1 vssd1 vccd1 vccd1 _13827__1111/HI net1111 sky130_fd_sc_hd__conb_1
XFILLER_0_143_548 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06150_ net900 vssd1 vssd1 vccd1 vccd1 _01393_ sky130_fd_sc_hd__inv_2
XFILLER_0_53_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold105 top.DUT.register\[14\]\[13\] vssd1 vssd1 vccd1 vccd1 net1221 sky130_fd_sc_hd__dlygate4sd3_1
Xhold116 _01364_ vssd1 vssd1 vccd1 vccd1 net1232 sky130_fd_sc_hd__dlygate4sd3_1
Xhold127 _01160_ vssd1 vssd1 vccd1 vccd1 net1243 sky130_fd_sc_hd__dlygate4sd3_1
Xhold138 top.DUT.register\[28\]\[31\] vssd1 vssd1 vccd1 vccd1 net1254 sky130_fd_sc_hd__dlygate4sd3_1
Xhold149 top.pad.button_control.r_counter\[1\] vssd1 vssd1 vccd1 vccd1 net1265 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08270__A net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_676 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout607 _04956_ vssd1 vssd1 vccd1 vccd1 net607 sky130_fd_sc_hd__buf_6
X_09840_ _04843_ _04851_ _04852_ _04151_ vssd1 vssd1 vccd1 vccd1 _04854_ sky130_fd_sc_hd__a31o_1
Xfanout618 _04954_ vssd1 vssd1 vccd1 vccd1 net618 sky130_fd_sc_hd__buf_4
Xfanout629 _04948_ vssd1 vssd1 vccd1 vccd1 net629 sky130_fd_sc_hd__buf_6
XFILLER_0_0_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_165_2924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07754__A2 net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08951__B2 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09771_ net826 _04395_ _04752_ top.a1.dataIn\[15\] vssd1 vssd1 vccd1 vccd1 _04792_
+ sky130_fd_sc_hd__a2bb2o_1
X_06983_ _02114_ _02116_ _02120_ _02121_ vssd1 vssd1 vccd1 vccd1 _02122_ sky130_fd_sc_hd__or4_1
X_08722_ _03476_ _03534_ _03676_ net279 _03839_ vssd1 vssd1 vccd1 vccd1 _03840_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_198_3412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07506__A2 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_198_3423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08653_ _03731_ _03773_ net290 vssd1 vssd1 vccd1 vccd1 _03774_ sky130_fd_sc_hd__mux2_1
XFILLER_0_178_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_105_2020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout172_A _04876_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07604_ top.DUT.register\[10\]\[6\] net770 net742 top.DUT.register\[2\]\[6\] vssd1
+ vssd1 vccd1 vccd1 _02743_ sky130_fd_sc_hd__a22o_1
X_08584_ _02614_ _03707_ vssd1 vssd1 vccd1 vccd1 _03708_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_138_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07535_ top.DUT.register\[30\]\[7\] net579 net459 top.DUT.register\[17\]\[7\] _02673_
+ vssd1 vssd1 vccd1 vccd1 _02674_ sky130_fd_sc_hd__a221o_1
XFILLER_0_76_443 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout437_A _01587_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07466_ top.DUT.register\[23\]\[15\] net672 net736 top.DUT.register\[16\]\[15\] _02604_
+ vssd1 vssd1 vccd1 vccd1 _02605_ sky130_fd_sc_hd__a221o_1
XFILLER_0_119_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06417_ top.DUT.register\[11\]\[30\] net525 net521 top.DUT.register\[10\]\[30\] vssd1
+ vssd1 vccd1 vccd1 _01556_ sky130_fd_sc_hd__a22o_1
XFILLER_0_45_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09205_ _04272_ _04273_ vssd1 vssd1 vccd1 vccd1 _04275_ sky130_fd_sc_hd__xnor2_1
XANTENNA__06493__A2 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07397_ top.DUT.register\[14\]\[9\] net583 net527 top.DUT.register\[26\]\[9\] vssd1
+ vssd1 vccd1 vccd1 _02536_ sky130_fd_sc_hd__a22o_1
XFILLER_0_60_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout604_A net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09975__S net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06348_ top.d_ready top.ru.state\[0\] net795 vssd1 vssd1 vccd1 vccd1 _00006_ sky130_fd_sc_hd__and3b_1
X_09136_ net806 _04201_ vssd1 vssd1 vccd1 vccd1 _04210_ sky130_fd_sc_hd__nor2_1
XFILLER_0_71_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09067_ _03936_ _04062_ _04141_ vssd1 vssd1 vccd1 vccd1 _04142_ sky130_fd_sc_hd__a21boi_4
XFILLER_0_114_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10914__S net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06279_ _01437_ _01439_ _01440_ _01441_ vssd1 vssd1 vccd1 vccd1 _01442_ sky130_fd_sc_hd__or4_4
XFILLER_0_130_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_116_2182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_2193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08018_ _02344_ _03153_ _03154_ _03156_ _01500_ vssd1 vssd1 vccd1 vccd1 _03157_ sky130_fd_sc_hd__o41a_4
XANTENNA__07993__A2 net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08180__A _01809_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold650 top.DUT.register\[11\]\[26\] vssd1 vssd1 vccd1 vccd1 net1766 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10329__A1 net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout594_X net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold661 top.DUT.register\[20\]\[0\] vssd1 vssd1 vccd1 vccd1 net1777 sky130_fd_sc_hd__dlygate4sd3_1
Xhold672 top.DUT.register\[20\]\[16\] vssd1 vssd1 vccd1 vccd1 net1788 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold683 top.DUT.register\[22\]\[15\] vssd1 vssd1 vccd1 vccd1 net1799 sky130_fd_sc_hd__dlygate4sd3_1
Xhold694 top.DUT.register\[7\]\[1\] vssd1 vssd1 vccd1 vccd1 net1810 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07745__A2 net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout761_X net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09969_ net1505 net174 net629 vssd1 vssd1 vccd1 vccd1 _00177_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout859_X net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12980_ clknet_leaf_55_clk _00572_ net1073 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[15\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_188_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11931_ _05758_ _05760_ _05792_ _05793_ _05789_ vssd1 vssd1 vccd1 vccd1 _05814_ sky130_fd_sc_hd__a221o_2
XFILLER_0_169_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06705__B1 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11862_ _05648_ _05676_ _05650_ vssd1 vssd1 vccd1 vccd1 _05745_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_200_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13601_ clknet_leaf_65_clk net1236 net1094 vssd1 vssd1 vccd1 vccd1 net93 sky130_fd_sc_hd__dfrtp_1
X_10813_ net192 net2106 net600 vssd1 vssd1 vccd1 vccd1 _00974_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11793_ _05655_ _05656_ _05643_ vssd1 vssd1 vccd1 vccd1 _05676_ sky130_fd_sc_hd__a21oi_2
XTAP_TAPCELL_ROW_45_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13532_ clknet_leaf_93_clk _01119_ net995 vssd1 vssd1 vccd1 vccd1 top.a1.data\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_10744_ net2000 net224 net421 vssd1 vssd1 vccd1 vccd1 _00905_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06427__X _01566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07130__B1 net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09670__A2 net139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_165_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13463_ clknet_leaf_128_clk _01055_ net913 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[30\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_11_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10096__S net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_180_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_608 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10675_ net1578 net207 net340 vssd1 vssd1 vccd1 vccd1 _00838_ sky130_fd_sc_hd__mux2_1
XFILLER_0_180_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12414_ clknet_leaf_103_clk top.ru.next_FetchedInstr\[26\] net976 vssd1 vssd1 vccd1
+ vccd1 top.a1.instruction\[26\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_35_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13394_ clknet_leaf_25_clk _00986_ net1014 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[28\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_211_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12345_ net2213 net904 net36 vssd1 vssd1 vccd1 vccd1 _01370_ sky130_fd_sc_hd__a21o_1
XFILLER_0_2_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_189_Left_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10824__S net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07984__A2 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12276_ top.lcd.cnt_500hz\[7\] _06094_ top.lcd.cnt_500hz\[8\] vssd1 vssd1 vccd1 vccd1
+ _06096_ sky130_fd_sc_hd__a21o_1
XFILLER_0_120_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12415__RESET_B net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11227_ net880 _01382_ vssd1 vssd1 vccd1 vccd1 _05120_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_56_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_208_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12190__B1 _05082_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07736__A2 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11158_ _01410_ _05085_ _05086_ _05087_ vssd1 vssd1 vccd1 vccd1 _01227_ sky130_fd_sc_hd__a31o_1
XANTENNA__06944__B1 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_147_2654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10109_ net1262 net154 net614 vssd1 vssd1 vccd1 vccd1 _00310_ sky130_fd_sc_hd__mux2_1
X_11089_ net66 net867 vssd1 vssd1 vccd1 vccd1 _05050_ sky130_fd_sc_hd__and2_1
XANTENNA__09125__S _04142_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11227__Y _05120_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_198_Left_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_172_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_160_2843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_159_Right_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_157_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11048__A2 net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_193_3342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13203__RESET_B net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07320_ top.DUT.register\[4\]\[12\] net667 net639 top.DUT.register\[8\]\[12\] _02458_
+ vssd1 vssd1 vccd1 vccd1 _02459_ sky130_fd_sc_hd__a221o_1
XANTENNA__11243__X _05136_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_190_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07251_ _02310_ _02389_ vssd1 vssd1 vccd1 vccd1 _02390_ sky130_fd_sc_hd__or2_1
XFILLER_0_73_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_143_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_619 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06202_ _01429_ _01431_ vssd1 vssd1 vccd1 vccd1 _00013_ sky130_fd_sc_hd__nand2_1
XFILLER_0_143_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07182_ top.DUT.register\[26\]\[10\] net527 _02320_ vssd1 vssd1 vccd1 vccd1 _02321_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_121_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_171_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09413__A2 _02679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_490 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10734__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09808__B _04471_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_721 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07975__A2 net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout404 net406 vssd1 vssd1 vccd1 vccd1 net404 sky130_fd_sc_hd__buf_4
XANTENNA__07188__B1 net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06232__B net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout426 net427 vssd1 vssd1 vccd1 vccd1 net426 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07727__A2 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09823_ _04487_ net486 net401 top.a1.dataIn\[20\] net397 vssd1 vssd1 vccd1 vccd1
+ _04839_ sky130_fd_sc_hd__a221o_2
Xfanout437 _01587_ vssd1 vssd1 vccd1 vccd1 net437 sky130_fd_sc_hd__clkbuf_4
Xfanout448 _01562_ vssd1 vssd1 vccd1 vccd1 net448 sky130_fd_sc_hd__buf_4
XANTENNA__06800__X _01939_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout459 net460 vssd1 vssd1 vccd1 vccd1 net459 sky130_fd_sc_hd__buf_4
XANTENNA__06935__B1 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout387_A net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09754_ top.a1.dataIn\[13\] _04752_ _04362_ net826 vssd1 vssd1 vccd1 vccd1 _04777_
+ sky130_fd_sc_hd__o2bb2a_1
X_06966_ top.DUT.register\[11\]\[23\] net526 _02102_ _02104_ vssd1 vssd1 vccd1 vccd1
+ _02105_ sky130_fd_sc_hd__a211o_1
X_08705_ net279 _03651_ _03823_ net283 _03819_ vssd1 vssd1 vccd1 vccd1 _03824_ sky130_fd_sc_hd__o221a_1
X_09685_ _04709_ _04720_ net34 vssd1 vssd1 vccd1 vccd1 _04721_ sky130_fd_sc_hd__o21a_1
XFILLER_0_146_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout554_A _01535_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_732 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06897_ top.DUT.register\[7\]\[18\] net661 net637 top.DUT.register\[6\]\[18\] vssd1
+ vssd1 vccd1 vccd1 _02036_ sky130_fd_sc_hd__a22o_1
XFILLER_0_55_80 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_87_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_93_clk clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_93_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_87_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_126_Right_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08636_ net274 _03577_ _03757_ net285 vssd1 vssd1 vccd1 vccd1 _03758_ sky130_fd_sc_hd__a22o_1
XFILLER_0_178_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_179_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_178_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10909__S net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout342_X net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08567_ _02655_ net431 net499 _02654_ vssd1 vssd1 vccd1 vccd1 _03692_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout721_A _01635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_202_Left_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07518_ _02656_ vssd1 vssd1 vccd1 vccd1 _02657_ sky130_fd_sc_hd__inv_2
X_08498_ net320 _03625_ _03621_ vssd1 vssd1 vccd1 vccd1 _03626_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_9_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07112__B1 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07449_ top.DUT.register\[30\]\[15\] net580 net536 top.DUT.register\[19\]\[15\] _02587_
+ vssd1 vssd1 vccd1 vccd1 _02588_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_118_2211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout607_X net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_2222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06407__B top.a1.instruction\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_40_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10460_ net150 net2096 net366 vssd1 vssd1 vccd1 vccd1 _00631_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_40_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09119_ _04191_ _04193_ vssd1 vssd1 vccd1 vccd1 _04194_ sky130_fd_sc_hd__nor2_1
X_10391_ net1518 net152 net376 vssd1 vssd1 vccd1 vccd1 _00566_ sky130_fd_sc_hd__mux2_1
XFILLER_0_161_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10644__S net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_131_2411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12130_ _06001_ _06004_ _05995_ vssd1 vssd1 vccd1 vccd1 _06013_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07966__A2 net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout976_X net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_211_Left_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12061_ _05927_ _05933_ _05934_ vssd1 vssd1 vccd1 vccd1 _05944_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_3_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold480 top.DUT.register\[19\]\[8\] vssd1 vssd1 vccd1 vccd1 net1596 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07179__B1 net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold491 top.DUT.register\[29\]\[16\] vssd1 vssd1 vccd1 vccd1 net1607 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08915__A1 net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11012_ net887 wb.prev_BUSY_O net840 vssd1 vssd1 vccd1 vccd1 _05043_ sky130_fd_sc_hd__and3b_1
XANTENNA__06926__B1 net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout960 net962 vssd1 vssd1 vccd1 vccd1 net960 sky130_fd_sc_hd__clkbuf_2
Xfanout971 net1007 vssd1 vssd1 vccd1 vccd1 net971 sky130_fd_sc_hd__clkbuf_2
Xfanout982 net983 vssd1 vssd1 vccd1 vccd1 net982 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_205_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout993 net1007 vssd1 vssd1 vccd1 vccd1 net993 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_129_2384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13826__1110 vssd1 vssd1 vccd1 vccd1 _13826__1110/HI net1110 sky130_fd_sc_hd__conb_1
X_12963_ clknet_leaf_53_clk _00555_ net1076 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[14\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1180 top.DUT.register\[16\]\[6\] vssd1 vssd1 vccd1 vccd1 net2296 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_84_clk clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_84_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_87_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1191 top.DUT.register\[13\]\[28\] vssd1 vssd1 vccd1 vccd1 net2307 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_206_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11914_ _05796_ vssd1 vssd1 vccd1 vccd1 _05797_ sky130_fd_sc_hd__inv_2
XFILLER_0_99_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_200_500 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12894_ clknet_leaf_20_clk _00486_ net1028 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[12\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_142_2573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07351__B1 net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_169_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11845_ top.a1.dataIn\[6\] net130 _05718_ vssd1 vssd1 vccd1 vccd1 _05728_ sky130_fd_sc_hd__and3_1
XANTENNA__10819__S net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09628__C1 _04668_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08085__A _02944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11776_ _05623_ _05658_ vssd1 vssd1 vccd1 vccd1 _05659_ sky130_fd_sc_hd__xnor2_2
XTAP_TAPCELL_ROW_175_3072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13515_ clknet_leaf_45_clk _01107_ net1069 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[31\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11223__B net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_684 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10727_ net1397 net141 net335 vssd1 vssd1 vccd1 vccd1 _00888_ sky130_fd_sc_hd__mux2_1
XFILLER_0_165_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13446_ clknet_leaf_33_clk _01038_ net1046 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[29\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08372__X _03505_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10658_ net152 net2015 net345 vssd1 vssd1 vccd1 vccd1 _00822_ sky130_fd_sc_hd__mux2_1
Xclkload14 clknet_leaf_119_clk vssd1 vssd1 vccd1 vccd1 clkload14/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_35_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload25 clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 clkload25/Y sky130_fd_sc_hd__clkinv_2
Xclkload36 clknet_leaf_109_clk vssd1 vssd1 vccd1 vccd1 clkload36/Y sky130_fd_sc_hd__inv_8
XANTENNA__10554__S net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload47 clknet_leaf_82_clk vssd1 vssd1 vccd1 vccd1 clkload47/Y sky130_fd_sc_hd__inv_6
X_13377_ clknet_leaf_19_clk _00969_ net1027 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[27\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_10589_ net1471 net164 net352 vssd1 vssd1 vccd1 vccd1 _00755_ sky130_fd_sc_hd__mux2_1
Xclkload58 clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 clkload58/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_140_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload69 clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 clkload69/Y sky130_fd_sc_hd__bufinv_16
X_12328_ top.pad.button_control.r_counter\[10\] _06127_ net791 vssd1 vssd1 vccd1 vccd1
+ _06129_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07429__A _02544_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09159__A1 _04216_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12259_ top.lcd.cnt_500hz\[0\] net686 vssd1 vssd1 vccd1 vccd1 _01335_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_71_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06917__B1 net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06820_ top.DUT.register\[4\]\[17\] net668 _01951_ _01954_ _01958_ vssd1 vssd1 vccd1
+ vccd1 _01959_ sky130_fd_sc_hd__a2111o_1
X_06751_ top.DUT.register\[14\]\[24\] net586 net506 top.DUT.register\[27\]\[24\] vssd1
+ vssd1 vccd1 vccd1 _01890_ sky130_fd_sc_hd__a22o_1
XFILLER_0_211_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_75_clk clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_75_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__09331__A1 net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06682_ _01815_ _01817_ _01819_ _01820_ vssd1 vssd1 vccd1 vccd1 _01821_ sky130_fd_sc_hd__or4_1
X_09470_ top.pc\[23\] _04514_ vssd1 vssd1 vccd1 vccd1 _04524_ sky130_fd_sc_hd__xor2_1
XANTENNA__08547__X _03673_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07342__B1 net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08421_ _03551_ vssd1 vssd1 vccd1 vccd1 _03552_ sky130_fd_sc_hd__inv_2
XFILLER_0_203_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_wire408_X net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06696__A2 net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10729__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_176_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_176_768 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08352_ _02851_ _03445_ _02850_ vssd1 vssd1 vccd1 vccd1 _03486_ sky130_fd_sc_hd__a21o_1
XANTENNA__07611__B _02749_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_40 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07303_ top.DUT.register\[14\]\[12\] net583 net539 top.DUT.register\[8\]\[12\] _02441_
+ vssd1 vssd1 vccd1 vccd1 _02442_ sky130_fd_sc_hd__a221o_1
XANTENNA__11133__B net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08283_ net276 _03417_ _03418_ vssd1 vssd1 vccd1 vccd1 _03419_ sky130_fd_sc_hd__o21a_1
XFILLER_0_190_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06227__B net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload8 clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 clkload8/Y sky130_fd_sc_hd__clkinv_8
XFILLER_0_27_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09378__X _04438_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07234_ top.DUT.register\[20\]\[10\] net663 net702 top.DUT.register\[3\]\[10\] _02367_
+ vssd1 vssd1 vccd1 vccd1 _02373_ sky130_fd_sc_hd__a221o_1
XFILLER_0_54_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_687 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07165_ _02289_ _02290_ _02294_ _02303_ vssd1 vssd1 vccd1 vccd1 _02304_ sky130_fd_sc_hd__or4_4
XFILLER_0_131_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10464__S net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1044_A net1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07096_ top.DUT.register\[8\]\[16\] net540 net460 top.DUT.register\[17\]\[16\] vssd1
+ vssd1 vccd1 vccd1 _02235_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_113_2141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06620__A2 net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout201 _04841_ vssd1 vssd1 vccd1 vccd1 net201 sky130_fd_sc_hd__clkbuf_2
Xfanout212 net214 vssd1 vssd1 vccd1 vccd1 net212 sky130_fd_sc_hd__buf_2
Xfanout223 _04805_ vssd1 vssd1 vccd1 vccd1 net223 sky130_fd_sc_hd__buf_2
Xfanout234 _05475_ vssd1 vssd1 vccd1 vccd1 net234 sky130_fd_sc_hd__buf_2
XANTENNA_fanout671_A _01597_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout245 net246 vssd1 vssd1 vccd1 vccd1 net245 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_208_3569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout256 _04737_ vssd1 vssd1 vccd1 vccd1 net256 sky130_fd_sc_hd__buf_1
X_09806_ net1268 net205 net634 vssd1 vssd1 vccd1 vccd1 _00139_ sky130_fd_sc_hd__mux2_1
Xfanout267 _04726_ vssd1 vssd1 vccd1 vccd1 net267 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_5_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout289 net294 vssd1 vssd1 vccd1 vccd1 net289 sky130_fd_sc_hd__clkbuf_4
X_07998_ top.DUT.register\[8\]\[31\] net641 net757 top.DUT.register\[1\]\[31\] _03136_
+ vssd1 vssd1 vccd1 vccd1 _03137_ sky130_fd_sc_hd__a221o_1
XFILLER_0_198_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07581__B1 net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09841__X _04855_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09737_ _03617_ net403 net488 _04762_ vssd1 vssd1 vccd1 vccd1 _04763_ sky130_fd_sc_hd__o211a_1
X_06949_ top.DUT.register\[26\]\[21\] net753 _02073_ _02078_ _02087_ vssd1 vssd1 vccd1
+ vccd1 _02088_ sky130_fd_sc_hd__a2111oi_2
Xclkbuf_leaf_66_clk clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_66_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout557_X net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_2_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09668_ _04194_ _04704_ vssd1 vssd1 vccd1 vccd1 _04705_ sky130_fd_sc_hd__nor2_1
XFILLER_0_179_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08619_ _02263_ net499 _03736_ net436 _03738_ vssd1 vssd1 vccd1 vccd1 _03742_ sky130_fd_sc_hd__a221o_1
XANTENNA__06687__A2 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10639__S net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09599_ net333 _04644_ vssd1 vssd1 vccd1 vccd1 _04645_ sky130_fd_sc_hd__xor2_1
XANTENNA_fanout724_X net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11630_ _05474_ _05479_ net234 vssd1 vssd1 vccd1 vccd1 _05513_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_65_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_194_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11561_ _05443_ vssd1 vssd1 vccd1 vccd1 _05444_ sky130_fd_sc_hd__inv_2
XFILLER_0_181_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08904__Y _04013_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13300_ clknet_leaf_55_clk _00892_ net1031 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[25\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_10512_ net2014 net225 net360 vssd1 vssd1 vccd1 vccd1 _00681_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_21_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11492_ _05360_ _05365_ _05373_ vssd1 vssd1 vccd1 vccd1 _05375_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_107_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13231_ clknet_leaf_22_clk _00823_ net1035 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[22\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_150_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10374__S net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10443_ net207 net1835 net367 vssd1 vssd1 vccd1 vccd1 _00614_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13162_ clknet_leaf_118_clk _00754_ net956 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[20\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_150_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_184 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06153__A top.a1.dataIn\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10374_ net1556 net214 net373 vssd1 vssd1 vccd1 vccd1 _00549_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12113_ _05986_ _05991_ _05992_ vssd1 vssd1 vccd1 vccd1 _05996_ sky130_fd_sc_hd__nand3_1
XANTENNA__06611__A2 net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13093_ clknet_leaf_35_clk _00685_ net1041 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[18\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_12044_ _05906_ _05908_ _05914_ _05926_ vssd1 vssd1 vccd1 vccd1 _05927_ sky130_fd_sc_hd__a31oi_2
XTAP_TAPCELL_ROW_53_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_144_2602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_2613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07572__B1 net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout790 _06112_ vssd1 vssd1 vccd1 vccd1 net790 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_189_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_57_clk clknet_4_12__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_57_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__09313__A1 net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_177_3101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09911__B _04620_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12946_ clknet_leaf_25_clk _00538_ net1014 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[14\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_62_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11120__A1 net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08808__A net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09864__A2 net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07712__A net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06678__A2 net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10549__S net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12877_ clknet_leaf_50_clk _00469_ net1058 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[11\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_158_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11828_ _05650_ _05677_ _05706_ vssd1 vssd1 vccd1 vccd1 _05711_ sky130_fd_sc_hd__or3b_2
XTAP_TAPCELL_ROW_190_3301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_173_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_117_Left_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11759_ _05640_ _05641_ vssd1 vssd1 vccd1 vccd1 _05642_ sky130_fd_sc_hd__nor2_1
XFILLER_0_83_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06615__X _01754_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_155_2764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_155_2775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08543__A net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload103 clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 clkload103/Y sky130_fd_sc_hd__inv_8
XFILLER_0_24_630 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10284__S net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13429_ clknet_leaf_29_clk _01021_ net1019 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[29\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06850__A2 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_302 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_188_3263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_58 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09063__D_N _03539_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08970_ _01829_ net692 net1229 net876 vssd1 vssd1 vccd1 vccd1 _00076_ sky130_fd_sc_hd__a2bb2o_1
X_07921_ _02544_ _02567_ vssd1 vssd1 vccd1 vccd1 _03060_ sky130_fd_sc_hd__nand2b_1
XANTENNA__09001__B1 _03454_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_126_Left_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07852_ top.DUT.register\[20\]\[0\] net564 net539 top.DUT.register\[8\]\[0\] vssd1
+ vssd1 vccd1 vccd1 _02991_ sky130_fd_sc_hd__a22o_1
XFILLER_0_194_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06803_ top.DUT.register\[14\]\[17\] net731 net636 top.DUT.register\[6\]\[17\] vssd1
+ vssd1 vccd1 vccd1 _01942_ sky130_fd_sc_hd__a22o_1
Xinput1 ACK_I vssd1 vssd1 vccd1 vccd1 net1 sky130_fd_sc_hd__clkbuf_2
X_07783_ _02915_ _02917_ _02919_ _02921_ vssd1 vssd1 vccd1 vccd1 _02922_ sky130_fd_sc_hd__or4_4
Xclkbuf_leaf_48_clk clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_48_clk
+ sky130_fd_sc_hd__clkbuf_8
X_09522_ top.pc\[26\] _04560_ vssd1 vssd1 vccd1 vccd1 _04573_ sky130_fd_sc_hd__or2_1
X_06734_ net808 net415 net438 vssd1 vssd1 vccd1 vccd1 _01873_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_84_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_203_3488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07315__B1 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10967__B _04998_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09855__A2 net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09453_ _04506_ _04507_ vssd1 vssd1 vccd1 vccd1 _04508_ sky130_fd_sc_hd__or2_1
X_06665_ top.DUT.register\[19\]\[26\] net537 net514 top.DUT.register\[24\]\[26\] vssd1
+ vssd1 vccd1 vccd1 _01804_ sky130_fd_sc_hd__a22o_1
XANTENNA__10459__S net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout252_A _04741_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_149_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08404_ _03535_ vssd1 vssd1 vccd1 vccd1 _03536_ sky130_fd_sc_hd__inv_2
X_09384_ net133 _04435_ _04443_ net900 vssd1 vssd1 vccd1 vccd1 _04444_ sky130_fd_sc_hd__o211a_1
XPHY_EDGE_ROW_135_Left_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_191_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06596_ top.DUT.register\[29\]\[28\] net725 _01730_ _01734_ vssd1 vssd1 vccd1 vccd1
+ _01735_ sky130_fd_sc_hd__a211o_1
XFILLER_0_136_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08335_ net297 _03468_ vssd1 vssd1 vccd1 vccd1 _03469_ sky130_fd_sc_hd__nand2_1
XFILLER_0_19_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12518__RESET_B net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout138_X net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout517_A _01558_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08266_ net274 _03395_ _03401_ net286 vssd1 vssd1 vccd1 vccd1 _03402_ sky130_fd_sc_hd__a22o_1
XANTENNA__07094__A2 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_490 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07217_ _02340_ _02355_ vssd1 vssd1 vccd1 vccd1 _02356_ sky130_fd_sc_hd__and2_1
XFILLER_0_131_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06841__A2 net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08197_ _03164_ _03182_ vssd1 vssd1 vccd1 vccd1 _03335_ sky130_fd_sc_hd__or2_1
XFILLER_0_104_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09983__S net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07148_ top.DUT.register\[7\]\[11\] net659 net714 top.DUT.register\[27\]\[11\] vssd1
+ vssd1 vccd1 vccd1 _02287_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_95_1866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_1877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout886_A top.ru.state\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07079_ _02208_ _02217_ vssd1 vssd1 vccd1 vccd1 _02218_ sky130_fd_sc_hd__or2_4
XFILLER_0_140_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_144_Left_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08900__B _04008_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10090_ net2109 net228 net612 vssd1 vssd1 vccd1 vccd1 _00291_ sky130_fd_sc_hd__mux2_1
Xfanout1007 net1098 vssd1 vssd1 vccd1 vccd1 net1007 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_7_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1018 net1020 vssd1 vssd1 vccd1 vccd1 net1018 sky130_fd_sc_hd__clkbuf_4
Xfanout1029 net1039 vssd1 vssd1 vccd1 vccd1 net1029 sky130_fd_sc_hd__buf_2
XANTENNA_fanout674_X net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_39_clk clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_39_clk
+ sky130_fd_sc_hd__clkbuf_8
X_12800_ clknet_leaf_17_clk _00392_ net1030 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[9\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_13780_ clknet_leaf_69_clk _01351_ net1097 vssd1 vssd1 vccd1 vccd1 top.pad.count\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_10992_ top.a1.dataInTemp\[7\] net785 vssd1 vssd1 vccd1 vccd1 _05028_ sky130_fd_sc_hd__or2_1
XANTENNA__11102__A1 net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12731_ clknet_leaf_119_clk _00323_ net931 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[7\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10369__S net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_153_Left_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_195_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_519 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12662_ clknet_leaf_3_clk _00254_ net941 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[5\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_182_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_172_3020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11613_ _05495_ _05492_ vssd1 vssd1 vccd1 vccd1 _05496_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_172_3031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12593_ clknet_leaf_108_clk _00185_ net977 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[3\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_182_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11544_ _05360_ _05422_ vssd1 vssd1 vccd1 vccd1 _05427_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07085__A2 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06832__A2 net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_2494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11475_ _05293_ _05329_ vssd1 vssd1 vccd1 vccd1 _05358_ sky130_fd_sc_hd__or2_1
X_13214_ clknet_leaf_54_clk _00806_ net1037 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[22\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_10426_ net1576 net155 net371 vssd1 vssd1 vccd1 vccd1 _00598_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_162_Left_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13145_ clknet_leaf_15_clk _00737_ net961 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[20\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_209_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10357_ net2307 net156 net378 vssd1 vssd1 vccd1 vccd1 _00533_ sky130_fd_sc_hd__mux2_1
XANTENNA__10832__S net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_150_2694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07793__B1 net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13076_ clknet_leaf_57_clk _00668_ net1075 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[18\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10288_ net1334 net169 net386 vssd1 vssd1 vccd1 vccd1 _00466_ sky130_fd_sc_hd__mux2_1
X_12027_ _05894_ _05898_ _05904_ vssd1 vssd1 vccd1 vccd1 _05910_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_183_3193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07545__B1 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09922__A net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06899__A2 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_171_Left_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11235__Y _05128_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12929_ clknet_leaf_17_clk _00521_ net1030 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[13\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10279__S net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_186_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_158_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_157_2804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06450_ top.a1.instruction\[6\] _01474_ vssd1 vssd1 vccd1 vccd1 _01589_ sky130_fd_sc_hd__and2_2
XFILLER_0_200_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12611__RESET_B net1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06381_ top.DUT.register\[22\]\[30\] net576 net573 top.DUT.register\[23\]\[30\] _01515_
+ vssd1 vssd1 vccd1 vccd1 _01520_ sky130_fd_sc_hd__a221o_1
XFILLER_0_7_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08120_ _03151_ _03181_ vssd1 vssd1 vccd1 vccd1 _03259_ sky130_fd_sc_hd__nor2_2
XANTENNA__08273__A1 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07076__A2 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10080__A1 net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06284__B1 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08051_ _01678_ net328 vssd1 vssd1 vccd1 vccd1 _03190_ sky130_fd_sc_hd__nand2_1
XFILLER_0_113_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_153_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_180_Left_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07002_ top.DUT.register\[3\]\[20\] net554 net529 top.DUT.register\[26\]\[20\] vssd1
+ vssd1 vccd1 vccd1 _02141_ sky130_fd_sc_hd__a22o_1
XFILLER_0_102_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_2100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09773__A1 _04403_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09773__B2 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10742__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08953_ _02566_ _04050_ top.ramstore\[9\] net873 vssd1 vssd1 vccd1 vccd1 _00059_
+ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_168_2966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07904_ _03041_ _03042_ vssd1 vssd1 vccd1 vccd1 _03043_ sky130_fd_sc_hd__nand2b_2
XTAP_TAPCELL_ROW_4_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_205_3517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07336__B _02452_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08884_ net296 _03676_ _03677_ net325 vssd1 vssd1 vccd1 vccd1 _03994_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_90_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_205_3528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07536__B1 net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06240__B net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1007_A net1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07000__A2 net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07835_ _02953_ net408 net823 vssd1 vssd1 vccd1 vccd1 _02974_ sky130_fd_sc_hd__mux2_2
XANTENNA_fanout467_A net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_2062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_211_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_108_2073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07766_ top.DUT.register\[30\]\[2\] net758 net754 top.DUT.register\[1\]\[2\] vssd1
+ vssd1 vccd1 vccd1 _02905_ sky130_fd_sc_hd__a22o_1
XFILLER_0_154_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_655 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09505_ top.pc\[24\] _04521_ top.pc\[25\] vssd1 vssd1 vccd1 vccd1 _04557_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06717_ top.DUT.register\[22\]\[25\] net647 net714 top.DUT.register\[27\]\[25\] _01855_
+ vssd1 vssd1 vccd1 vccd1 _01856_ sky130_fd_sc_hd__a221o_1
XFILLER_0_154_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_195_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout634_A _04714_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07697_ top.DUT.register\[25\]\[4\] net457 net449 top.DUT.register\[21\]\[4\] _02835_
+ vssd1 vssd1 vccd1 vccd1 _02836_ sky130_fd_sc_hd__a221o_1
XFILLER_0_78_176 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_149_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_327 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09436_ net901 top.pc\[20\] _04481_ _04492_ net891 vssd1 vssd1 vccd1 vccd1 _00100_
+ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_121_2262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06648_ _01786_ vssd1 vssd1 vccd1 vccd1 _01787_ sky130_fd_sc_hd__inv_2
XFILLER_0_164_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09367_ net899 top.pc\[16\] _04427_ net892 vssd1 vssd1 vccd1 vccd1 _00096_ sky130_fd_sc_hd__o211a_1
XANTENNA__10917__S net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06579_ top.DUT.register\[22\]\[28\] net577 net521 top.DUT.register\[10\]\[28\] vssd1
+ vssd1 vccd1 vccd1 _01718_ sky130_fd_sc_hd__a22o_1
XFILLER_0_170_70 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08318_ _03174_ _03451_ net311 vssd1 vssd1 vccd1 vccd1 _03453_ sky130_fd_sc_hd__mux2_1
XFILLER_0_164_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07067__A2 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_1906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_760 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09298_ _04360_ _04361_ vssd1 vssd1 vccd1 vccd1 _04362_ sky130_fd_sc_hd__or2_1
XFILLER_0_117_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_555 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06814__A2 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08249_ net423 _03377_ _03385_ _03334_ _03383_ vssd1 vssd1 vccd1 vccd1 _03386_ sky130_fd_sc_hd__a221o_1
XANTENNA__08451__A2_N net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_279 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11260_ net1269 net813 _05152_ net1078 vssd1 vssd1 vccd1 vccd1 _01264_ sky130_fd_sc_hd__o211a_1
XFILLER_0_15_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09213__B1 net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout889_X net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11020__B1 _05044_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10211_ net199 net2050 net394 vssd1 vssd1 vccd1 vccd1 _00391_ sky130_fd_sc_hd__mux2_1
XANTENNA__08567__A2 net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10652__S net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11191_ net1226 net587 net473 _05102_ vssd1 vssd1 vccd1 vccd1 _01245_ sky130_fd_sc_hd__a22o_1
XFILLER_0_101_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08630__B net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10142_ net152 net2172 net610 vssd1 vssd1 vccd1 vccd1 _00342_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_50_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13140__RESET_B net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10073_ top.DUT.register\[5\]\[26\] net165 net618 vssd1 vssd1 vccd1 vccd1 _00275_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__07527__B1 net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input28_A DAT_I[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13832_ net1116 vssd1 vssd1 vccd1 vccd1 gpio_out[31] sky130_fd_sc_hd__buf_2
XANTENNA__08358__A _03342_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_187_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10099__S net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_186_126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_463 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13763_ clknet_leaf_72_clk _01334_ vssd1 vssd1 vccd1 vccd1 top.lcd.currentState\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_10975_ top.a1.dataInTemp\[3\] net785 vssd1 vssd1 vccd1 vccd1 _05015_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_48_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12714_ clknet_leaf_118_clk _00306_ net955 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[6\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_636 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13694_ clknet_leaf_89_clk _01265_ vssd1 vssd1 vccd1 vccd1 net123 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_167_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12645_ clknet_leaf_35_clk _00237_ net1040 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[4\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_139_2534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10827__S net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_150_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08255__A1 net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08093__A _03230_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08255__B2 _03391_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12576_ clknet_leaf_80_clk _00168_ net1072 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[2\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xwire240 _05469_ vssd1 vssd1 vccd1 vccd1 net240 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_142_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_152_2723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11527_ _05376_ _05401_ vssd1 vssd1 vccd1 vccd1 _05410_ sky130_fd_sc_hd__xnor2_1
XANTENNA__11231__B _05123_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06805__A2 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold309 top.DUT.register\[9\]\[5\] vssd1 vssd1 vccd1 vccd1 net1425 sky130_fd_sc_hd__dlygate4sd3_1
X_11458_ _05338_ _05339_ vssd1 vssd1 vccd1 vccd1 _05341_ sky130_fd_sc_hd__nor2_1
XFILLER_0_7_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13228__RESET_B net1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_185_3222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10409_ net1448 net212 net369 vssd1 vssd1 vccd1 vccd1 _00581_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_295 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11389_ top.a1.dataIn\[27\] _05271_ _05269_ vssd1 vssd1 vccd1 vccd1 _05272_ sky130_fd_sc_hd__mux2_1
XANTENNA__07766__B1 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13128_ clknet_leaf_7_clk _00720_ net946 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[19\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07230__A2 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06341__A net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_175_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_187_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13059_ clknet_leaf_49_clk _00651_ net1060 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[17\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1009 top.DUT.register\[15\]\[11\] vssd1 vssd1 vccd1 vccd1 net2125 sky130_fd_sc_hd__dlygate4sd3_1
X_07620_ top.DUT.register\[2\]\[5\] net559 net539 top.DUT.register\[8\]\[5\] vssd1
+ vssd1 vccd1 vccd1 _02759_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_163_2885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09371__B _04420_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_163_2896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_200_3447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07551_ top.DUT.register\[28\]\[7\] net766 net726 top.DUT.register\[18\]\[7\] vssd1
+ vssd1 vccd1 vccd1 _02690_ sky130_fd_sc_hd__a22o_1
XFILLER_0_159_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06502_ top.DUT.register\[22\]\[30\] net649 net763 top.DUT.register\[9\]\[30\] vssd1
+ vssd1 vccd1 vccd1 _01641_ sky130_fd_sc_hd__a22o_1
XFILLER_0_75_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_196_3384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08494__A1 _02880_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07297__A2 net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07482_ top.DUT.register\[12\]\[14\] net533 net520 top.DUT.register\[10\]\[14\] vssd1
+ vssd1 vccd1 vccd1 _02621_ sky130_fd_sc_hd__a22o_1
XFILLER_0_174_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09691__B1 net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09221_ _04288_ _04289_ vssd1 vssd1 vccd1 vccd1 _04290_ sky130_fd_sc_hd__nor2_1
X_06433_ _01571_ vssd1 vssd1 vccd1 vccd1 _01572_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_17_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10737__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_173_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_161_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09152_ top.pc\[3\] _02904_ _04213_ vssd1 vssd1 vccd1 vccd1 _04225_ sky130_fd_sc_hd__a21oi_1
X_06364_ net896 top.a1.instruction\[5\] top.a1.instruction\[6\] _01502_ vssd1 vssd1
+ vccd1 vccd1 _01503_ sky130_fd_sc_hd__and4b_2
XFILLER_0_133_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_173_376 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_161_527 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08103_ _03240_ _03241_ vssd1 vssd1 vccd1 vccd1 _03242_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_79_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11141__B net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09083_ top.a1.instruction\[24\] top.a1.instruction\[25\] top.a1.instruction\[26\]
+ top.a1.instruction\[27\] vssd1 vssd1 vccd1 vccd1 _04158_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_79_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06295_ top.lcd.nextState\[0\] top.lcd.currentState\[0\] net815 vssd1 vssd1 vccd1
+ vccd1 _01453_ sky130_fd_sc_hd__mux2_1
XFILLER_0_140_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06235__B net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08034_ net276 _03172_ vssd1 vssd1 vccd1 vccd1 _03173_ sky130_fd_sc_hd__or2_1
Xhold810 top.DUT.register\[17\]\[5\] vssd1 vssd1 vccd1 vccd1 net1926 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold821 top.DUT.register\[9\]\[4\] vssd1 vssd1 vccd1 vccd1 net1937 sky130_fd_sc_hd__dlygate4sd3_1
Xhold832 top.DUT.register\[16\]\[29\] vssd1 vssd1 vccd1 vccd1 net1948 sky130_fd_sc_hd__dlygate4sd3_1
Xhold843 top.DUT.register\[9\]\[28\] vssd1 vssd1 vccd1 vccd1 net1959 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09746__A1 top.a1.dataIn\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10472__S net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold854 top.DUT.register\[17\]\[21\] vssd1 vssd1 vccd1 vccd1 net1970 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07757__B1 net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold865 top.DUT.register\[12\]\[18\] vssd1 vssd1 vccd1 vccd1 net1981 sky130_fd_sc_hd__dlygate4sd3_1
Xhold876 top.DUT.register\[27\]\[9\] vssd1 vssd1 vccd1 vccd1 net1992 sky130_fd_sc_hd__dlygate4sd3_1
Xhold887 top.DUT.register\[22\]\[22\] vssd1 vssd1 vccd1 vccd1 net2003 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_51_clk_A clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07221__A2 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold898 top.DUT.register\[18\]\[16\] vssd1 vssd1 vccd1 vccd1 net2014 sky130_fd_sc_hd__dlygate4sd3_1
X_09985_ net251 net2258 net623 vssd1 vssd1 vccd1 vccd1 _00190_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout584_A _01513_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08936_ net424 _04042_ _04043_ _04033_ vssd1 vssd1 vccd1 vccd1 _04044_ sky130_fd_sc_hd__a211o_1
XANTENNA__07509__B1 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08867_ net308 _03899_ _03976_ _03977_ net285 vssd1 vssd1 vccd1 vccd1 _03978_ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout372_X net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout751_A _01621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_66_clk_A clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout849_A net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07818_ top.DUT.register\[24\]\[0\] net644 net738 top.DUT.register\[12\]\[0\] _02956_
+ vssd1 vssd1 vccd1 vccd1 _02957_ sky130_fd_sc_hd__a221o_1
X_08798_ _01920_ _03893_ _01918_ vssd1 vssd1 vccd1 vccd1 _03912_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07082__A _02198_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_603 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07749_ top.DUT.register\[30\]\[3\] net581 net446 top.DUT.register\[1\]\[3\] _02887_
+ vssd1 vssd1 vccd1 vccd1 _02888_ sky130_fd_sc_hd__a221o_1
XFILLER_0_168_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout637_X net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10760_ top.DUT.register\[26\]\[0\] net145 net483 vssd1 vssd1 vccd1 vccd1 _00921_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_177_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11084__A3 net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08906__A net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09419_ net137 _04463_ _04476_ vssd1 vssd1 vccd1 vccd1 _04477_ sky130_fd_sc_hd__o21ai_1
X_10691_ top.DUT.register\[23\]\[29\] net154 net341 vssd1 vssd1 vccd1 vccd1 _00854_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10647__S net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_101_1954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_124_clk_A clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12430_ clknet_leaf_85_clk _00026_ net998 vssd1 vssd1 vccd1 vccd1 top.ramaddr\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_101_1965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_180_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_544 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09434__B1 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_173 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08788__A2 net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12361_ clknet_leaf_94_clk top.ru.next_FetchedData\[5\] net982 vssd1 vssd1 vccd1
+ vccd1 top.a1.dataIn\[5\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_145_590 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_683 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11312_ top.a1.row1\[63\] _05136_ _05197_ _05117_ vssd1 vssd1 vccd1 vccd1 _05198_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_134_2453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12292_ top.lcd.cnt_500hz\[13\] _06104_ _06106_ net687 vssd1 vssd1 vccd1 vccd1 _01348_
+ sky130_fd_sc_hd__o211a_1
XANTENNA__07460__A2 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09737__A1 _03617_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10382__S net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11243_ top.lcd.nextState\[3\] _05128_ _05135_ vssd1 vssd1 vccd1 vccd1 _05136_ sky130_fd_sc_hd__and3_4
XANTENNA__09456__B _04499_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06432__Y _01571_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07748__B1 net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_19_clk_A clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11174_ top.a1.state\[1\] top.a1.state\[0\] _05002_ _05082_ vssd1 vssd1 vccd1 vccd1
+ _05097_ sky130_fd_sc_hd__or4_1
X_10125_ net213 net1652 net607 vssd1 vssd1 vccd1 vccd1 _00325_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_180_3141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_180_3152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10056_ net1654 net232 net615 vssd1 vssd1 vccd1 vccd1 _00258_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_199_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13815_ net1100 vssd1 vssd1 vccd1 vccd1 gpio_out[2] sky130_fd_sc_hd__buf_2
XANTENNA__11226__B _05118_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_187_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08973__A2_N net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_202_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13746_ clknet_leaf_99_clk _01317_ vssd1 vssd1 vccd1 vccd1 top.lcd.cnt_20ms\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__07279__A2 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10958_ net904 _04996_ vssd1 vssd1 vccd1 vccd1 _05001_ sky130_fd_sc_hd__or2_1
XFILLER_0_128_502 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08816__A _03909_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10557__S net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13677_ clknet_leaf_90_clk _01253_ net999 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_72_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10889_ net2025 net267 net480 vssd1 vssd1 vccd1 vccd1 _01050_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_14_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12628_ clknet_leaf_56_clk _00220_ net1073 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[4\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12559_ clknet_leaf_32_clk _00151_ net1023 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[1\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07987__B1 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_182 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold106 top.ramstore\[4\] vssd1 vssd1 vccd1 vccd1 net1222 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold117 top.pad.button_control.r_counter\[14\] vssd1 vssd1 vccd1 vccd1 net1233 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08551__A net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_9_Right_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold128 top.a1.row1\[120\] vssd1 vssd1 vccd1 vccd1 net1244 sky130_fd_sc_hd__dlygate4sd3_1
Xhold139 top.ramstore\[11\] vssd1 vssd1 vccd1 vccd1 net1255 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10292__S net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_74_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_688 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout608 _04956_ vssd1 vssd1 vccd1 vccd1 net608 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08400__B2 _02830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout619 net622 vssd1 vssd1 vccd1 vccd1 net619 sky130_fd_sc_hd__buf_8
XTAP_TAPCELL_ROW_165_2914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_165_2925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_107_Right_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08951__A2 net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09770_ _04790_ _04789_ vssd1 vssd1 vccd1 vccd1 _04791_ sky130_fd_sc_hd__and2b_1
X_06982_ top.DUT.register\[4\]\[23\] net668 net739 top.DUT.register\[12\]\[23\] _02117_
+ vssd1 vssd1 vccd1 vccd1 _02121_ sky130_fd_sc_hd__a221o_1
X_08721_ net283 _03838_ vssd1 vssd1 vccd1 vccd1 _03839_ sky130_fd_sc_hd__or2_1
XFILLER_0_28_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_198_3413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08652_ _03214_ _03219_ vssd1 vssd1 vccd1 vccd1 _03773_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_105_2021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07603_ top.DUT.register\[8\]\[6\] net639 _02730_ _02741_ vssd1 vssd1 vccd1 vccd1
+ _02742_ sky130_fd_sc_hd__a211o_1
X_08583_ _02657_ _03684_ _03071_ vssd1 vssd1 vccd1 vccd1 _03707_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_44_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07534_ top.DUT.register\[22\]\[7\] net575 net551 top.DUT.register\[3\]\[7\] vssd1
+ vssd1 vccd1 vccd1 _02673_ sky130_fd_sc_hd__a22o_1
XANTENNA__07901__Y _03040_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08285__X _03421_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10975__B net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_455 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10467__S net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07465_ top.DUT.register\[13\]\[15\] net775 net767 top.DUT.register\[28\]\[15\] vssd1
+ vssd1 vccd1 vccd1 _02604_ sky130_fd_sc_hd__a22o_1
XFILLER_0_17_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1074_A net1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11152__A _04657_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09204_ _04272_ _04273_ vssd1 vssd1 vccd1 vccd1 _04274_ sky130_fd_sc_hd__nand2_1
X_06416_ net683 _01512_ _01521_ vssd1 vssd1 vccd1 vccd1 _01555_ sky130_fd_sc_hd__and3_1
XFILLER_0_119_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_173_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07690__A2 _02808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06246__A top.ramload\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07396_ top.DUT.register\[15\]\[9\] net679 net675 top.DUT.register\[31\]\[9\] vssd1
+ vssd1 vccd1 vccd1 _02535_ sky130_fd_sc_hd__a22o_1
XFILLER_0_72_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09135_ net138 _04208_ vssd1 vssd1 vccd1 vccd1 _04209_ sky130_fd_sc_hd__nor2_1
X_06347_ _01389_ _01473_ _01487_ vssd1 vssd1 vccd1 vccd1 _01489_ sky130_fd_sc_hd__and3_2
XFILLER_0_71_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07978__B1 net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09557__A _01722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09066_ _04022_ _04042_ _04093_ _04140_ vssd1 vssd1 vccd1 vccd1 _04141_ sky130_fd_sc_hd__o31a_1
X_06278_ top.lcd.cnt_500hz\[5\] top.lcd.cnt_500hz\[7\] top.lcd.cnt_500hz\[6\] top.lcd.cnt_500hz\[4\]
+ vssd1 vssd1 vccd1 vccd1 _01441_ sky130_fd_sc_hd__or4b_1
XANTENNA__07442__A2 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_116_2183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08017_ _01391_ _01392_ net893 vssd1 vssd1 vccd1 vccd1 _03156_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout799_A _04150_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold640 top.DUT.register\[27\]\[15\] vssd1 vssd1 vccd1 vccd1 net1756 sky130_fd_sc_hd__dlygate4sd3_1
Xhold651 top.DUT.register\[29\]\[2\] vssd1 vssd1 vccd1 vccd1 net1767 sky130_fd_sc_hd__dlygate4sd3_1
Xhold662 top.DUT.register\[24\]\[11\] vssd1 vssd1 vccd1 vccd1 net1778 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09991__S net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09844__X _04858_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold673 top.DUT.register\[3\]\[21\] vssd1 vssd1 vccd1 vccd1 net1789 sky130_fd_sc_hd__dlygate4sd3_1
Xhold684 top.DUT.register\[27\]\[23\] vssd1 vssd1 vccd1 vccd1 net1800 sky130_fd_sc_hd__dlygate4sd3_1
Xhold695 top.DUT.register\[6\]\[30\] vssd1 vssd1 vccd1 vccd1 net1811 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout966_A net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout587_X net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10930__S _04972_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09968_ net1743 net177 net629 vssd1 vssd1 vccd1 vccd1 _00176_ sky130_fd_sc_hd__mux2_1
XANTENNA__12856__CLK clknet_leaf_128_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07805__A _02934_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08919_ _04009_ _04027_ vssd1 vssd1 vccd1 vccd1 _04028_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout754_X net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09899_ top.pc\[28\] _04605_ vssd1 vssd1 vccd1 vccd1 _04907_ sky130_fd_sc_hd__nand2_1
X_11930_ _05774_ _05810_ _05811_ vssd1 vssd1 vccd1 vccd1 _05813_ sky130_fd_sc_hd__or3_1
XFILLER_0_197_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11861_ _05708_ _05743_ _05677_ vssd1 vssd1 vccd1 vccd1 _05744_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11046__B net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13600_ clknet_leaf_64_clk net1198 net1092 vssd1 vssd1 vccd1 vccd1 net92 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_197_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_192_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10812_ net202 net1986 net600 vssd1 vssd1 vccd1 vccd1 _00973_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_196_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11792_ _05642_ _05669_ _05670_ _05640_ vssd1 vssd1 vccd1 vccd1 _05675_ sky130_fd_sc_hd__a22o_1
XFILLER_0_67_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_45_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13531_ clknet_leaf_93_clk _01118_ net998 vssd1 vssd1 vccd1 vccd1 top.a1.data\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_10743_ net2081 net190 net419 vssd1 vssd1 vccd1 vccd1 _00904_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_165_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10377__S net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13462_ clknet_leaf_4_clk _01054_ net940 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[30\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_192_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_165_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06156__A top.a1.dataIn\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10674_ net1338 net213 net339 vssd1 vssd1 vccd1 vccd1 _00837_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_458 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07681__A2 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12413_ clknet_leaf_110_clk top.ru.next_FetchedInstr\[25\] net989 vssd1 vssd1 vccd1
+ vccd1 top.a1.instruction\[25\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_125_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_209_Right_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_211_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13393_ clknet_leaf_113_clk _00985_ net991 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[28\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_152_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07969__B1 net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07539__X _02678_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12344_ net2027 net904 net35 vssd1 vssd1 vccd1 vccd1 _01369_ sky130_fd_sc_hd__a21o_1
XANTENNA__09467__A top.pc\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07433__A2 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12275_ top.lcd.cnt_500hz\[7\] _06094_ _06095_ vssd1 vssd1 vccd1 vccd1 _01342_ sky130_fd_sc_hd__o21a_1
XANTENNA__09186__B _02778_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06162__Y _01405_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_591 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11226_ net878 _05118_ vssd1 vssd1 vccd1 vccd1 _05119_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_56_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_208_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11157_ _05085_ top.a1.row1\[56\] vssd1 vssd1 vccd1 vccd1 _05087_ sky130_fd_sc_hd__and2b_1
XANTENNA__10840__S net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_147_2644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_147_2655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10108_ top.DUT.register\[6\]\[28\] net156 net614 vssd1 vssd1 vccd1 vccd1 _00309_
+ sky130_fd_sc_hd__mux2_1
X_11088_ net908 net1291 net863 _05049_ vssd1 vssd1 vccd1 vccd1 _01195_ sky130_fd_sc_hd__a31o_1
X_10039_ net1787 net171 net619 vssd1 vssd1 vccd1 vccd1 _00242_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_160_2844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_400 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_800 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_175_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_193_3343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10287__S net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13729_ clknet_leaf_96_clk _01300_ vssd1 vssd1 vccd1 vccd1 top.a1.dataInTemp\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07250_ _02388_ vssd1 vssd1 vccd1 vccd1 _02389_ sky130_fd_sc_hd__inv_2
XANTENNA__13161__CLK clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07672__A2 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06201_ _01431_ vssd1 vssd1 vccd1 vccd1 _01432_ sky130_fd_sc_hd__inv_2
XFILLER_0_121_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06880__B1 net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07181_ top.DUT.register\[15\]\[10\] net679 net675 top.DUT.register\[31\]\[10\] vssd1
+ vssd1 vccd1 vccd1 _02320_ sky130_fd_sc_hd__a22o_1
XFILLER_0_14_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_143_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_300 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07424__A2 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08621__A1 net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_733 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06632__B1 net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08909__C1 net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout405 net406 vssd1 vssd1 vccd1 vccd1 net405 sky130_fd_sc_hd__buf_2
Xfanout427 _03259_ vssd1 vssd1 vccd1 vccd1 net427 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12181__B2 _05879_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09822_ net829 _04480_ vssd1 vssd1 vccd1 vccd1 _04838_ sky130_fd_sc_hd__nor2_1
XANTENNA__10750__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout438 _01587_ vssd1 vssd1 vccd1 vccd1 net438 sky130_fd_sc_hd__buf_2
Xfanout449 _01562_ vssd1 vssd1 vccd1 vccd1 net449 sky130_fd_sc_hd__clkbuf_8
XANTENNA__06935__B2 top.DUT.register\[11\]\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09753_ _01579_ _04172_ vssd1 vssd1 vccd1 vccd1 _04776_ sky130_fd_sc_hd__nor2_1
X_06965_ top.DUT.register\[20\]\[23\] net566 net465 top.DUT.register\[13\]\[23\] _02103_
+ vssd1 vssd1 vccd1 vccd1 _02104_ sky130_fd_sc_hd__a221o_1
X_08704_ _03732_ _03822_ net308 vssd1 vssd1 vccd1 vccd1 _03823_ sky130_fd_sc_hd__mux2_1
X_09684_ _04712_ _04718_ vssd1 vssd1 vccd1 vccd1 _04720_ sky130_fd_sc_hd__nand2_1
X_06896_ top.DUT.register\[11\]\[18\] net712 _02029_ _02031_ _02034_ vssd1 vssd1 vccd1
+ vccd1 _02035_ sky130_fd_sc_hd__a2111o_1
XANTENNA__08688__B2 _03807_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08635_ _03675_ _03756_ net310 vssd1 vssd1 vccd1 vccd1 _03757_ sky130_fd_sc_hd__mux2_1
XFILLER_0_179_744 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_92 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06699__B1 net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_87_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout547_A net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08566_ net319 _03690_ vssd1 vssd1 vccd1 vccd1 _03691_ sky130_fd_sc_hd__nor2_2
XFILLER_0_194_736 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11153__Y _05083_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07517_ _02654_ _02655_ vssd1 vssd1 vccd1 vccd1 _02656_ sky130_fd_sc_hd__and2b_1
XFILLER_0_194_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10197__S net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08497_ net316 _03427_ vssd1 vssd1 vccd1 vccd1 _03625_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout714_A _01637_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout335_X net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09986__S net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07448_ top.DUT.register\[16\]\[15\] net545 net510 top.DUT.register\[4\]\[15\] vssd1
+ vssd1 vccd1 vccd1 _02587_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_118_2212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_118_2223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06871__B1 net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_40_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10925__S net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07379_ top.DUT.register\[28\]\[8\] net766 net719 top.DUT.register\[19\]\[8\] vssd1
+ vssd1 vccd1 vccd1 _02518_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout502_X net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_160 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_631 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09118_ _04190_ _04192_ vssd1 vssd1 vccd1 vccd1 _04193_ sky130_fd_sc_hd__or2_1
XANTENNA__08612__A1 net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10390_ net1717 _04916_ net376 vssd1 vssd1 vccd1 vccd1 _00565_ sky130_fd_sc_hd__mux2_1
XANTENNA__07415__A2 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08612__B2 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_2412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06623__B1 net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09049_ _04080_ _04123_ vssd1 vssd1 vccd1 vccd1 _04124_ sky130_fd_sc_hd__nand2_1
Xclkbuf_4_4__f_clk clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_4__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_60_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12060_ _05942_ vssd1 vssd1 vccd1 vccd1 _05943_ sky130_fd_sc_hd__inv_2
Xhold470 top.DUT.register\[8\]\[7\] vssd1 vssd1 vccd1 vccd1 net1586 sky130_fd_sc_hd__dlygate4sd3_1
Xhold481 top.DUT.register\[13\]\[1\] vssd1 vssd1 vccd1 vccd1 net1597 sky130_fd_sc_hd__dlygate4sd3_1
X_11011_ wb.curr_state\[1\] net1 vssd1 vssd1 vccd1 vccd1 _05042_ sky130_fd_sc_hd__nand2_1
Xhold492 top.DUT.register\[30\]\[12\] vssd1 vssd1 vccd1 vccd1 net1608 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08915__A2 net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10660__S net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout950 net951 vssd1 vssd1 vccd1 vccd1 net950 sky130_fd_sc_hd__clkbuf_2
Xfanout961 net962 vssd1 vssd1 vccd1 vccd1 net961 sky130_fd_sc_hd__clkbuf_4
Xfanout972 net973 vssd1 vssd1 vccd1 vccd1 net972 sky130_fd_sc_hd__clkbuf_4
Xfanout983 net987 vssd1 vssd1 vccd1 vccd1 net983 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_99_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_129_2374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout994 net1000 vssd1 vssd1 vccd1 vccd1 net994 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_129_2385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12962_ clknet_leaf_11_clk _00554_ net948 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[14\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08918__X _04027_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1170 top.ramload\[10\] vssd1 vssd1 vccd1 vccd1 net2286 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_input10_A DAT_I[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11913_ _05729_ _05753_ vssd1 vssd1 vccd1 vccd1 _05796_ sky130_fd_sc_hd__xnor2_1
Xhold1181 top.ramload\[30\] vssd1 vssd1 vccd1 vccd1 net2297 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09750__A top.pc\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1192 top.ramload\[26\] vssd1 vssd1 vccd1 vccd1 net2308 sky130_fd_sc_hd__dlygate4sd3_1
X_12893_ clknet_leaf_118_clk _00485_ net954 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[12\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_206_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_142_2574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11844_ net130 _05718_ top.a1.dataIn\[6\] vssd1 vssd1 vccd1 vccd1 _05727_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_67_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07270__A _02399_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11775_ _05655_ _05656_ _05629_ vssd1 vssd1 vccd1 vccd1 _05658_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_200_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_172_408 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_175_3073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13514_ clknet_leaf_121_clk _01106_ net934 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[31\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_10726_ net1914 net148 net335 vssd1 vssd1 vccd1 vccd1 _00887_ sky130_fd_sc_hd__mux2_1
XANTENNA__07654__A2 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13445_ clknet_leaf_34_clk _01037_ net1040 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[29\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_10657_ _04916_ net2228 net345 vssd1 vssd1 vccd1 vccd1 _00821_ sky130_fd_sc_hd__mux2_1
XANTENNA__10835__S net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_119 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload15 clknet_leaf_121_clk vssd1 vssd1 vccd1 vccd1 clkload15/Y sky130_fd_sc_hd__inv_8
XANTENNA__07269__X _02408_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload26 clknet_leaf_112_clk vssd1 vssd1 vccd1 vccd1 clkload26/Y sky130_fd_sc_hd__inv_8
XFILLER_0_141_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload37 clknet_leaf_110_clk vssd1 vssd1 vccd1 vccd1 clkload37/Y sky130_fd_sc_hd__inv_8
XANTENNA__07406__A2 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13376_ clknet_leaf_17_clk _00968_ net965 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[27\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_58_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10588_ net1349 net170 net350 vssd1 vssd1 vccd1 vccd1 _00754_ sky130_fd_sc_hd__mux2_1
Xclkload48 clknet_leaf_86_clk vssd1 vssd1 vccd1 vccd1 clkload48/Y sky130_fd_sc_hd__inv_8
XFILLER_0_50_152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload59 clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 clkload59/Y sky130_fd_sc_hd__inv_6
X_12327_ _06127_ _06128_ vssd1 vssd1 vccd1 vccd1 _01361_ sky130_fd_sc_hd__nor2_1
XANTENNA__06614__B1 net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08958__A1_N _02652_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_39_Left_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07429__B _02567_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_192_Right_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12258_ net979 net815 _06059_ vssd1 vssd1 vccd1 vccd1 _06086_ sky130_fd_sc_hd__and3_1
XFILLER_0_121_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11209_ net845 _05099_ vssd1 vssd1 vccd1 vccd1 _05111_ sky130_fd_sc_hd__and2_1
XANTENNA__10570__S net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12189_ top.a1.row2\[15\] net851 _05083_ vssd1 vssd1 vccd1 vccd1 _01297_ sky130_fd_sc_hd__o21a_1
XFILLER_0_207_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06750_ top.DUT.register\[23\]\[24\] net574 _01888_ vssd1 vssd1 vccd1 vccd1 _01889_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_210_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06681_ top.DUT.register\[30\]\[26\] net761 net642 top.DUT.register\[8\]\[26\] _01813_
+ vssd1 vssd1 vccd1 vccd1 _01820_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_48_Left_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_203_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_69_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08420_ _03231_ _03251_ vssd1 vssd1 vccd1 vccd1 _03551_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_69_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07451__Y _02590_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07893__A2 net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08276__A net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08351_ net429 _03473_ _03484_ vssd1 vssd1 vccd1 vccd1 _03485_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_86_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07302_ top.DUT.register\[23\]\[12\] net572 net564 top.DUT.register\[20\]\[12\] vssd1
+ vssd1 vccd1 vccd1 _02441_ sky130_fd_sc_hd__a22o_1
XFILLER_0_128_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08282_ _02995_ net287 _03288_ vssd1 vssd1 vccd1 vccd1 _03418_ sky130_fd_sc_hd__or3_1
XFILLER_0_18_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07645__A2 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_156_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload9 clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 clkload9/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_143_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07233_ top.DUT.register\[9\]\[10\] net762 net706 top.DUT.register\[15\]\[10\] vssd1
+ vssd1 vccd1 vccd1 _02372_ sky130_fd_sc_hd__a22o_1
XANTENNA__10745__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09819__B _04487_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07164_ top.DUT.register\[29\]\[11\] net722 _02296_ _02298_ _02302_ vssd1 vssd1 vccd1
+ vccd1 _02303_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_144_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07095_ top.DUT.register\[2\]\[16\] net560 _02233_ vssd1 vssd1 vccd1 vccd1 _02234_
+ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_113_2142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06243__B net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1037_A net1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09394__X _04453_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12377__RESET_B net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout202 _04841_ vssd1 vssd1 vccd1 vccd1 net202 sky130_fd_sc_hd__buf_2
XANTENNA_fanout497_A net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13057__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout213 net214 vssd1 vssd1 vccd1 vccd1 net213 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__10480__S net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout224 _04805_ vssd1 vssd1 vccd1 vccd1 net224 sky130_fd_sc_hd__buf_1
Xfanout235 _04757_ vssd1 vssd1 vccd1 vccd1 net235 sky130_fd_sc_hd__buf_2
Xfanout246 _04749_ vssd1 vssd1 vccd1 vccd1 net246 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_208_3559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout257 net258 vssd1 vssd1 vccd1 vccd1 net257 sky130_fd_sc_hd__clkbuf_2
XANTENNA_input2_A DAT_I[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09805_ _03787_ net404 net489 _04822_ vssd1 vssd1 vccd1 vccd1 _04823_ sky130_fd_sc_hd__o211a_1
Xfanout268 _04726_ vssd1 vssd1 vccd1 vccd1 net268 sky130_fd_sc_hd__buf_1
Xfanout279 _03239_ vssd1 vssd1 vccd1 vccd1 net279 sky130_fd_sc_hd__clkbuf_4
X_07997_ top.DUT.register\[25\]\[31\] net780 net752 top.DUT.register\[26\]\[31\] vssd1
+ vssd1 vccd1 vccd1 _03136_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout285_X net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout664_A _01605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06948_ _02080_ _02082_ _02084_ _02086_ vssd1 vssd1 vccd1 vccd1 _02087_ sky130_fd_sc_hd__or4_1
X_09736_ top.pc\[10\] net799 _04754_ _04761_ vssd1 vssd1 vccd1 vccd1 _04762_ sky130_fd_sc_hd__a211o_1
Xclkbuf_4_12__f_clk clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_12__leaf_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_179_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09667_ _04191_ _04193_ vssd1 vssd1 vccd1 vccd1 _04704_ sky130_fd_sc_hd__and2_1
X_06879_ top.DUT.register\[19\]\[18\] net537 net509 top.DUT.register\[4\]\[18\] vssd1
+ vssd1 vccd1 vccd1 _02018_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_2_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout452_X net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout831_A net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08618_ _02265_ _03185_ net492 _02266_ _03740_ vssd1 vssd1 vccd1 vccd1 _03741_ sky130_fd_sc_hd__o221a_1
XFILLER_0_139_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_179_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12200__S _06049_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09598_ top.a1.instruction\[31\] net822 net422 vssd1 vssd1 vccd1 vccd1 _04644_ sky130_fd_sc_hd__a21o_2
XANTENNA__07884__A2 net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08549_ _03627_ _03674_ net289 vssd1 vssd1 vccd1 vccd1 _03675_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_403 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout717_X net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07097__B1 net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11560_ _05431_ _05440_ _05442_ vssd1 vssd1 vccd1 vccd1 _05443_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_119_151 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08833__B2 net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_255 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_406 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10511_ net2042 net190 net358 vssd1 vssd1 vccd1 vccd1 _00680_ sky130_fd_sc_hd__mux2_1
XANTENNA__10655__S net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11491_ _05366_ _05373_ vssd1 vssd1 vccd1 vccd1 _05374_ sky130_fd_sc_hd__nor2_1
XFILLER_0_17_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_21_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13230_ clknet_leaf_41_clk _00822_ net1057 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[22\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_10442_ net211 net2078 net365 vssd1 vssd1 vccd1 vccd1 _00613_ sky130_fd_sc_hd__mux2_1
X_13161_ clknet_leaf_50_clk _00753_ net1058 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[20\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_10373_ net1511 net221 net373 vssd1 vssd1 vccd1 vccd1 _00548_ sky130_fd_sc_hd__mux2_1
X_12112_ _05994_ vssd1 vssd1 vccd1 vccd1 _05995_ sky130_fd_sc_hd__inv_2
X_13092_ clknet_leaf_36_clk _00684_ net1049 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[18\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10390__S net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12043_ _05913_ _05919_ _05922_ _05925_ vssd1 vssd1 vccd1 vccd1 _05926_ sky130_fd_sc_hd__a31oi_1
XTAP_TAPCELL_ROW_53_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07021__B1 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_144_2603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout780 _01603_ vssd1 vssd1 vccd1 vccd1 net780 sky130_fd_sc_hd__clkbuf_8
Xfanout791 _06112_ vssd1 vssd1 vccd1 vccd1 net791 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_189_316 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09313__A2 top.pc\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12945_ clknet_leaf_121_clk _00537_ net977 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[14\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_177_3102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08808__B net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07712__B _02849_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12876_ clknet_leaf_63_clk _00468_ net1091 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[11\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07875__A2 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_158_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11827_ _05708_ _05709_ vssd1 vssd1 vccd1 vccd1 _05710_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_190_3302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07088__B1 net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11758_ _05595_ _05622_ vssd1 vssd1 vccd1 vccd1 _05641_ sky130_fd_sc_hd__xor2_4
XANTENNA__07627__A2 net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06835__B1 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10709_ net1802 net208 net335 vssd1 vssd1 vccd1 vccd1 _00870_ sky130_fd_sc_hd__mux2_1
XANTENNA__10565__S net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_155_2765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11689_ _05537_ _05570_ vssd1 vssd1 vccd1 vccd1 _05572_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_70_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload104 clknet_leaf_61_clk vssd1 vssd1 vccd1 vccd1 clkload104/Y sky130_fd_sc_hd__inv_8
XTAP_TAPCELL_ROW_155_2776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_181_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_66 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13428_ clknet_leaf_79_clk _01020_ net1073 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[29\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_178_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11187__A2 net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08588__B1 net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13359_ clknet_leaf_22_clk _00951_ net1056 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[26\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_178_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_188_3264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_68 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12470__RESET_B net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07920_ _02659_ _03057_ vssd1 vssd1 vccd1 vccd1 _03059_ sky130_fd_sc_hd__or2_1
XANTENNA__11229__A_N top.lcd.nextState\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07012__B1 net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07851_ top.DUT.register\[14\]\[0\] net584 net443 top.DUT.register\[1\]\[0\] _02989_
+ vssd1 vssd1 vccd1 vccd1 _02990_ sky130_fd_sc_hd__a221o_1
X_06802_ top.DUT.register\[15\]\[17\] net707 net699 top.DUT.register\[31\]\[17\] vssd1
+ vssd1 vccd1 vccd1 _01941_ sky130_fd_sc_hd__a22o_1
X_07782_ top.DUT.register\[20\]\[2\] net663 net647 top.DUT.register\[22\]\[2\] _02920_
+ vssd1 vssd1 vccd1 vccd1 _02921_ sky130_fd_sc_hd__a221o_1
Xinput2 DAT_I[0] vssd1 vssd1 vccd1 vccd1 net2 sky130_fd_sc_hd__clkbuf_1
X_09521_ top.pc\[26\] _04560_ vssd1 vssd1 vccd1 vccd1 _04572_ sky130_fd_sc_hd__and2_1
X_06733_ top.DUT.register\[26\]\[25\] net751 _01857_ _01862_ _01871_ vssd1 vssd1 vccd1
+ vccd1 _01872_ sky130_fd_sc_hd__a2111oi_1
XANTENNA__07903__A net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_203_3489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09452_ top.pc\[21\] _04478_ top.pc\[22\] vssd1 vssd1 vccd1 vccd1 _04507_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_149_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_210_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06664_ top.DUT.register\[13\]\[26\] net464 net544 top.DUT.register\[16\]\[26\] _01802_
+ vssd1 vssd1 vccd1 vccd1 _01803_ sky130_fd_sc_hd__a221o_1
XANTENNA__07866__A2 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06519__A _01571_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08403_ net324 net333 vssd1 vssd1 vccd1 vccd1 _03535_ sky130_fd_sc_hd__nor2_2
X_09383_ _04436_ _04440_ _04441_ _04442_ net811 vssd1 vssd1 vccd1 vccd1 _04443_ sky130_fd_sc_hd__a311o_1
XFILLER_0_149_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06595_ top.DUT.register\[7\]\[28\] net661 net658 top.DUT.register\[21\]\[28\] _01727_
+ vssd1 vssd1 vccd1 vccd1 _01734_ sky130_fd_sc_hd__a221o_1
XFILLER_0_93_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08334_ net302 _03306_ _03467_ vssd1 vssd1 vccd1 vccd1 _03468_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07618__A2 net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08815__A1 net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06826__B1 net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08265_ _03398_ _03400_ net312 vssd1 vssd1 vccd1 vccd1 _03401_ sky130_fd_sc_hd__mux2_1
XANTENNA__10475__S net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07216_ _02350_ _02352_ _02354_ _02349_ vssd1 vssd1 vccd1 vccd1 _02355_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_104_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_794 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08196_ _03164_ _03182_ vssd1 vssd1 vccd1 vccd1 _03334_ sky130_fd_sc_hd__nor2_4
XFILLER_0_14_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07147_ _02276_ _02285_ vssd1 vssd1 vccd1 vccd1 _02286_ sky130_fd_sc_hd__nor2_8
XFILLER_0_15_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09240__A1 net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09240__B2 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_1867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_1878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07078_ _02213_ _02214_ _02215_ _02216_ vssd1 vssd1 vccd1 vccd1 _02217_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout781_A _01603_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout879_A top.lcd.nextState\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1008 net1016 vssd1 vssd1 vccd1 vccd1 net1008 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_7_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1019 net1020 vssd1 vssd1 vccd1 vccd1 net1019 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07003__B1 net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11319__B net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout667_X net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_303 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09719_ net407 _04747_ vssd1 vssd1 vccd1 vccd1 _04748_ sky130_fd_sc_hd__or2_1
X_10991_ top.a1.data\[3\] net783 vssd1 vssd1 vccd1 vccd1 _05027_ sky130_fd_sc_hd__or2_1
XFILLER_0_198_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12730_ clknet_leaf_0_clk _00322_ net916 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[7\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_26_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12661_ clknet_leaf_31_clk _00253_ net1020 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[5\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_194_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11612_ _05465_ _05481_ vssd1 vssd1 vccd1 vccd1 _05495_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_77_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08806__A1 net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_172_3021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12592_ clknet_leaf_28_clk _00184_ net1010 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[2\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_172_3032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11543_ _05372_ _05412_ vssd1 vssd1 vccd1 vccd1 _05426_ sky130_fd_sc_hd__xnor2_2
XANTENNA__06817__B1 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10385__S net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_761 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11474_ _05349_ _05354_ _05355_ _05356_ vssd1 vssd1 vccd1 vccd1 _05357_ sky130_fd_sc_hd__a211o_1
XANTENNA__07490__B1 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_2495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13213_ clknet_leaf_119_clk _00805_ net930 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[22\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_10425_ net1320 net157 net370 vssd1 vssd1 vccd1 vccd1 _00597_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07242__B1 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13144_ clknet_leaf_128_clk _00736_ net921 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[20\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09475__A _01585_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10356_ net1993 net160 net378 vssd1 vssd1 vccd1 vccd1 _00532_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_150_2695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06596__A2 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13075_ clknet_leaf_120_clk _00667_ net932 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[18\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_10287_ net1713 net175 net387 vssd1 vssd1 vccd1 vccd1 _00465_ sky130_fd_sc_hd__mux2_1
X_12026_ top.a1.dataIn\[4\] _05879_ vssd1 vssd1 vccd1 vccd1 _05909_ sky130_fd_sc_hd__xnor2_2
XTAP_TAPCELL_ROW_183_3194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09883__B1_N _04892_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_66_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12928_ clknet_leaf_79_clk _00520_ net1073 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[13\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07848__A2 net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10852__A1 net156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_157_2805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12859_ clknet_leaf_124_clk _00451_ net923 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[11\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_374 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06380_ net684 _01516_ _01518_ vssd1 vssd1 vccd1 vccd1 _01519_ sky130_fd_sc_hd__and3_4
XFILLER_0_90_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06808__B1 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08050_ _01722_ net328 vssd1 vssd1 vccd1 vccd1 _03189_ sky130_fd_sc_hd__or2_1
XANTENNA__06284__A1 top.lcd.nextState\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07481__B1 net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07001_ top.DUT.register\[13\]\[20\] net464 net505 top.DUT.register\[27\]\[20\] _02139_
+ vssd1 vssd1 vccd1 vccd1 _02140_ sky130_fd_sc_hd__a221o_1
XFILLER_0_153_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_141_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07233__B1 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_2101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06587__A2 net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08952_ _02521_ _04050_ net1292 net877 vssd1 vssd1 vccd1 vccd1 _00058_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_168_2967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09672__X _04708_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07903_ net295 _03040_ vssd1 vssd1 vccd1 vccd1 _03042_ sky130_fd_sc_hd__nand2_1
XFILLER_0_209_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08883_ _01702_ _03992_ vssd1 vssd1 vccd1 vccd1 _03993_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_205_3518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout195_A _04850_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07834_ net408 vssd1 vssd1 vccd1 vccd1 _02973_ sky130_fd_sc_hd__inv_2
X_07765_ net805 _01582_ _02903_ vssd1 vssd1 vccd1 vccd1 _02904_ sky130_fd_sc_hd__a21o_2
XTAP_TAPCELL_ROW_108_2063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout362_A net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06716_ top.DUT.register\[4\]\[25\] net667 net664 top.DUT.register\[20\]\[25\] vssd1
+ vssd1 vccd1 vccd1 _01855_ sky130_fd_sc_hd__a22o_1
XANTENNA__11096__A1 net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09504_ top.pc\[24\] top.pc\[25\] _04521_ vssd1 vssd1 vccd1 vccd1 _04556_ sky130_fd_sc_hd__and3_1
XFILLER_0_79_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_189_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_177_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07839__A2 net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07696_ top.DUT.register\[30\]\[4\] net581 net520 top.DUT.register\[10\]\[4\] vssd1
+ vssd1 vccd1 vccd1 _02835_ sky130_fd_sc_hd__a22o_1
XFILLER_0_195_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09435_ net133 _04486_ _04490_ _04491_ net901 vssd1 vssd1 vccd1 vccd1 _04492_ sky130_fd_sc_hd__o221ai_1
XFILLER_0_149_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06647_ _01764_ _01784_ vssd1 vssd1 vccd1 vccd1 _01786_ sky130_fd_sc_hd__and2_1
XFILLER_0_78_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_121_2263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_339 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06511__A2 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout627_A _04948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_176_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_164_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09366_ net137 _04412_ _04426_ vssd1 vssd1 vccd1 vccd1 _04427_ sky130_fd_sc_hd__o21ai_1
X_06578_ top.DUT.register\[23\]\[28\] net573 net509 top.DUT.register\[4\]\[28\] _01716_
+ vssd1 vssd1 vccd1 vccd1 _01717_ sky130_fd_sc_hd__a221o_1
XANTENNA__12739__RESET_B net1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08317_ _03451_ vssd1 vssd1 vccd1 vccd1 _03452_ sky130_fd_sc_hd__inv_2
XFILLER_0_117_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09297_ top.pc\[12\] _04326_ top.pc\[13\] vssd1 vssd1 vccd1 vccd1 _04361_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_97_1907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_772 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09994__S net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08248_ _02947_ _03384_ vssd1 vssd1 vccd1 vccd1 _03385_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_62_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_160_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08179_ _01854_ net329 vssd1 vssd1 vccd1 vccd1 _03317_ sky130_fd_sc_hd__or2_1
XANTENNA__10933__S net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10210_ net207 net1553 net394 vssd1 vssd1 vccd1 vccd1 _00390_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_37_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11190_ top.a1.dataInTemp\[10\] top.a1.data\[10\] net785 vssd1 vssd1 vccd1 vccd1
+ _05102_ sky130_fd_sc_hd__mux2_1
XFILLER_0_113_680 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06578__A2 net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10141_ net157 net2188 net610 vssd1 vssd1 vccd1 vccd1 _00341_ sky130_fd_sc_hd__mux2_1
XANTENNA__11308__C1 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_50_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10072_ net1380 net171 net615 vssd1 vssd1 vccd1 vccd1 _00274_ sky130_fd_sc_hd__mux2_1
XANTENNA__09921__C1 _04927_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13831_ net1115 vssd1 vssd1 vccd1 vccd1 gpio_out[30] sky130_fd_sc_hd__buf_2
XFILLER_0_202_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06750__A2 net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10974_ net1165 _05014_ net589 vssd1 vssd1 vccd1 vccd1 _01116_ sky130_fd_sc_hd__mux2_1
X_13762_ clknet_leaf_70_clk _01333_ vssd1 vssd1 vccd1 vccd1 top.lcd.currentState\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__06159__A top.a1.dataIn\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_186_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12713_ clknet_leaf_50_clk _00305_ net1058 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[6\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_48_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_648 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13693_ clknet_leaf_73_clk _01264_ vssd1 vssd1 vccd1 vccd1 net122 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_84_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06502__A2 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_194_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_139_2524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12644_ clknet_leaf_36_clk _00236_ net1050 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[4\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_139_2535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_61_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12575_ clknet_leaf_20_clk _00167_ net1028 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[2\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08255__A2 top.pc\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09757__X _04780_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11526_ _05402_ _05408_ vssd1 vssd1 vccd1 vccd1 _05409_ sky130_fd_sc_hd__nor2_1
XANTENNA__07463__B1 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_152_2724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10843__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11457_ _05339_ vssd1 vssd1 vccd1 vccd1 _05340_ sky130_fd_sc_hd__inv_2
XANTENNA__12762__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10408_ net2125 net222 net369 vssd1 vssd1 vccd1 vccd1 _00580_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_185_3223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11388_ _05239_ _05270_ vssd1 vssd1 vccd1 vccd1 _05271_ sky130_fd_sc_hd__and2_1
XANTENNA__06569__A2 net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10339_ net1941 net227 net377 vssd1 vssd1 vccd1 vccd1 _00515_ sky130_fd_sc_hd__mux2_1
X_13127_ clknet_leaf_6_clk _00719_ net937 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[19\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_13058_ clknet_leaf_25_clk _00650_ net1012 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[17\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_12009_ _05890_ _05891_ vssd1 vssd1 vccd1 vccd1 _05892_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_163_2886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_191_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_163_2897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13268__CLK clknet_4_12__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06741__A2 net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07550_ top.DUT.register\[23\]\[7\] net671 net718 top.DUT.register\[19\]\[7\] vssd1
+ vssd1 vccd1 vccd1 _02689_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_200_3448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06501_ net787 _01596_ _01607_ vssd1 vssd1 vccd1 vccd1 _01640_ sky130_fd_sc_hd__and3_4
XFILLER_0_88_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_186_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07481_ top.DUT.register\[3\]\[14\] net553 net548 top.DUT.register\[18\]\[14\] _02619_
+ vssd1 vssd1 vccd1 vccd1 _02620_ sky130_fd_sc_hd__a221o_1
XFILLER_0_75_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09691__A1 _03353_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_196_3385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09220_ top.pc\[8\] _02682_ vssd1 vssd1 vccd1 vccd1 _04289_ sky130_fd_sc_hd__nor2_1
XFILLER_0_173_300 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06432_ _01545_ _01570_ vssd1 vssd1 vccd1 vccd1 _01571_ sky130_fd_sc_hd__nor2_2
XANTENNA__11703__A top.a1.dataIn\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12832__RESET_B net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_238 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09151_ net138 _04223_ vssd1 vssd1 vccd1 vccd1 _04224_ sky130_fd_sc_hd__nor2_1
X_06363_ top.a1.instruction\[0\] top.a1.instruction\[1\] top.a1.instruction\[2\] vssd1
+ vssd1 vccd1 vccd1 _01502_ sky130_fd_sc_hd__and3_1
XANTENNA__08246__A2 net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08102_ _02590_ net328 vssd1 vssd1 vccd1 vccd1 _03241_ sky130_fd_sc_hd__nand2_1
XFILLER_0_173_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09082_ top.a1.instruction\[6\] top.a1.instruction\[11\] top.a1.instruction\[19\]
+ top.a1.instruction\[21\] vssd1 vssd1 vccd1 vccd1 _04157_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_79_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07454__B1 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06294_ _01331_ _01451_ vssd1 vssd1 vccd1 vccd1 _01452_ sky130_fd_sc_hd__nor2_1
X_08033_ net301 _02994_ vssd1 vssd1 vccd1 vccd1 _03172_ sky130_fd_sc_hd__nand2_2
XFILLER_0_4_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_140_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10753__S net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold800 top.DUT.register\[25\]\[4\] vssd1 vssd1 vccd1 vccd1 net1916 sky130_fd_sc_hd__dlygate4sd3_1
Xhold811 top.DUT.register\[7\]\[18\] vssd1 vssd1 vccd1 vccd1 net1927 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_431 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold822 top.DUT.register\[23\]\[16\] vssd1 vssd1 vccd1 vccd1 net1938 sky130_fd_sc_hd__dlygate4sd3_1
Xhold833 top.DUT.register\[5\]\[24\] vssd1 vssd1 vccd1 vccd1 net1949 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09746__A2 _04752_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_1826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold844 top.DUT.register\[5\]\[3\] vssd1 vssd1 vccd1 vccd1 net1960 sky130_fd_sc_hd__dlygate4sd3_1
Xhold855 top.DUT.register\[24\]\[25\] vssd1 vssd1 vccd1 vccd1 net1971 sky130_fd_sc_hd__dlygate4sd3_1
Xhold866 top.DUT.register\[17\]\[27\] vssd1 vssd1 vccd1 vccd1 net1982 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08954__B1 _02383_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold877 top.DUT.register\[13\]\[27\] vssd1 vssd1 vccd1 vccd1 net1993 sky130_fd_sc_hd__dlygate4sd3_1
Xhold888 top.DUT.register\[24\]\[0\] vssd1 vssd1 vccd1 vccd1 net2004 sky130_fd_sc_hd__dlygate4sd3_1
Xhold899 top.DUT.register\[22\]\[29\] vssd1 vssd1 vccd1 vccd1 net2015 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06251__B net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09984_ net255 net2099 net625 vssd1 vssd1 vccd1 vccd1 _00189_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08935_ net436 _04038_ _04040_ _03144_ vssd1 vssd1 vccd1 vccd1 _04043_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout577_A net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08706__B1 net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06980__A2 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07634__Y _02773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_707 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08866_ net289 _03189_ _03197_ net306 vssd1 vssd1 vccd1 vccd1 _03977_ sky130_fd_sc_hd__a31o_1
X_07817_ top.DUT.register\[21\]\[0\] net655 _02954_ _02955_ vssd1 vssd1 vccd1 vccd1
+ _02956_ sky130_fd_sc_hd__a211o_1
XANTENNA__06193__B1 net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08797_ net1732 net830 net800 _03911_ vssd1 vssd1 vccd1 vccd1 _00042_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout365_X net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout744_A _01623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09989__S net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07748_ top.DUT.register\[22\]\[3\] net576 net528 top.DUT.register\[26\]\[3\] vssd1
+ vssd1 vccd1 vccd1 _02887_ sky130_fd_sc_hd__a22o_1
XANTENNA__11316__C _01442_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12635__CLK clknet_leaf_120_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07679_ top.DUT.register\[22\]\[4\] net649 net716 top.DUT.register\[27\]\[4\] vssd1
+ vssd1 vccd1 vccd1 _02818_ sky130_fd_sc_hd__a22o_1
XANTENNA__10928__S net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout532_X net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09682__A1 top.a1.instruction\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09418_ net133 _04468_ _04475_ net811 net901 vssd1 vssd1 vccd1 vccd1 _04476_ sky130_fd_sc_hd__o221a_1
XFILLER_0_192_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10690_ net1715 net158 net341 vssd1 vssd1 vccd1 vccd1 _00853_ sky130_fd_sc_hd__mux2_1
XANTENNA__07693__B1 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_176_182 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_4_3__f_clk_A clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_1955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_101_1966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12502__RESET_B net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09349_ top.pc\[15\] top.pc\[16\] _04377_ vssd1 vssd1 vccd1 vccd1 _04410_ sky130_fd_sc_hd__and3_1
XFILLER_0_180_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_43_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_191_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12360_ clknet_leaf_95_clk top.ru.next_FetchedData\[4\] net981 vssd1 vssd1 vccd1
+ vccd1 top.a1.dataIn\[4\] sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_43_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07445__B1 net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06799__A2 net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11311_ top.a1.row2\[15\] _05135_ top.lcd.nextState\[5\] vssd1 vssd1 vccd1 vccd1
+ _05197_ sky130_fd_sc_hd__or3b_1
XFILLER_0_90_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_134_2454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13779__RESET_B net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12291_ _06105_ vssd1 vssd1 vccd1 vccd1 _06106_ sky130_fd_sc_hd__inv_2
XANTENNA__10663__S net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11242_ net879 _05131_ vssd1 vssd1 vccd1 vccd1 _05135_ sky130_fd_sc_hd__nor2_1
XANTENNA__09737__A2 net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11173_ top.a1.row1\[63\] _05085_ _05096_ net851 vssd1 vssd1 vccd1 vccd1 _01233_
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_38_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10124_ net220 net1946 net607 vssd1 vssd1 vccd1 vccd1 _00324_ sky130_fd_sc_hd__mux2_1
XANTENNA__13361__RESET_B net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_180_3142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10055_ net1542 net238 net616 vssd1 vssd1 vccd1 vccd1 _00257_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_180_3153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08369__A _03230_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06723__A2 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_740 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13814_ net1099 vssd1 vssd1 vccd1 vccd1 gpio_out[1] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_11_Left_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_187_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13745_ clknet_leaf_99_clk _01316_ vssd1 vssd1 vccd1 vccd1 top.lcd.cnt_20ms\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_10957_ _04657_ _04998_ vssd1 vssd1 vccd1 vccd1 _05000_ sky130_fd_sc_hd__or2_1
XANTENNA__10838__S net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08816__B _03929_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_195_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07684__B1 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_49 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13676_ clknet_leaf_90_clk _01252_ net999 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_10888_ net1862 net144 net479 vssd1 vssd1 vccd1 vccd1 _01049_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_14_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12627_ clknet_leaf_123_clk _00219_ net927 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[4\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_66_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07436__B1 net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12558_ clknet_leaf_39_clk _00150_ net1054 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[1\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_11509_ _05388_ _05389_ vssd1 vssd1 vccd1 vccd1 _05392_ sky130_fd_sc_hd__xor2_2
XPHY_EDGE_ROW_20_Left_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10573__S net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold107 _01164_ vssd1 vssd1 vccd1 vccd1 net1223 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12489_ clknet_leaf_74_clk top.a1.nextHex\[7\] net1077 vssd1 vssd1 vccd1 vccd1 top.a1.hexop\[3\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold118 top.a1.row1\[10\] vssd1 vssd1 vccd1 vccd1 net1234 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09189__B1 net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold129 top.ramload\[6\] vssd1 vssd1 vccd1 vccd1 net1245 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13449__RESET_B net1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09728__A2 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10145__Y _04957_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_186_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout609 _04956_ vssd1 vssd1 vccd1 vccd1 net609 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_95_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_165_2915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_165_2926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06981_ top.DUT.register\[28\]\[23\] net767 net760 top.DUT.register\[30\]\[23\] _02119_
+ vssd1 vssd1 vccd1 vccd1 _02120_ sky130_fd_sc_hd__a221o_1
XANTENNA_clkbuf_4_14__f_clk_A clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11257__X _05150_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08720_ _03756_ _03837_ net310 vssd1 vssd1 vccd1 vccd1 _03838_ sky130_fd_sc_hd__mux2_1
XANTENNA__08279__A _03187_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08651_ net322 _03373_ vssd1 vssd1 vccd1 vccd1 _03772_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_198_3414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07911__A1 _02880_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07602_ top.DUT.register\[23\]\[6\] net671 net746 top.DUT.register\[17\]\[6\] _02731_
+ vssd1 vssd1 vccd1 vccd1 _02741_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_105_2022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08582_ net2311 net832 net802 _03706_ vssd1 vssd1 vccd1 vccd1 _00032_ sky130_fd_sc_hd__a22o_1
XFILLER_0_49_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07470__X _02609_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07533_ top.DUT.register\[21\]\[7\] net447 net507 top.DUT.register\[4\]\[7\] _02671_
+ vssd1 vssd1 vccd1 vccd1 _02672_ sky130_fd_sc_hd__a221o_1
XFILLER_0_44_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10748__S net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09664__A1 top.a1.halfData\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout158_A _04916_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07464_ top.DUT.register\[29\]\[15\] net723 _02591_ _02602_ vssd1 vssd1 vccd1 vccd1
+ _02603_ sky130_fd_sc_hd__a211o_1
XANTENNA__07675__B1 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_33_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06415_ net683 _01518_ _01521_ vssd1 vssd1 vccd1 vccd1 _01554_ sky130_fd_sc_hd__and3_4
X_09203_ _04254_ _04255_ _04257_ vssd1 vssd1 vccd1 vccd1 _04273_ sky130_fd_sc_hd__a21o_1
XANTENNA__11152__B net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07395_ _02527_ _02529_ _02531_ _02533_ vssd1 vssd1 vccd1 vccd1 _02534_ sky130_fd_sc_hd__or4_2
XANTENNA_fanout325_A net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06246__B net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09134_ top.pc\[2\] top.pc\[3\] vssd1 vssd1 vccd1 vccd1 _04208_ sky130_fd_sc_hd__xnor2_1
X_06346_ top.a1.instruction\[4\] _01484_ vssd1 vssd1 vccd1 vccd1 _01488_ sky130_fd_sc_hd__or2_1
XFILLER_0_115_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09065_ _03444_ _04134_ _04139_ _04119_ _04129_ vssd1 vssd1 vccd1 vccd1 _04140_ sky130_fd_sc_hd__o311a_1
XANTENNA__10483__S net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06277_ top.lcd.cnt_500hz\[8\] _01404_ top.lcd.cnt_500hz\[13\] top.lcd.cnt_500hz\[12\]
+ vssd1 vssd1 vccd1 vccd1 _01440_ sky130_fd_sc_hd__or4_1
XANTENNA__09557__B _04605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_194 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_403 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08016_ _03149_ _03148_ vssd1 vssd1 vccd1 vccd1 _03155_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_116_2184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold630 top.DUT.register\[31\]\[6\] vssd1 vssd1 vccd1 vccd1 net1746 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06262__A top.ramload\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout694_A net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold641 top.DUT.register\[25\]\[13\] vssd1 vssd1 vccd1 vccd1 net1757 sky130_fd_sc_hd__dlygate4sd3_1
Xhold652 top.DUT.register\[9\]\[16\] vssd1 vssd1 vccd1 vccd1 net1768 sky130_fd_sc_hd__dlygate4sd3_1
Xhold663 top.DUT.register\[16\]\[0\] vssd1 vssd1 vccd1 vccd1 net1779 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold674 top.DUT.register\[27\]\[29\] vssd1 vssd1 vccd1 vccd1 net1790 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold685 top.DUT.register\[5\]\[17\] vssd1 vssd1 vccd1 vccd1 net1801 sky130_fd_sc_hd__dlygate4sd3_1
Xhold696 top.DUT.register\[9\]\[25\] vssd1 vssd1 vccd1 vccd1 net1812 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09573__A _01678_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09967_ net2194 net182 net628 vssd1 vssd1 vccd1 vccd1 _00175_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout861_A net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout482_X net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08918_ _01657_ net502 _04026_ vssd1 vssd1 vccd1 vccd1 _04027_ sky130_fd_sc_hd__a21o_1
XANTENNA__07805__B _02943_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09898_ net2163 net161 net634 vssd1 vssd1 vccd1 vccd1 _00148_ sky130_fd_sc_hd__mux2_1
XFILLER_0_197_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08849_ _01788_ net501 _03185_ _01786_ vssd1 vssd1 vccd1 vccd1 _03961_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_99_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06705__A2 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12500__Q top.pc\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout747_X net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11860_ _05716_ _05718_ _05705_ _05707_ _05710_ vssd1 vssd1 vccd1 vccd1 _05743_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_86_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_196_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10811_ net184 net2094 net600 vssd1 vssd1 vccd1 vccd1 _00972_ sky130_fd_sc_hd__mux2_1
XFILLER_0_169_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10658__S net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11791_ _05642_ _05669_ _05670_ _05640_ vssd1 vssd1 vccd1 vccd1 _05674_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_184_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_45_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13530_ clknet_leaf_92_clk _01117_ net998 vssd1 vssd1 vccd1 vccd1 top.a1.data\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_10742_ net1371 net198 net419 vssd1 vssd1 vccd1 vccd1 _00903_ sky130_fd_sc_hd__mux2_1
XANTENNA__07130__A2 net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_165_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13461_ clknet_leaf_34_clk _01053_ net1040 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[30\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_10673_ net2273 net219 net338 vssd1 vssd1 vccd1 vccd1 _00836_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_11_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_173_Right_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_165_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12412_ clknet_leaf_108_clk top.ru.next_FetchedInstr\[24\] net975 vssd1 vssd1 vccd1
+ vccd1 top.a1.instruction\[24\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__07418__B1 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13392_ clknet_leaf_28_clk _00984_ net1011 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[27\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_12343_ net1123 _06137_ net791 vssd1 vssd1 vccd1 vccd1 _01368_ sky130_fd_sc_hd__o21a_1
XANTENNA__10393__S net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_572 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12274_ top.lcd.cnt_500hz\[7\] _06094_ net686 vssd1 vssd1 vccd1 vccd1 _06095_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_105_296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06172__A top.a1.halfData\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11225_ top.lcd.nextState\[5\] _05117_ vssd1 vssd1 vccd1 vccd1 _05118_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_56_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12190__A2 net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09483__A net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11156_ top.a1.halfData\[5\] net888 _01415_ _01418_ _01377_ vssd1 vssd1 vccd1 vccd1
+ _05086_ sky130_fd_sc_hd__o32a_1
XANTENNA__06944__A2 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_207_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10107_ net2248 net161 net613 vssd1 vssd1 vccd1 vccd1 _00308_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_147_2645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_147_2656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11087_ net65 net867 vssd1 vssd1 vccd1 vccd1 _05049_ sky130_fd_sc_hd__and2_1
XANTENNA__08099__A net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10038_ net1786 net173 net620 vssd1 vssd1 vccd1 vccd1 _00241_ sky130_fd_sc_hd__mux2_1
XFILLER_0_188_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11237__B top.lcd.nextState\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_160_2845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12495__RESET_B net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10568__S net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11989_ _05866_ _05869_ _05870_ vssd1 vssd1 vccd1 vccd1 _05872_ sky130_fd_sc_hd__and3_1
XFILLER_0_58_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_193_3344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13728_ clknet_leaf_93_clk _01299_ vssd1 vssd1 vccd1 vccd1 top.a1.dataInTemp\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_50_clk_A clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_692 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13659_ clknet_leaf_92_clk _01235_ net995 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[105\]
+ sky130_fd_sc_hd__dfrtp_1
X_06200_ wb.curr_state\[0\] _01430_ vssd1 vssd1 vccd1 vccd1 _01431_ sky130_fd_sc_hd__nand2_1
XANTENNA__07409__B1 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_140_Right_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07180_ _02312_ _02314_ _02316_ _02318_ vssd1 vssd1 vccd1 vccd1 _02319_ sky130_fd_sc_hd__or4_2
XFILLER_0_41_312 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_65_clk_A clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_197_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07188__A2 net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout406 _04717_ vssd1 vssd1 vccd1 vccd1 net406 sky130_fd_sc_hd__clkbuf_4
X_09821_ _04833_ _04836_ vssd1 vssd1 vccd1 vccd1 _04837_ sky130_fd_sc_hd__xor2_1
Xfanout428 net430 vssd1 vssd1 vccd1 vccd1 net428 sky130_fd_sc_hd__clkbuf_4
Xfanout439 _01566_ vssd1 vssd1 vccd1 vccd1 net439 sky130_fd_sc_hd__clkbuf_8
XANTENNA__06935__A2 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_123_clk_A clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09752_ _04772_ _04773_ _04151_ vssd1 vssd1 vccd1 vccd1 _04775_ sky130_fd_sc_hd__a21o_1
X_06964_ top.DUT.register\[18\]\[23\] net548 net533 top.DUT.register\[12\]\[23\] vssd1
+ vssd1 vccd1 vccd1 _02103_ sky130_fd_sc_hd__a22o_1
X_08703_ _03821_ vssd1 vssd1 vccd1 vccd1 _03822_ sky130_fd_sc_hd__inv_2
XFILLER_0_198_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_146_62 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06895_ top.DUT.register\[10\]\[18\] net772 net642 top.DUT.register\[8\]\[18\] _02033_
+ vssd1 vssd1 vccd1 vccd1 _02034_ sky130_fd_sc_hd__a221o_1
X_09683_ top.a1.instruction\[7\] top.a1.instruction\[8\] top.a1.instruction\[9\] net786
+ vssd1 vssd1 vccd1 vccd1 _04719_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_87_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08634_ _03714_ _03755_ net289 vssd1 vssd1 vccd1 vccd1 _03756_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_87_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07896__B1 net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07360__A2 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08565_ _03504_ _03689_ net296 vssd1 vssd1 vccd1 vccd1 _03690_ sky130_fd_sc_hd__mux2_1
XANTENNA__10478__S net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout442_A _01566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08456__B _03534_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_194_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07648__B1 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07516_ _02633_ _02653_ vssd1 vssd1 vccd1 vccd1 _02655_ sky130_fd_sc_hd__nand2_1
XANTENNA_clkbuf_leaf_18_clk_A clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08496_ _02307_ net431 net499 _02309_ vssd1 vssd1 vccd1 vccd1 _03624_ sky130_fd_sc_hd__a22o_1
XFILLER_0_18_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07112__A2 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_146_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07447_ top.DUT.register\[6\]\[15\] net568 net440 top.DUT.register\[5\]\[15\] _02585_
+ vssd1 vssd1 vccd1 vccd1 _02586_ sky130_fd_sc_hd__a221o_1
XFILLER_0_162_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout230_X net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout707_A _01640_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_2213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_539 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07378_ top.DUT.register\[13\]\[8\] net774 net743 top.DUT.register\[2\]\[8\] _02516_
+ vssd1 vssd1 vccd1 vccd1 _02517_ sky130_fd_sc_hd__a221o_1
XANTENNA_clkbuf_3_5_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06329_ _01475_ vssd1 vssd1 vccd1 vccd1 _01476_ sky130_fd_sc_hd__inv_2
X_09117_ _03000_ _03040_ vssd1 vssd1 vccd1 vccd1 _04192_ sky130_fd_sc_hd__and2_1
XANTENNA__07359__Y _02498_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_2413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09048_ net320 _03625_ _04120_ _04122_ vssd1 vssd1 vccd1 vccd1 _04123_ sky130_fd_sc_hd__o211a_1
XANTENNA__09855__X _04868_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07820__B1 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12823__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout697_X net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10941__S net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold460 top.DUT.register\[15\]\[29\] vssd1 vssd1 vccd1 vccd1 net1576 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08972__A2_N net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold471 top.DUT.register\[11\]\[23\] vssd1 vssd1 vccd1 vccd1 net1587 sky130_fd_sc_hd__dlygate4sd3_1
Xhold482 top.DUT.register\[1\]\[28\] vssd1 vssd1 vccd1 vccd1 net1598 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07179__A2 net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11010_ wb.curr_state\[1\] net1 vssd1 vssd1 vccd1 vccd1 _05041_ sky130_fd_sc_hd__and2_1
Xhold493 top.DUT.register\[16\]\[4\] vssd1 vssd1 vccd1 vccd1 net1609 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06387__B1 net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06926__A2 net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout940 net943 vssd1 vssd1 vccd1 vccd1 net940 sky130_fd_sc_hd__clkbuf_4
Xfanout951 net952 vssd1 vssd1 vccd1 vccd1 net951 sky130_fd_sc_hd__clkbuf_2
Xfanout962 net965 vssd1 vssd1 vccd1 vccd1 net962 sky130_fd_sc_hd__buf_2
Xfanout973 net974 vssd1 vssd1 vccd1 vccd1 net973 sky130_fd_sc_hd__clkbuf_4
Xfanout984 net985 vssd1 vssd1 vccd1 vccd1 net984 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_129_2375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout995 net997 vssd1 vssd1 vccd1 vccd1 net995 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_129_2386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12961_ clknet_leaf_17_clk _00553_ net965 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[14\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_99_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1160 top.DUT.register\[8\]\[9\] vssd1 vssd1 vccd1 vccd1 net2276 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1171 top.DUT.register\[10\]\[29\] vssd1 vssd1 vccd1 vccd1 net2287 sky130_fd_sc_hd__dlygate4sd3_1
X_11912_ _05770_ _05788_ vssd1 vssd1 vccd1 vccd1 _05795_ sky130_fd_sc_hd__xnor2_1
Xhold1182 top.DUT.register\[24\]\[18\] vssd1 vssd1 vccd1 vccd1 net2298 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07887__B1 net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12892_ clknet_leaf_130_clk _00484_ net909 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[12\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1193 top.ramload\[20\] vssd1 vssd1 vccd1 vccd1 net2309 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_206_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07351__A2 net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_142_2575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10388__S net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11843_ _05723_ _05725_ vssd1 vssd1 vccd1 vccd1 _05726_ sky130_fd_sc_hd__nor2_1
XANTENNA__12176__A1_N _05083_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_540 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07270__B _02408_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11774_ _05655_ _05656_ vssd1 vssd1 vccd1 vccd1 _05657_ sky130_fd_sc_hd__nand2_1
XFILLER_0_95_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_175_3074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13513_ clknet_leaf_51_clk _01105_ net1036 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[31\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_10725_ net2120 net153 net336 vssd1 vssd1 vccd1 vccd1 _00886_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13444_ clknet_leaf_36_clk _01036_ net1050 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[29\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13723__RESET_B net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10656_ net162 net1851 net344 vssd1 vssd1 vccd1 vccd1 _00820_ sky130_fd_sc_hd__mux2_1
XFILLER_0_192_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload16 clknet_leaf_122_clk vssd1 vssd1 vccd1 vccd1 clkload16/Y sky130_fd_sc_hd__inv_8
X_10587_ net1648 net174 net352 vssd1 vssd1 vccd1 vccd1 _00753_ sky130_fd_sc_hd__mux2_1
Xclkload27 clknet_leaf_114_clk vssd1 vssd1 vccd1 vccd1 clkload27/Y sky130_fd_sc_hd__inv_8
X_13375_ clknet_leaf_15_clk _00967_ net961 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[27\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_140_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkload38 clknet_leaf_95_clk vssd1 vssd1 vccd1 vccd1 clkload38/Y sky130_fd_sc_hd__inv_6
XTAP_TAPCELL_ROW_58_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload49 clknet_leaf_111_clk vssd1 vssd1 vccd1 vccd1 clkload49/X sky130_fd_sc_hd__clkbuf_8
X_12326_ top.pad.button_control.r_counter\[9\] _06126_ net791 vssd1 vssd1 vccd1 vccd1
+ _06128_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_23_378 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12405__Q top.a1.instruction\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10851__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12257_ net1121 _06084_ _06085_ vssd1 vssd1 vccd1 vccd1 _01328_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12191__X _06049_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09925__B _04628_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08367__A1 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11208_ _05110_ net1261 net471 vssd1 vssd1 vccd1 vccd1 _01254_ sky130_fd_sc_hd__mux2_1
X_12188_ top.a1.row2\[43\] net847 net797 _05657_ vssd1 vssd1 vccd1 vccd1 _01296_ sky130_fd_sc_hd__a22o_1
XANTENNA__10174__A1 net156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06917__A2 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11139_ net61 net868 vssd1 vssd1 vccd1 vccd1 _05075_ sky130_fd_sc_hd__and2_1
XFILLER_0_207_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09941__A net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_183_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09867__A1 net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_204_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06680_ top.DUT.register\[4\]\[26\] net670 net776 top.DUT.register\[13\]\[26\] _01818_
+ vssd1 vssd1 vccd1 vccd1 _01819_ sky130_fd_sc_hd__a221o_1
XANTENNA__07878__B1 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07342__A2 net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10298__S net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_69_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06550__B1 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08276__B _02899_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_175_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08350_ net436 _03477_ _03483_ net427 _03479_ vssd1 vssd1 vccd1 vccd1 _03484_ sky130_fd_sc_hd__a221o_1
XFILLER_0_86_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07301_ top.DUT.register\[24\]\[12\] net511 net447 top.DUT.register\[21\]\[12\] _02439_
+ vssd1 vssd1 vccd1 vccd1 _02440_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_82_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08281_ _03285_ _03289_ vssd1 vssd1 vccd1 vccd1 _03417_ sky130_fd_sc_hd__nand2_1
XFILLER_0_191_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_190_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07232_ top.DUT.register\[17\]\[10\] net746 net722 top.DUT.register\[29\]\[10\] vssd1
+ vssd1 vccd1 vccd1 _02371_ sky130_fd_sc_hd__a22o_1
XANTENNA__11711__A top.a1.dataIn\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07163_ top.DUT.register\[3\]\[11\] net702 _02299_ _02301_ vssd1 vssd1 vccd1 vccd1
+ _02302_ sky130_fd_sc_hd__a211o_1
XFILLER_0_143_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07802__B1 net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07094_ top.DUT.register\[15\]\[16\] net680 net676 top.DUT.register\[31\]\[16\] vssd1
+ vssd1 vccd1 vccd1 _02233_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_113_2143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10761__S net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout203 net206 vssd1 vssd1 vccd1 vccd1 net203 sky130_fd_sc_hd__buf_2
Xfanout214 _04771_ vssd1 vssd1 vccd1 vccd1 net214 sky130_fd_sc_hd__clkbuf_2
XANTENNA__06540__A _01678_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout225 _04805_ vssd1 vssd1 vccd1 vccd1 net225 sky130_fd_sc_hd__buf_2
Xfanout236 _04757_ vssd1 vssd1 vccd1 vccd1 net236 sky130_fd_sc_hd__buf_1
Xfanout247 _04749_ vssd1 vssd1 vccd1 vccd1 net247 sky130_fd_sc_hd__clkbuf_2
X_09804_ _04151_ _04821_ _04816_ vssd1 vssd1 vccd1 vccd1 _04822_ sky130_fd_sc_hd__o21ai_1
Xfanout258 _04737_ vssd1 vssd1 vccd1 vccd1 net258 sky130_fd_sc_hd__clkbuf_2
Xfanout269 _04726_ vssd1 vssd1 vccd1 vccd1 net269 sky130_fd_sc_hd__buf_2
X_07996_ top.DUT.register\[28\]\[31\] net767 _03129_ _03134_ vssd1 vssd1 vccd1 vccd1
+ _03135_ sky130_fd_sc_hd__a211o_1
XANTENNA__07581__A2 net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09851__A top.pc\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09735_ net826 _04312_ _04752_ top.a1.dataIn\[10\] vssd1 vssd1 vccd1 vccd1 _04761_
+ sky130_fd_sc_hd__a2bb2o_1
X_06947_ top.DUT.register\[20\]\[21\] net666 net716 top.DUT.register\[27\]\[21\] _02085_
+ vssd1 vssd1 vccd1 vccd1 _02086_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout657_A _01609_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07869__B1 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09666_ top.pc\[1\] _02952_ _04201_ net806 vssd1 vssd1 vccd1 vccd1 _04703_ sky130_fd_sc_hd__o22a_1
X_06878_ top.DUT.register\[15\]\[18\] net681 net677 top.DUT.register\[31\]\[18\] vssd1
+ vssd1 vccd1 vccd1 _02017_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_2_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_715 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08617_ net323 _03739_ vssd1 vssd1 vccd1 vccd1 _03740_ sky130_fd_sc_hd__or2_1
XANTENNA__06541__B1 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout445_X net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09597_ _04627_ _04631_ _04629_ vssd1 vssd1 vccd1 vccd1 _04643_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout824_A net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09997__S net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10001__S net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08548_ _03273_ _03278_ vssd1 vssd1 vccd1 vccd1 _03674_ sky130_fd_sc_hd__nand2_1
XFILLER_0_77_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_415 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_595 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout612_X net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10936__S net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08479_ _02387_ net431 net499 _02386_ vssd1 vssd1 vccd1 vccd1 _03608_ sky130_fd_sc_hd__a22o_1
XFILLER_0_147_472 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11621__A top.a1.dataIn\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10510_ net1988 net198 net358 vssd1 vssd1 vccd1 vccd1 _00679_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11490_ _05370_ _05371_ _05367_ _05368_ vssd1 vssd1 vccd1 vccd1 _05373_ sky130_fd_sc_hd__a211o_1
XANTENNA__06715__A _01853_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_598 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_464 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10441_ net219 net2275 net365 vssd1 vssd1 vccd1 vccd1 _00612_ sky130_fd_sc_hd__mux2_1
X_10372_ net2089 net230 net373 vssd1 vssd1 vccd1 vccd1 _00547_ sky130_fd_sc_hd__mux2_1
X_13160_ clknet_leaf_27_clk _00752_ net1008 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[20\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_12111_ _05970_ _05993_ vssd1 vssd1 vccd1 vccd1 _05994_ sky130_fd_sc_hd__xor2_2
X_13091_ clknet_leaf_49_clk _00683_ net1061 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[18\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10671__S net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12042_ _05887_ _05888_ net125 vssd1 vssd1 vccd1 vccd1 _05925_ sky130_fd_sc_hd__o21ba_1
Xhold290 top.DUT.register\[11\]\[30\] vssd1 vssd1 vccd1 vccd1 net1406 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10156__A1 net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_144_2604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07572__A2 net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout770 _01614_ vssd1 vssd1 vccd1 vccd1 net770 sky130_fd_sc_hd__clkbuf_8
Xfanout781 _01603_ vssd1 vssd1 vccd1 vccd1 net781 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_205_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout792 _01590_ vssd1 vssd1 vccd1 vccd1 net792 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_189_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12719__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12944_ clknet_leaf_29_clk _00536_ net1017 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[13\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_201_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_177_3103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11120__A3 net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12875_ clknet_leaf_45_clk _00467_ net1065 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[11\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06532__B1 net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11826_ _05673_ net131 _05675_ vssd1 vssd1 vccd1 vccd1 _05709_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_190_3303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11757_ _05599_ _05639_ vssd1 vssd1 vccd1 vccd1 _05640_ sky130_fd_sc_hd__xor2_2
XANTENNA__10846__S net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10708_ net1410 net213 net334 vssd1 vssd1 vccd1 vccd1 _00869_ sky130_fd_sc_hd__mux2_1
XFILLER_0_181_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_165_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_153_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11688_ _05537_ _05570_ vssd1 vssd1 vccd1 vccd1 _05571_ sky130_fd_sc_hd__nand2_1
XANTENNA__06625__A _01754_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_155_2766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_155_2777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload105 clknet_leaf_62_clk vssd1 vssd1 vccd1 vccd1 clkload105/Y sky130_fd_sc_hd__clkinv_8
X_13427_ clknet_leaf_122_clk _01019_ net934 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[29\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11250__B _05118_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10639_ net228 net1704 net342 vssd1 vssd1 vccd1 vccd1 _00803_ sky130_fd_sc_hd__mux2_1
XFILLER_0_180_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_188 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09785__B1 net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13358_ clknet_leaf_41_clk _00950_ net1047 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[26\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06599__B1 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_188_3265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_140_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12309_ top.pad.button_control.r_counter\[3\] _06114_ vssd1 vssd1 vccd1 vccd1 _06117_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_11_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10581__S net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13289_ clknet_leaf_21_clk _00881_ net1034 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[24\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_18_Right_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_194_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07850_ top.DUT.register\[12\]\[0\] net531 net523 top.DUT.register\[11\]\[0\] vssd1
+ vssd1 vccd1 vccd1 _02989_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_3_Left_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06801_ _01930_ _01939_ vssd1 vssd1 vccd1 vccd1 _01940_ sky130_fd_sc_hd__nor2_4
X_07781_ top.DUT.register\[8\]\[2\] net639 net702 top.DUT.register\[3\]\[2\] vssd1
+ vssd1 vccd1 vccd1 _02920_ sky130_fd_sc_hd__a22o_1
Xinput3 DAT_I[10] vssd1 vssd1 vccd1 vccd1 net3 sky130_fd_sc_hd__clkbuf_1
X_09520_ top.pc\[25\] _04543_ _04553_ vssd1 vssd1 vccd1 vccd1 _04571_ sky130_fd_sc_hd__a21o_1
X_06732_ _01865_ _01866_ _01868_ _01870_ vssd1 vssd1 vccd1 vccd1 _01871_ sky130_fd_sc_hd__or4_1
XANTENNA__09390__B _04438_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07903__B _03040_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire413_X net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07315__A2 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06663_ top.DUT.register\[2\]\[26\] net562 net518 top.DUT.register\[7\]\[26\] vssd1
+ vssd1 vccd1 vccd1 _01802_ sky130_fd_sc_hd__a22o_1
X_09451_ top.pc\[21\] top.pc\[22\] _04478_ vssd1 vssd1 vccd1 vccd1 _04506_ sky130_fd_sc_hd__and3_1
XANTENNA__06523__B1 net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08402_ net324 net315 vssd1 vssd1 vccd1 vccd1 _03534_ sky130_fd_sc_hd__or2_4
XFILLER_0_47_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06594_ _01724_ _01726_ _01731_ _01732_ vssd1 vssd1 vccd1 vccd1 _01733_ sky130_fd_sc_hd__or4_1
XFILLER_0_47_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09382_ _04440_ _04441_ _04436_ vssd1 vssd1 vccd1 vccd1 _04442_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_27_Right_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08333_ net313 _03320_ vssd1 vssd1 vccd1 vccd1 _03467_ sky130_fd_sc_hd__or2_1
XFILLER_0_176_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10756__S net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_125_clk clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_125_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_157_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout238_A _04757_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_634 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08264_ net276 _03295_ _03399_ vssd1 vssd1 vccd1 vccd1 _03400_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_191_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07215_ _01477_ _01488_ _02353_ vssd1 vssd1 vccd1 vccd1 _02354_ sky130_fd_sc_hd__o21a_1
X_08195_ net316 net302 vssd1 vssd1 vccd1 vccd1 _03333_ sky130_fd_sc_hd__or2_1
XANTENNA__06254__B net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout405_A net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08579__A1 _03342_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07146_ _02278_ _02280_ _02282_ _02284_ vssd1 vssd1 vccd1 vccd1 _02285_ sky130_fd_sc_hd__or4_2
XFILLER_0_14_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11178__A3 net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08579__B2 net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_95_1868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10491__S net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07077_ top.DUT.register\[21\]\[22\] net656 net718 top.DUT.register\[19\]\[22\] _02210_
+ vssd1 vssd1 vccd1 vccd1 _02216_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_36_Right_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_168_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06270__A top.ramload\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout774_A net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1009 net1016 vssd1 vssd1 vccd1 vccd1 net1009 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout395_X net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_hold185_A top.edg2.flip1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08751__B2 net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06762__B1 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout562_X net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07979_ top.DUT.register\[3\]\[31\] net553 net506 top.DUT.register\[27\]\[31\] vssd1
+ vssd1 vccd1 vccd1 _03118_ sky130_fd_sc_hd__a22o_1
X_09718_ top.a1.dataIn\[7\] net795 net799 top.pc\[7\] _04746_ vssd1 vssd1 vccd1 vccd1
+ _04747_ sky130_fd_sc_hd__a221o_1
X_10990_ net1285 _05026_ net589 vssd1 vssd1 vccd1 vccd1 _01120_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07306__A2 net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11102__A3 net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09700__B1 net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09649_ _04686_ _04687_ _04688_ _04690_ vssd1 vssd1 vccd1 vccd1 _04691_ sky130_fd_sc_hd__or4_1
XANTENNA__06514__B1 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08957__A1_N _02428_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_45_Right_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout827_X net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12660_ clknet_leaf_58_clk _00252_ net1075 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[5\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08925__A net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11611_ _05493_ vssd1 vssd1 vccd1 vccd1 _05494_ sky130_fd_sc_hd__inv_2
XFILLER_0_93_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13315__RESET_B net1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10666__S net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_182_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_172_3022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_116_clk clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_116_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_108_612 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12591_ clknet_leaf_21_clk _00183_ net1033 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[2\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_148_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_67_Left_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_182_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_172_3033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11542_ _05419_ _05420_ _05424_ vssd1 vssd1 vccd1 vccd1 _05425_ sky130_fd_sc_hd__a21o_1
XFILLER_0_9_180 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xwire412 _02260_ vssd1 vssd1 vccd1 vccd1 net412 sky130_fd_sc_hd__buf_2
XFILLER_0_37_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_208_Left_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_163_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11473_ _05319_ _05322_ _05321_ vssd1 vssd1 vccd1 vccd1 _05356_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_137_2496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13212_ clknet_leaf_130_clk _00804_ net910 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[22\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_10424_ net2130 net162 net370 vssd1 vssd1 vccd1 vccd1 _00596_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_54_Right_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13143_ clknet_leaf_2_clk _00735_ net914 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[20\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_10355_ net1515 net167 net378 vssd1 vssd1 vccd1 vccd1 _00531_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09475__B _02111_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_150_2696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07793__A2 net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10286_ net1587 net178 net388 vssd1 vssd1 vccd1 vccd1 _00464_ sky130_fd_sc_hd__mux2_1
X_13074_ clknet_leaf_31_clk _00666_ net1021 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[18\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_76_Left_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12025_ _05882_ _05907_ vssd1 vssd1 vccd1 vccd1 _05908_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_183_3184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_183_3195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07545__A2 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06753__B1 net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_63_Right_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12927_ clknet_leaf_15_clk _00519_ net961 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[13\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06505__B1 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12858_ clknet_leaf_5_clk _00450_ net936 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[11\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_85_Left_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_157_2806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_201_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11809_ _05668_ net131 _05659_ vssd1 vssd1 vccd1 vccd1 _05692_ sky130_fd_sc_hd__a21o_1
XANTENNA__13056__RESET_B net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_185_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13047__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_107_clk clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_107_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__10576__S net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12789_ clknet_leaf_31_clk _00381_ net1023 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[9\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_77 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_773 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06284__A2 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07000_ top.DUT.register\[10\]\[20\] net521 net442 top.DUT.register\[5\]\[20\] vssd1
+ vssd1 vccd1 vccd1 _02139_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_72_Right_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_141_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_110_2102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08951_ net1207 net873 _02701_ net693 vssd1 vssd1 vccd1 vccd1 _00057_ sky130_fd_sc_hd__a22o_1
XANTENNA__12620__RESET_B net1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_168_2968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07902_ net295 _03040_ vssd1 vssd1 vccd1 vccd1 _03041_ sky130_fd_sc_hd__nor2_1
X_08882_ _01744_ _03974_ _01743_ vssd1 vssd1 vccd1 vccd1 _03992_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_4_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_205_3519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07536__A2 net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07833_ top.DUT.register\[27\]\[0\] net715 _02964_ _02967_ _02971_ vssd1 vssd1 vccd1
+ vccd1 _02972_ sky130_fd_sc_hd__a2111oi_1
XANTENNA__10540__A1 net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06744__B1 net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_81_Right_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout188_A net191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07764_ net410 _02854_ _02902_ net804 vssd1 vssd1 vccd1 vccd1 _02903_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_108_2064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09503_ _04553_ _04554_ vssd1 vssd1 vccd1 vccd1 _04555_ sky130_fd_sc_hd__or2_1
X_06715_ _01853_ vssd1 vssd1 vccd1 vccd1 _01854_ sky130_fd_sc_hd__inv_2
X_07695_ top.DUT.register\[19\]\[4\] net537 net461 top.DUT.register\[17\]\[4\] _02833_
+ vssd1 vssd1 vccd1 vccd1 _02834_ sky130_fd_sc_hd__a221o_1
XFILLER_0_2_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06249__B net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout355_A net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1097_A net1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09434_ _04472_ _04488_ _04489_ net811 vssd1 vssd1 vccd1 vccd1 _04491_ sky130_fd_sc_hd__a31o_1
X_06646_ _01764_ _01784_ vssd1 vssd1 vccd1 vccd1 _01785_ sky130_fd_sc_hd__and2b_1
XFILLER_0_94_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_121_2264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_707 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_148 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09365_ net132 _04418_ _04425_ net811 net900 vssd1 vssd1 vccd1 vccd1 _04426_ sky130_fd_sc_hd__o221a_1
XANTENNA__10486__S net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06577_ top.DUT.register\[16\]\[28\] net545 net537 top.DUT.register\[19\]\[28\] vssd1
+ vssd1 vccd1 vccd1 _01716_ sky130_fd_sc_hd__a22o_1
XFILLER_0_90_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08316_ _03379_ _03449_ net292 vssd1 vssd1 vccd1 vccd1 _03451_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06265__A top.ramload\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09296_ top.pc\[12\] top.pc\[13\] _04326_ vssd1 vssd1 vccd1 vccd1 _04360_ sky130_fd_sc_hd__and3_1
XFILLER_0_117_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_191_378 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_90_Right_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_97_1908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08247_ _03042_ _03179_ _03041_ vssd1 vssd1 vccd1 vccd1 _03384_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_132_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08178_ _01764_ net329 _03315_ vssd1 vssd1 vccd1 vccd1 _03316_ sky130_fd_sc_hd__o21a_1
XFILLER_0_160_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09213__A2 top.pc\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout891_A net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout989_A net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11020__A2 net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07129_ top.DUT.register\[16\]\[11\] net543 net539 top.DUT.register\[8\]\[11\] vssd1
+ vssd1 vccd1 vccd1 _02268_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_37_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10140_ net162 net1548 net610 vssd1 vssd1 vccd1 vccd1 _00340_ sky130_fd_sc_hd__mux2_1
XANTENNA__07775__A2 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09863__X _04875_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_180 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout777_X net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10071_ net1949 net175 net618 vssd1 vssd1 vccd1 vccd1 _00273_ sky130_fd_sc_hd__mux2_1
XANTENNA__07527__A2 net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07383__X _02522_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13830_ net1114 vssd1 vssd1 vccd1 vccd1 gpio_out[29] sky130_fd_sc_hd__buf_2
X_13761_ clknet_leaf_70_clk _01332_ vssd1 vssd1 vccd1 vccd1 top.lcd.currentState\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_10973_ top.a1.dataIn\[2\] net849 _05011_ _05013_ vssd1 vssd1 vccd1 vccd1 _05014_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_69_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12712_ clknet_leaf_8_clk _00304_ net947 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[6\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_179_191 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13692_ clknet_leaf_72_clk _00004_ vssd1 vssd1 vccd1 vccd1 top.lcd.nextState\[5\]
+ sky130_fd_sc_hd__dfxtp_2
XANTENNA__07160__B1 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12643_ clknet_leaf_60_clk _00235_ net1088 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[4\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_139_2525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06446__Y _01585_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_139_2536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06175__A top.a1.halfData\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12574_ clknet_leaf_18_clk _00166_ net1026 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[2\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_170_507 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_250 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11525_ _05376_ _05401_ vssd1 vssd1 vccd1 vccd1 _05408_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_152_2725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09486__A top.pc\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11456_ _05292_ _05332_ vssd1 vssd1 vccd1 vccd1 _05339_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_33_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_150_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_827 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10407_ net228 net2068 _04984_ vssd1 vssd1 vccd1 vccd1 _00579_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11387_ top.a1.dataIn\[26\] _05238_ top.a1.dataIn\[27\] vssd1 vssd1 vccd1 vccd1 _05270_
+ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_185_3224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07766__A2 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13126_ clknet_leaf_40_clk _00718_ net1053 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[19\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_103_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10338_ net1633 net233 net380 vssd1 vssd1 vccd1 vccd1 _00514_ sky130_fd_sc_hd__mux2_1
XANTENNA__06974__B1 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12413__Q top.a1.instruction\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13057_ clknet_leaf_16_clk _00649_ net963 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[17\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_10269_ net2182 net244 net385 vssd1 vssd1 vccd1 vccd1 _00447_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08715__A1 _02156_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12008_ _05865_ _05872_ net126 vssd1 vssd1 vccd1 vccd1 _05891_ sky130_fd_sc_hd__nand3_1
XANTENNA__06726__B1 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_788 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_163_2887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_163_2898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_99 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_187_Right_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08479__B1 net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_93_Left_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_200_3449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06500_ top.DUT.register\[27\]\[30\] net716 net712 top.DUT.register\[11\]\[30\] vssd1
+ vssd1 vccd1 vccd1 _01639_ sky130_fd_sc_hd__a22o_1
XFILLER_0_48_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07480_ top.DUT.register\[6\]\[14\] net568 net536 top.DUT.register\[19\]\[14\] vssd1
+ vssd1 vccd1 vccd1 _02619_ sky130_fd_sc_hd__a22o_1
XANTENNA__07151__B1 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_707 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_196_3386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09691__A2 net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_186_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_174_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_201_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06431_ _01551_ _01557_ _01563_ _01569_ vssd1 vssd1 vccd1 vccd1 _01570_ sky130_fd_sc_hd__or4_1
XFILLER_0_57_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_173_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_17_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06362_ net896 _01473_ vssd1 vssd1 vccd1 vccd1 _01501_ sky130_fd_sc_hd__nand2_2
XFILLER_0_72_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09150_ _04221_ _04222_ vssd1 vssd1 vccd1 vccd1 _04223_ sky130_fd_sc_hd__or2_1
XFILLER_0_44_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08101_ _02633_ net299 vssd1 vssd1 vccd1 vccd1 _03240_ sky130_fd_sc_hd__nand2_1
XFILLER_0_71_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09081_ top.a1.instruction\[7\] top.a1.instruction\[8\] vssd1 vssd1 vccd1 vccd1 _04156_
+ sky130_fd_sc_hd__nand2_1
X_06293_ _01330_ vssd1 vssd1 vccd1 vccd1 _01451_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_79_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08032_ net319 net315 vssd1 vssd1 vccd1 vccd1 _03171_ sky130_fd_sc_hd__or2_2
XANTENNA__09396__A _02016_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold801 top.DUT.register\[14\]\[30\] vssd1 vssd1 vccd1 vccd1 net1917 sky130_fd_sc_hd__dlygate4sd3_1
Xhold812 top.DUT.register\[13\]\[12\] vssd1 vssd1 vccd1 vccd1 net1928 sky130_fd_sc_hd__dlygate4sd3_1
Xhold823 top.DUT.register\[30\]\[16\] vssd1 vssd1 vccd1 vccd1 net1939 sky130_fd_sc_hd__dlygate4sd3_1
Xhold834 top.DUT.register\[7\]\[15\] vssd1 vssd1 vccd1 vccd1 net1950 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_1827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold845 top.DUT.register\[16\]\[3\] vssd1 vssd1 vccd1 vccd1 net1961 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07757__A2 net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold856 top.DUT.register\[7\]\[30\] vssd1 vssd1 vccd1 vccd1 net1972 sky130_fd_sc_hd__dlygate4sd3_1
Xhold867 top.DUT.register\[23\]\[30\] vssd1 vssd1 vccd1 vccd1 net1983 sky130_fd_sc_hd__dlygate4sd3_1
Xhold878 top.DUT.register\[5\]\[28\] vssd1 vssd1 vccd1 vccd1 net1994 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08954__B2 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09983_ net260 net1775 net624 vssd1 vssd1 vccd1 vccd1 _00188_ sky130_fd_sc_hd__mux2_1
Xhold889 top.DUT.register\[7\]\[4\] vssd1 vssd1 vccd1 vccd1 net2005 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06965__B1 net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08934_ _03102_ _03145_ vssd1 vssd1 vccd1 vccd1 _04042_ sky130_fd_sc_hd__xor2_1
XFILLER_0_110_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1012_A net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07509__A2 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08865_ net277 _03937_ vssd1 vssd1 vccd1 vccd1 _03976_ sky130_fd_sc_hd__and2_1
XANTENNA__06717__B1 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07816_ top.DUT.register\[15\]\[0\] net706 net698 top.DUT.register\[31\]\[0\] vssd1
+ vssd1 vccd1 vccd1 _02955_ sky130_fd_sc_hd__a22o_1
XFILLER_0_165_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08796_ net883 top.pc\[24\] net694 _03910_ vssd1 vssd1 vccd1 vccd1 _03911_ sky130_fd_sc_hd__a22o_1
XANTENNA__07390__B1 net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07747_ top.DUT.register\[3\]\[3\] net553 net453 top.DUT.register\[29\]\[3\] _02885_
+ vssd1 vssd1 vccd1 vccd1 _02886_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_154_Right_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout358_X net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09131__A1 top.pc\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07142__B1 net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07678_ _02811_ _02814_ _02815_ _02816_ vssd1 vssd1 vccd1 vccd1 _02817_ sky130_fd_sc_hd__or4_2
XANTENNA__09682__A2 top.a1.instruction\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_177_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_0_Right_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_36_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09417_ _04469_ _04474_ vssd1 vssd1 vccd1 vccd1 _04475_ sky130_fd_sc_hd__xor2_1
XFILLER_0_149_375 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06629_ top.DUT.register\[2\]\[27\] net745 net701 top.DUT.register\[31\]\[27\] vssd1
+ vssd1 vccd1 vccd1 _01768_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout525_X net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_176_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09348_ net903 top.pc\[15\] _04409_ net892 vssd1 vssd1 vccd1 vccd1 _00095_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_101_1956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_1967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_43_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10944__S net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09279_ net903 top.pc\[11\] _04344_ net892 vssd1 vssd1 vccd1 vccd1 _00091_ sky130_fd_sc_hd__o211a_1
X_11310_ top.a1.row1\[15\] _05130_ _05123_ vssd1 vssd1 vccd1 vccd1 _05196_ sky130_fd_sc_hd__o21a_1
XANTENNA__07996__A2 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12290_ top.lcd.cnt_500hz\[13\] top.lcd.cnt_500hz\[12\] _06101_ vssd1 vssd1 vccd1
+ vccd1 _06105_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_134_2455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11241_ net880 _01382_ _05128_ _05133_ vssd1 vssd1 vccd1 vccd1 _05134_ sky130_fd_sc_hd__and4_1
XFILLER_0_30_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07748__A2 net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11172_ _05090_ _05095_ _05085_ vssd1 vssd1 vccd1 vccd1 _05096_ sky130_fd_sc_hd__a21bo_1
XANTENNA__06956__B1 net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10123_ net229 net1532 net607 vssd1 vssd1 vccd1 vccd1 _00323_ sky130_fd_sc_hd__mux2_1
XANTENNA__09753__B _04172_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10054_ net1842 net245 net615 vssd1 vssd1 vccd1 vccd1 _00256_ sky130_fd_sc_hd__mux2_1
XANTENNA_input33_A DAT_I[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_180_3143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_199_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_203_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13813_ top.lcd.lcd_rs vssd1 vssd1 vccd1 vccd1 net111 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08656__Y _03777_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_774 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_121_Right_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_187_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_262 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13744_ clknet_leaf_100_clk _01315_ vssd1 vssd1 vccd1 vccd1 top.lcd.cnt_20ms\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_10956_ _04657_ _04998_ vssd1 vssd1 vccd1 vccd1 _04999_ sky130_fd_sc_hd__nor2_1
XANTENNA__07133__B1 net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13675_ clknet_leaf_90_clk _01251_ net999 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_10887_ net140 net2203 net596 vssd1 vssd1 vccd1 vccd1 _01048_ sky130_fd_sc_hd__mux2_1
XFILLER_0_155_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12626_ clknet_leaf_23_clk _00218_ net1015 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[4\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_159_Left_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12557_ clknet_leaf_42_clk _00149_ net1064 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[1\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10854__S net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_182_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11508_ _05385_ _05386_ _05390_ vssd1 vssd1 vccd1 vccd1 _05391_ sky130_fd_sc_hd__mux2_1
XANTENNA__07987__A2 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_540 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12488_ clknet_leaf_74_clk _00009_ net1077 vssd1 vssd1 vccd1 vccd1 top.a1.hexop\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold108 top.ramload\[4\] vssd1 vssd1 vccd1 vccd1 net1224 sky130_fd_sc_hd__dlygate4sd3_1
Xhold119 top.ramstore\[28\] vssd1 vssd1 vccd1 vccd1 net1235 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11439_ _05272_ _05309_ vssd1 vssd1 vccd1 vccd1 _05322_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_123_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08936__A1 net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09944__A net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_186_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_74_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06947__B1 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10743__A1 net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_192_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13109_ clknet_leaf_32_clk _00701_ net1044 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[19\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_165_2916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_168_Left_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06980_ top.DUT.register\[2\]\[23\] net744 net717 top.DUT.register\[27\]\[23\] vssd1
+ vssd1 vccd1 vccd1 _02119_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_165_2927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11299__A2 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08650_ _02049_ _03769_ vssd1 vssd1 vccd1 vccd1 _03771_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_198_3415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07372__B1 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07601_ _02734_ _02737_ _02738_ _02739_ vssd1 vssd1 vccd1 vccd1 _02740_ sky130_fd_sc_hd__or4_1
XANTENNA__07911__A2 _02899_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_2023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08581_ net885 top.pc\[14\] net696 _03705_ vssd1 vssd1 vccd1 vccd1 _03706_ sky130_fd_sc_hd__a22o_1
XANTENNA__08566__Y _03691_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07532_ top.DUT.register\[28\]\[7\] net555 net511 top.DUT.register\[24\]\[7\] vssd1
+ vssd1 vccd1 vccd1 _02671_ sky130_fd_sc_hd__a22o_1
XFILLER_0_88_295 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07463_ top.DUT.register\[22\]\[15\] net648 net727 top.DUT.register\[18\]\[15\] _02595_
+ vssd1 vssd1 vccd1 vccd1 _02602_ sky130_fd_sc_hd__a221o_1
XANTENNA__08872__B1 net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09202_ top.pc\[7\] _02728_ vssd1 vssd1 vccd1 vccd1 _04272_ sky130_fd_sc_hd__xnor2_1
X_06414_ net684 _01521_ _01523_ vssd1 vssd1 vccd1 vccd1 _01553_ sky130_fd_sc_hd__and3_4
XANTENNA__09678__X _04714_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07394_ top.DUT.register\[13\]\[9\] net463 net507 top.DUT.register\[4\]\[9\] _02532_
+ vssd1 vssd1 vccd1 vccd1 _02533_ sky130_fd_sc_hd__a221o_1
X_09133_ _01503_ _02359_ _04183_ vssd1 vssd1 vccd1 vccd1 _04207_ sky130_fd_sc_hd__o21a_1
XANTENNA__10764__S net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06345_ net896 _01479_ _01485_ vssd1 vssd1 vccd1 vccd1 _01487_ sky130_fd_sc_hd__nor3_1
XFILLER_0_97_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout220_A _04766_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_220 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout318_A _02830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07978__A2 net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09064_ _04136_ _04137_ _04138_ vssd1 vssd1 vccd1 vccd1 _04139_ sky130_fd_sc_hd__or3_1
XFILLER_0_4_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06276_ top.lcd.cnt_500hz\[11\] _01438_ vssd1 vssd1 vccd1 vccd1 _01439_ sky130_fd_sc_hd__nand2_1
XFILLER_0_114_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08015_ _03149_ _03148_ vssd1 vssd1 vccd1 vccd1 _03154_ sky130_fd_sc_hd__and2b_1
XFILLER_0_102_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_116_2185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold620 top.DUT.register\[17\]\[9\] vssd1 vssd1 vccd1 vccd1 net1736 sky130_fd_sc_hd__dlygate4sd3_1
Xhold631 top.DUT.register\[27\]\[6\] vssd1 vssd1 vccd1 vccd1 net1747 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06262__B net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold642 top.DUT.register\[23\]\[19\] vssd1 vssd1 vccd1 vccd1 net1758 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08927__A1 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12184__B1 net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold653 top.DUT.register\[28\]\[2\] vssd1 vssd1 vccd1 vccd1 net1769 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold664 top.DUT.register\[14\]\[31\] vssd1 vssd1 vccd1 vccd1 net1780 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06938__B1 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold675 top.DUT.register\[18\]\[12\] vssd1 vssd1 vccd1 vccd1 net1791 sky130_fd_sc_hd__dlygate4sd3_1
Xhold686 top.DUT.register\[24\]\[13\] vssd1 vssd1 vccd1 vccd1 net1802 sky130_fd_sc_hd__dlygate4sd3_1
Xhold697 top.DUT.register\[12\]\[6\] vssd1 vssd1 vccd1 vccd1 net1813 sky130_fd_sc_hd__dlygate4sd3_1
X_09966_ net2280 net192 net630 vssd1 vssd1 vccd1 vccd1 _00174_ sky130_fd_sc_hd__mux2_1
XANTENNA__09573__B _04620_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08917_ net425 _04022_ _04025_ _04015_ vssd1 vssd1 vccd1 vccd1 _04026_ sky130_fd_sc_hd__a211o_1
XFILLER_0_85_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09897_ _04903_ _04905_ net490 _04896_ vssd1 vssd1 vccd1 vccd1 _04906_ sky130_fd_sc_hd__o211a_2
XANTENNA_fanout854_A net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_96_clk clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_96_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout475_X net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08848_ net324 _03631_ _03959_ vssd1 vssd1 vccd1 vccd1 _03960_ sky130_fd_sc_hd__o21a_1
XANTENNA__10004__S net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_1_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10939__S net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08779_ _01920_ _03893_ vssd1 vssd1 vccd1 vccd1 _03894_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout642_X net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_196_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10810_ net204 net2243 net600 vssd1 vssd1 vccd1 vccd1 _00971_ sky130_fd_sc_hd__mux2_1
X_11790_ _05668_ _05672_ vssd1 vssd1 vccd1 vccd1 _05673_ sky130_fd_sc_hd__nand2_1
XANTENNA__07115__B1 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_45_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07666__A1 top.a1.instruction\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10741_ net1757 net208 net419 vssd1 vssd1 vccd1 vccd1 _00902_ sky130_fd_sc_hd__mux2_1
XANTENNA__07666__B2 top.a1.instruction\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06437__B net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13460_ clknet_leaf_56_clk _01052_ net1074 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[30\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_165_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10672_ net2291 net228 net338 vssd1 vssd1 vccd1 vccd1 _00835_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_356 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12411_ clknet_leaf_109_clk top.ru.next_FetchedInstr\[23\] net975 vssd1 vssd1 vccd1
+ vccd1 top.a1.instruction\[23\] sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_11_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08615__B1 _03737_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13391_ clknet_leaf_32_clk _00983_ net1024 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[27\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_63_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10674__S net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_20_clk clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_20_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__07969__A2 net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12342_ _06137_ net791 _06136_ vssd1 vssd1 vccd1 vccd1 _01367_ sky130_fd_sc_hd__and3b_1
XANTENNA__06453__A top.a1.instruction\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10973__A1 top.a1.dataIn\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_584 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06641__A2 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12273_ _06094_ net686 _06093_ vssd1 vssd1 vccd1 vccd1 _01341_ sky130_fd_sc_hd__and3b_1
X_11224_ top.lcd.nextState\[3\] top.lcd.nextState\[4\] vssd1 vssd1 vccd1 vccd1 _05117_
+ sky130_fd_sc_hd__and2b_1
XANTENNA__10262__X _04978_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11155_ net844 _05084_ vssd1 vssd1 vccd1 vccd1 _05085_ sky130_fd_sc_hd__and2b_2
X_10106_ net1504 net166 net614 vssd1 vssd1 vccd1 vccd1 _00307_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_147_2646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11086_ net908 net1572 net863 _05048_ vssd1 vssd1 vccd1 vccd1 _01194_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_147_2657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08099__B net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_87_clk clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_87_clk
+ sky130_fd_sc_hd__clkbuf_8
X_10037_ net2034 net176 net622 vssd1 vssd1 vccd1 vccd1 _00240_ sky130_fd_sc_hd__mux2_1
XANTENNA__07354__B1 net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_160_2846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10849__S net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_172_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_188_768 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11534__A top.a1.dataIn\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_203_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11988_ _05870_ vssd1 vssd1 vccd1 vccd1 _05871_ sky130_fd_sc_hd__inv_2
XANTENNA__07106__B1 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_193_3334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11253__B top.lcd.nextState\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13727_ clknet_leaf_90_clk _01298_ net1005 vssd1 vssd1 vccd1 vccd1 top.a1.row2\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_10939_ net1577 net186 net592 vssd1 vssd1 vccd1 vccd1 _01100_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_193_3345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13658_ clknet_leaf_90_clk _01234_ net998 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[104\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_30_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_171_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12609_ clknet_leaf_15_clk _00201_ net961 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[3\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10584__S net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06880__A2 net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13589_ clknet_leaf_46_clk net1206 net1090 vssd1 vssd1 vccd1 vccd1 net80 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_143_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_11_clk clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_11_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_205_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_197_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06632__A2 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08909__A1 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09674__A top.a1.instruction\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout407 _04716_ vssd1 vssd1 vccd1 vccd1 net407 sky130_fd_sc_hd__clkbuf_4
X_09820_ _04834_ _04835_ vssd1 vssd1 vccd1 vccd1 _04836_ sky130_fd_sc_hd__nor2_1
Xfanout418 net421 vssd1 vssd1 vccd1 vccd1 net418 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_39_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout429 net430 vssd1 vssd1 vccd1 vccd1 net429 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07593__B1 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09751_ _04772_ _04773_ vssd1 vssd1 vccd1 vccd1 _04774_ sky130_fd_sc_hd__nor2_1
X_06963_ top.DUT.register\[15\]\[23\] net681 net677 top.DUT.register\[31\]\[23\] vssd1
+ vssd1 vccd1 vccd1 _02102_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_78_clk clknet_4_12__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_78_clk
+ sky130_fd_sc_hd__clkbuf_8
X_08702_ net277 _03773_ _03820_ vssd1 vssd1 vccd1 vccd1 _03821_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09680__Y _04716_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09682_ top.a1.instruction\[7\] top.a1.instruction\[8\] net786 vssd1 vssd1 vccd1
+ vccd1 _04718_ sky130_fd_sc_hd__o21ai_1
X_06894_ top.DUT.register\[24\]\[18\] net645 net720 top.DUT.register\[19\]\[18\] _02032_
+ vssd1 vssd1 vccd1 vccd1 _02033_ sky130_fd_sc_hd__a221o_1
XANTENNA__07345__B1 net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_146_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08633_ _03271_ _03310_ vssd1 vssd1 vccd1 vccd1 _03755_ sky130_fd_sc_hd__nand2_1
XANTENNA__07922__A _02498_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08665__A1_N _03334_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06699__A2 net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10759__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11444__A top.a1.dataIn\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_571 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout268_A _04726_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08564_ _03688_ vssd1 vssd1 vccd1 vccd1 _03689_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07515_ _02633_ _02653_ vssd1 vssd1 vccd1 vccd1 _02654_ sky130_fd_sc_hd__nor2_1
X_08495_ _03621_ _03622_ vssd1 vssd1 vccd1 vccd1 _03623_ sky130_fd_sc_hd__nor2_2
XANTENNA_fanout435_A net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06257__B net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09849__A top.pc\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07446_ top.DUT.register\[29\]\[15\] net452 net444 top.DUT.register\[1\]\[15\] vssd1
+ vssd1 vccd1 vccd1 _02585_ sky130_fd_sc_hd__a22o_1
XFILLER_0_119_367 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_2214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10494__S net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06871__A2 net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout602_A _04957_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07377_ top.DUT.register\[25\]\[8\] net779 net723 top.DUT.register\[29\]\[8\] vssd1
+ vssd1 vccd1 vccd1 _02516_ sky130_fd_sc_hd__a22o_1
XFILLER_0_91_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_40_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09116_ _02952_ _02994_ vssd1 vssd1 vccd1 vccd1 _04191_ sky130_fd_sc_hd__nand2_1
XFILLER_0_32_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06328_ _01390_ _01474_ vssd1 vssd1 vccd1 vccd1 _01475_ sky130_fd_sc_hd__nand2_2
XFILLER_0_161_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_2414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06623__A2 net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09047_ net281 _03471_ _03644_ net320 net271 vssd1 vssd1 vccd1 vccd1 _04122_ sky130_fd_sc_hd__o221a_1
X_06259_ top.ramload\[20\] net853 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedData\[20\]
+ sky130_fd_sc_hd__and2_1
Xhold450 top.DUT.register\[31\]\[20\] vssd1 vssd1 vccd1 vccd1 net1566 sky130_fd_sc_hd__dlygate4sd3_1
Xhold461 top.DUT.register\[31\]\[19\] vssd1 vssd1 vccd1 vccd1 net1577 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout592_X net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout971_A net1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold472 top.DUT.register\[19\]\[14\] vssd1 vssd1 vccd1 vccd1 net1588 sky130_fd_sc_hd__dlygate4sd3_1
Xhold483 top.DUT.register\[14\]\[16\] vssd1 vssd1 vccd1 vccd1 net1599 sky130_fd_sc_hd__dlygate4sd3_1
Xhold494 top.DUT.register\[3\]\[22\] vssd1 vssd1 vccd1 vccd1 net1610 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout930 net931 vssd1 vssd1 vccd1 vccd1 net930 sky130_fd_sc_hd__clkbuf_4
Xfanout941 net943 vssd1 vssd1 vccd1 vccd1 net941 sky130_fd_sc_hd__buf_2
Xfanout952 net967 vssd1 vssd1 vccd1 vccd1 net952 sky130_fd_sc_hd__clkbuf_2
X_09949_ net1478 net255 net629 vssd1 vssd1 vccd1 vccd1 _00157_ sky130_fd_sc_hd__mux2_1
Xfanout963 net964 vssd1 vssd1 vccd1 vccd1 net963 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_205_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_69_clk clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_69_clk
+ sky130_fd_sc_hd__clkbuf_8
Xfanout974 net1007 vssd1 vssd1 vccd1 vccd1 net974 sky130_fd_sc_hd__buf_2
XANTENNA__12511__Q top.pc\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout985 net986 vssd1 vssd1 vccd1 vccd1 net985 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_129_2376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout996 net997 vssd1 vssd1 vccd1 vccd1 net996 sky130_fd_sc_hd__clkbuf_4
X_12960_ clknet_leaf_17_clk _00552_ net965 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[14\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_129_2387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1150 top.DUT.register\[30\]\[20\] vssd1 vssd1 vccd1 vccd1 net2266 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1161 top.DUT.register\[30\]\[27\] vssd1 vssd1 vccd1 vccd1 net2277 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11911_ _05792_ _05793_ vssd1 vssd1 vccd1 vccd1 _05794_ sky130_fd_sc_hd__nand2_1
Xhold1172 top.DUT.register\[10\]\[9\] vssd1 vssd1 vccd1 vccd1 net2288 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1183 top.DUT.register\[14\]\[27\] vssd1 vssd1 vccd1 vccd1 net2299 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10669__S net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12891_ clknet_leaf_125_clk _00483_ net923 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[12\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1194 top.DUT.register\[27\]\[10\] vssd1 vssd1 vccd1 vccd1 net2310 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11842_ _05698_ _05724_ vssd1 vssd1 vccd1 vccd1 _05725_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_142_2576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09628__A2 _04657_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06448__A net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_185_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_200_547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11773_ _05616_ _05631_ vssd1 vssd1 vccd1 vccd1 _05656_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_138_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13512_ clknet_leaf_25_clk _01104_ net1009 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[31\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_10724_ net1674 net156 net336 vssd1 vssd1 vccd1 vccd1 _00885_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_175_3064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_175_3075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_193_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13443_ clknet_leaf_54_clk _01035_ net1038 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[29\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_22_clk_X clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10655_ net165 net2198 net345 vssd1 vssd1 vccd1 vccd1 _00819_ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_635 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkload17 clknet_leaf_123_clk vssd1 vssd1 vccd1 vccd1 clkload17/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_106_551 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13374_ clknet_leaf_54_clk _00966_ net1037 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[27\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload28 clknet_leaf_115_clk vssd1 vssd1 vccd1 vccd1 clkload28/Y sky130_fd_sc_hd__clkinv_2
X_10586_ net1374 net177 net351 vssd1 vssd1 vccd1 vccd1 _00752_ sky130_fd_sc_hd__mux2_1
Xclkload39 clknet_leaf_96_clk vssd1 vssd1 vccd1 vccd1 clkload39/Y sky130_fd_sc_hd__bufinv_16
XTAP_TAPCELL_ROW_58_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12325_ top.pad.button_control.r_counter\[9\] _06126_ vssd1 vssd1 vccd1 vccd1 _06127_
+ sky130_fd_sc_hd__and2_1
XANTENNA__06614__A2 net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06470__X _01609_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12256_ net1121 _06084_ net979 vssd1 vssd1 vccd1 vccd1 _06085_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_71_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11207_ net845 _05022_ _05034_ vssd1 vssd1 vccd1 vccd1 _05110_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_71_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09564__B2 _04051_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12187_ top.a1.row2\[42\] net847 net797 net131 vssd1 vssd1 vccd1 vccd1 _01295_ sky130_fd_sc_hd__a22o_1
XFILLER_0_76_49 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07575__B1 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_207_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11138_ net906 net1305 net861 _05074_ vssd1 vssd1 vccd1 vccd1 _01220_ sky130_fd_sc_hd__a31o_1
X_11069_ net85 net870 net834 net1166 vssd1 vssd1 vccd1 vccd1 _01180_ sky130_fd_sc_hd__a22o_1
XFILLER_0_92_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_0_clk clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_0_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_183_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10579__S net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_5__f_clk_X clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10960__C_N top.edg2.flip1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_703 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07300_ top.DUT.register\[12\]\[12\] net531 net515 top.DUT.register\[7\]\[12\] vssd1
+ vssd1 vccd1 vccd1 _02439_ sky130_fd_sc_hd__a22o_1
XFILLER_0_46_427 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_82_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08280_ net431 _03411_ _03413_ net495 _03415_ vssd1 vssd1 vccd1 vccd1 _03416_ sky130_fd_sc_hd__a221o_1
X_07231_ top.DUT.register\[22\]\[10\] net647 net758 top.DUT.register\[30\]\[10\] _02369_
+ vssd1 vssd1 vccd1 vccd1 _02370_ sky130_fd_sc_hd__a221o_1
XFILLER_0_73_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_123 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07162_ top.DUT.register\[4\]\[11\] net667 net754 top.DUT.register\[1\]\[11\] _02300_
+ vssd1 vssd1 vccd1 vccd1 _02301_ sky130_fd_sc_hd__a221o_1
XFILLER_0_144_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07093_ _02225_ _02227_ _02229_ _02231_ vssd1 vssd1 vccd1 vccd1 _02232_ sky130_fd_sc_hd__or4_4
XTAP_TAPCELL_ROW_113_2144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06380__X _01519_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13433__RESET_B net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout204 net206 vssd1 vssd1 vccd1 vccd1 net204 sky130_fd_sc_hd__buf_2
Xfanout215 net218 vssd1 vssd1 vccd1 vccd1 net215 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07566__B1 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout226 _04805_ vssd1 vssd1 vccd1 vccd1 net226 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout237 _04757_ vssd1 vssd1 vccd1 vccd1 net237 sky130_fd_sc_hd__clkbuf_2
X_09803_ _04819_ _04820_ vssd1 vssd1 vccd1 vccd1 _04821_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09691__X _04726_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07030__A2 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout248 _04749_ vssd1 vssd1 vccd1 vccd1 net248 sky130_fd_sc_hd__buf_1
Xfanout259 net262 vssd1 vssd1 vccd1 vccd1 net259 sky130_fd_sc_hd__clkbuf_2
X_07995_ top.DUT.register\[22\]\[31\] net649 net760 top.DUT.register\[30\]\[31\] _03130_
+ vssd1 vssd1 vccd1 vccd1 _03134_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout385_A _04978_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09734_ net2265 net232 net631 vssd1 vssd1 vccd1 vccd1 _00130_ sky130_fd_sc_hd__mux2_1
X_06946_ top.DUT.register\[25\]\[21\] net781 net748 top.DUT.register\[17\]\[21\] vssd1
+ vssd1 vccd1 vccd1 _02085_ sky130_fd_sc_hd__a22o_1
XANTENNA__09851__B _01584_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07318__B1 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11114__A1 net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09665_ top.a1.halfData\[5\] _01471_ _04693_ net1086 vssd1 vssd1 vccd1 vccd1 _00119_
+ sky130_fd_sc_hd__o211a_1
XANTENNA__10489__S net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06877_ _02009_ _02011_ _02013_ _02015_ vssd1 vssd1 vccd1 vccd1 _02016_ sky130_fd_sc_hd__or4_2
XANTENNA_fanout552_A _01535_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06539__Y _01678_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08616_ _03121_ net426 vssd1 vssd1 vccd1 vccd1 _03739_ sky130_fd_sc_hd__nand2_1
XANTENNA__06268__A top.ramload\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12512__SET_B net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09596_ net902 top.pc\[30\] _04642_ net890 vssd1 vssd1 vccd1 vccd1 _00110_ sky130_fd_sc_hd__o211a_1
XFILLER_0_167_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12386__RESET_B net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08547_ _03470_ _03533_ _03670_ vssd1 vssd1 vccd1 vccd1 _03673_ sky130_fd_sc_hd__a21o_1
XFILLER_0_167_749 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout340_X net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout817_A _05044_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07097__A2 net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08294__A1 net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08478_ net434 _03606_ vssd1 vssd1 vccd1 vccd1 _03607_ sky130_fd_sc_hd__nor2_1
XFILLER_0_37_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09491__B1 _04543_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08294__B2 net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_484 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07429_ _02544_ _02567_ vssd1 vssd1 vccd1 vccd1 _02568_ sky130_fd_sc_hd__nand2_1
XFILLER_0_190_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout605_X net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10440_ net228 net1911 net365 vssd1 vssd1 vccd1 vccd1 _00611_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_21_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09794__A1 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10371_ net1753 net232 net373 vssd1 vssd1 vccd1 vccd1 _00546_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12110_ _05972_ _05978_ _05983_ _05992_ vssd1 vssd1 vccd1 vccd1 _05993_ sky130_fd_sc_hd__a22o_1
X_13090_ clknet_leaf_9_clk _00682_ net948 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[18\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_103_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09546__A1 net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12041_ _05913_ _05919_ vssd1 vssd1 vccd1 vccd1 _05924_ sky130_fd_sc_hd__nand2_1
Xhold280 top.DUT.register\[26\]\[5\] vssd1 vssd1 vccd1 vccd1 net1396 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold291 top.DUT.register\[25\]\[31\] vssd1 vssd1 vccd1 vccd1 net1407 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07557__B1 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07021__A2 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout760 _01617_ vssd1 vssd1 vccd1 vccd1 net760 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_144_2605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout771 _01614_ vssd1 vssd1 vccd1 vccd1 net771 sky130_fd_sc_hd__clkbuf_4
Xfanout782 _01509_ vssd1 vssd1 vccd1 vccd1 net782 sky130_fd_sc_hd__buf_2
XANTENNA__08658__A _02047_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout793 net794 vssd1 vssd1 vccd1 vccd1 net793 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07309__B1 net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12943_ clknet_leaf_41_clk _00535_ net1056 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[13\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_64_clk_A clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_177_3104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12874_ clknet_leaf_117_clk _00466_ net958 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[11\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_62_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_29_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_158_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11825_ _05673_ _05675_ net131 vssd1 vssd1 vccd1 vccd1 _05708_ sky130_fd_sc_hd__nand3_1
XANTENNA__08809__B1 net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09489__A net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11756_ _05597_ _05620_ vssd1 vssd1 vccd1 vccd1 _05639_ sky130_fd_sc_hd__nand2_1
XANTENNA__07088__A2 net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_200_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_79_clk_A clknet_4_12__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10707_ net1778 net221 net334 vssd1 vssd1 vccd1 vccd1 _00868_ sky130_fd_sc_hd__mux2_1
XANTENNA__06835__A2 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11687_ _05529_ _05535_ _05549_ vssd1 vssd1 vccd1 vccd1 _05570_ sky130_fd_sc_hd__o21a_1
XFILLER_0_55_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_122_clk_A clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06625__B _01763_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_155_2767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13426_ clknet_leaf_23_clk _01018_ net1014 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[29\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_155_2778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10638_ net231 net2192 net342 vssd1 vssd1 vccd1 vccd1 _00802_ sky130_fd_sc_hd__mux2_1
XANTENNA__11250__C _05130_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload106 clknet_leaf_63_clk vssd1 vssd1 vccd1 vccd1 clkload106/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_181_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_307 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_430 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08588__A2 net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13357_ clknet_leaf_41_clk _00949_ net1057 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[26\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10862__S net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10569_ net1881 net243 net350 vssd1 vssd1 vccd1 vccd1 _00735_ sky130_fd_sc_hd__mux2_1
XANTENNA__09936__B _04644_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07796__B1 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12308_ top.pad.button_control.r_counter\[3\] _06114_ vssd1 vssd1 vccd1 vccd1 _06116_
+ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_188_3266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13288_ clknet_leaf_7_clk _00880_ net946 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[24\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11259__A _05121_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12239_ _06074_ net978 _06073_ vssd1 vssd1 vccd1 vccd1 _01321_ sky130_fd_sc_hd__and3b_1
XANTENNA__07548__B1 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_17_clk_A clknet_4_12__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_194_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07012__A2 net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12897__RESET_B net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_207_3550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06800_ _01932_ _01934_ _01936_ _01938_ vssd1 vssd1 vccd1 vccd1 _01939_ sky130_fd_sc_hd__or4_4
X_07780_ top.DUT.register\[12\]\[2\] net738 net714 top.DUT.register\[27\]\[2\] _02918_
+ vssd1 vssd1 vccd1 vccd1 _02919_ sky130_fd_sc_hd__a221o_1
Xinput4 DAT_I[11] vssd1 vssd1 vccd1 vccd1 net4 sky130_fd_sc_hd__clkbuf_1
XANTENNA__07472__A _02590_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06731_ top.DUT.register\[30\]\[25\] net758 net730 top.DUT.register\[14\]\[25\] _01869_
+ vssd1 vssd1 vccd1 vccd1 _01870_ sky130_fd_sc_hd__a221o_1
XFILLER_0_189_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08512__A2 net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09450_ net901 top.pc\[21\] _04505_ net891 vssd1 vssd1 vccd1 vccd1 _00101_ sky130_fd_sc_hd__o211a_1
X_06662_ top.DUT.register\[10\]\[26\] net521 _01800_ vssd1 vssd1 vccd1 vccd1 _01801_
+ sky130_fd_sc_hd__a21o_1
XANTENNA__10102__S net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07720__B1 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_203_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08401_ net324 net316 vssd1 vssd1 vccd1 vccd1 _03533_ sky130_fd_sc_hd__nor2_1
XFILLER_0_188_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12813__CLK clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09381_ _01930_ _01939_ _04438_ vssd1 vssd1 vccd1 vccd1 _04441_ sky130_fd_sc_hd__or3_1
X_06593_ top.DUT.register\[10\]\[28\] net773 net717 top.DUT.register\[27\]\[28\] _01728_
+ vssd1 vssd1 vccd1 vccd1 _01732_ sky130_fd_sc_hd__a221o_1
XANTENNA__08971__A2_N net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08332_ net280 _03464_ _03465_ net283 vssd1 vssd1 vccd1 vccd1 _03466_ sky130_fd_sc_hd__o22a_1
XFILLER_0_191_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06375__X _01514_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06287__B1 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08263_ net276 _03287_ vssd1 vssd1 vccd1 vccd1 _03399_ sky130_fd_sc_hd__nor2_1
XANTENNA__06826__A2 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_646 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout133_A net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07214_ _01485_ _01588_ _02346_ _01475_ _02338_ vssd1 vssd1 vccd1 vccd1 _02353_ sky130_fd_sc_hd__o221a_1
XPHY_EDGE_ROW_104_Left_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08194_ net307 _03331_ vssd1 vssd1 vccd1 vccd1 _03332_ sky130_fd_sc_hd__nor2_1
XFILLER_0_6_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09225__B1 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07145_ top.DUT.register\[28\]\[11\] net555 net451 top.DUT.register\[29\]\[11\] _02283_
+ vssd1 vssd1 vccd1 vccd1 _02284_ sky130_fd_sc_hd__a221o_1
XANTENNA__10772__S net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07787__B1 net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_1869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07076_ top.DUT.register\[4\]\[22\] net668 net734 top.DUT.register\[16\]\[22\] _02209_
+ vssd1 vssd1 vccd1 vccd1 _02215_ sky130_fd_sc_hd__a221o_1
XFILLER_0_112_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06270__B net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_7_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07003__A2 net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout767_A net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout388_X net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_113_Left_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_199_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07978_ top.DUT.register\[9\]\[31\] net468 net465 top.DUT.register\[13\]\[31\] _03116_
+ vssd1 vssd1 vccd1 vccd1 _03117_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_126_2335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08478__A net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09717_ net829 _04270_ vssd1 vssd1 vccd1 vccd1 _04746_ sky130_fd_sc_hd__nor2_1
X_06929_ _02061_ _02063_ _02065_ _02067_ vssd1 vssd1 vccd1 vccd1 _02068_ sky130_fd_sc_hd__or4_2
XFILLER_0_97_603 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout934_A net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout555_X net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09700__A1 _03430_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09648_ _04675_ _04689_ vssd1 vssd1 vccd1 vccd1 _04690_ sky130_fd_sc_hd__nor2_1
XFILLER_0_195_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_179_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_167_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_26_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10947__S net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout722_X net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09579_ _04624_ _04626_ top.pc\[29\] _04051_ vssd1 vssd1 vccd1 vccd1 _00109_ sky130_fd_sc_hd__o2bb2a_1
X_11610_ _05467_ _05482_ vssd1 vssd1 vccd1 vccd1 _05493_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_194_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_182_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12590_ clknet_leaf_39_clk _00182_ net1054 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[2\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_65_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_172_3023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_624 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11541_ _05364_ _05399_ _05422_ _05423_ vssd1 vssd1 vccd1 vccd1 _05424_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__11271__B1 _05136_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_122_Left_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06817__A2 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xwire413 _02088_ vssd1 vssd1 vccd1 vccd1 net413 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_9_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11472_ _05321_ _05322_ _05350_ vssd1 vssd1 vccd1 vccd1 _05355_ sky130_fd_sc_hd__and3_1
XFILLER_0_163_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07490__A2 net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13211_ clknet_leaf_125_clk _00803_ net924 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[22\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_137_2497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10423_ net1344 net166 net371 vssd1 vssd1 vccd1 vccd1 _00595_ sky130_fd_sc_hd__mux2_1
XANTENNA__10682__S net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07778__B1 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13142_ clknet_leaf_4_clk _00734_ net940 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[20\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07242__A2 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10354_ net1744 net168 net380 vssd1 vssd1 vccd1 vccd1 _00530_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_150_2697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13073_ clknet_leaf_116_clk _00665_ net988 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[18\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_10285_ net1908 net181 net385 vssd1 vssd1 vccd1 vccd1 _00463_ sky130_fd_sc_hd__mux2_1
X_12024_ _05886_ _05904_ vssd1 vssd1 vccd1 vccd1 _05907_ sky130_fd_sc_hd__xor2_1
XPHY_EDGE_ROW_131_Left_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_168_Right_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_183_3185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_183_3196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07292__A _02409_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_205_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12926_ clknet_leaf_20_clk _00518_ net1029 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[13\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_186_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_66_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_202_3480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09711__S net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10857__S net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12857_ clknet_leaf_10_clk _00449_ net949 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[11\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_158_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_157_2807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12986__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_680 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_708 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11808_ _05659_ _05668_ _05690_ vssd1 vssd1 vccd1 vccd1 _05691_ sky130_fd_sc_hd__nand3_4
XFILLER_0_56_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_140_Left_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_173_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12788_ clknet_leaf_55_clk _00380_ net1073 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[9\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_173_538 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11739_ _05589_ _05620_ vssd1 vssd1 vccd1 vccd1 _05622_ sky130_fd_sc_hd__and2_2
XANTENNA__06808__A2 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_89 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07481__A2 net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11014__B1 _05044_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10592__S net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13409_ clknet_leaf_18_clk _01001_ net1027 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[28\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07769__B1 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07233__A2 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_110_2103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08950_ net1267 net873 _02748_ net693 vssd1 vssd1 vccd1 vccd1 _00056_ sky130_fd_sc_hd__a22o_1
X_07901_ _03030_ _03039_ vssd1 vssd1 vccd1 vccd1 _03040_ sky130_fd_sc_hd__nor2_8
XTAP_TAPCELL_ROW_168_2969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08881_ net1305 net830 net800 _03991_ vssd1 vssd1 vccd1 vccd1 _00046_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_4_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_135_Right_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07832_ top.DUT.register\[16\]\[0\] net737 _02968_ _02970_ vssd1 vssd1 vccd1 vccd1
+ _02971_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_90_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07763_ net820 _02901_ _02359_ vssd1 vssd1 vccd1 vccd1 _02902_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_108_2065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09502_ _04551_ _04552_ vssd1 vssd1 vccd1 vccd1 _04554_ sky130_fd_sc_hd__nor2_1
XFILLER_0_2_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06714_ _01843_ _01852_ vssd1 vssd1 vccd1 vccd1 _01853_ sky130_fd_sc_hd__nor2_4
XFILLER_0_78_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_189_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07694_ top.DUT.register\[20\]\[4\] net565 net505 top.DUT.register\[27\]\[4\] vssd1
+ vssd1 vccd1 vccd1 _02833_ sky130_fd_sc_hd__a22o_1
XANTENNA__11096__A3 net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09694__B1 net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_524 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09433_ _04472_ _04489_ _04488_ vssd1 vssd1 vccd1 vccd1 _04490_ sky130_fd_sc_hd__a21oi_1
X_06645_ net808 _01783_ net437 vssd1 vssd1 vccd1 vccd1 _01784_ sky130_fd_sc_hd__o21a_1
XANTENNA__10767__S net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_2254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_2265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08745__B net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout348_A _04991_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09364_ _04423_ _04424_ vssd1 vssd1 vccd1 vccd1 _04425_ sky130_fd_sc_hd__xnor2_1
XANTENNA__08249__A1 net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06576_ top.DUT.register\[7\]\[28\] net518 net442 top.DUT.register\[5\]\[28\] _01714_
+ vssd1 vssd1 vccd1 vccd1 _01715_ sky130_fd_sc_hd__a221o_1
XFILLER_0_59_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08249__B2 _03334_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08315_ _03449_ vssd1 vssd1 vccd1 vccd1 _03450_ sky130_fd_sc_hd__inv_2
XFILLER_0_170_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_164_549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09295_ net897 top.pc\[12\] _04359_ net889 vssd1 vssd1 vccd1 vccd1 _00092_ sky130_fd_sc_hd__o211a_1
XFILLER_0_145_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout515_A _01558_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout136_X net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06265__B net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09857__A top.pc\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08246_ _02945_ net499 net494 _02947_ _03382_ vssd1 vssd1 vccd1 vccd1 _03383_ sky130_fd_sc_hd__a221o_1
XANTENNA__06680__B1 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08177_ _01722_ net329 vssd1 vssd1 vccd1 vccd1 _03315_ sky130_fd_sc_hd__nand2_1
XFILLER_0_6_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07128_ _02050_ _02223_ _02266_ vssd1 vssd1 vccd1 vccd1 _02267_ sky130_fd_sc_hd__nand3b_1
XTAP_TAPCELL_ROW_37_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout884_A net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13291__CLK clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10007__S net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07059_ _02188_ _02197_ vssd1 vssd1 vccd1 vccd1 _02198_ sky130_fd_sc_hd__nor2_8
XFILLER_0_100_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12748__RESET_B net1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10070_ net1657 net178 net617 vssd1 vssd1 vccd1 vccd1 _00272_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout672_X net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_102_Right_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10195__A_N net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13760_ clknet_leaf_71_clk _01331_ vssd1 vssd1 vccd1 vccd1 top.lcd.currentState\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_168_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10972_ top.a1.halfData\[2\] _04667_ _05012_ net843 vssd1 vssd1 vccd1 vccd1 _05013_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__08488__A1 net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09685__B1 net34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08488__B2 _03334_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12711_ clknet_leaf_6_clk _00303_ net937 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[6\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10677__S net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13691_ clknet_leaf_70_clk _00003_ vssd1 vssd1 vccd1 vccd1 top.lcd.nextState\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_48_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12642_ clknet_leaf_10_clk _00234_ net949 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[4\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06456__A top.a1.instruction\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_139_2526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_566 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_139_2537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11244__B1 _05136_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12573_ clknet_leaf_119_clk _00165_ net953 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[2\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_182_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08942__Y _04049_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07999__B1 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_519 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11524_ _05406_ vssd1 vssd1 vccd1 vccd1 _05407_ sky130_fd_sc_hd__inv_2
XFILLER_0_80_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08660__A1 _02049_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07463__A2 net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_262 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08660__B2 _03258_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_152_2726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11455_ _05305_ _05336_ vssd1 vssd1 vccd1 vccd1 _05338_ sky130_fd_sc_hd__xnor2_2
XANTENNA__09486__B _01584_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10406_ net1661 net232 net369 vssd1 vssd1 vccd1 vccd1 _00578_ sky130_fd_sc_hd__mux2_1
XANTENNA__08412__A1 net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_150_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11386_ _05249_ _05250_ _05236_ _05242_ _05244_ vssd1 vssd1 vccd1 vccd1 _05269_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_1_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_185_3214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_185_3225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13125_ clknet_leaf_35_clk _00717_ net1041 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[19\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10337_ net1738 net238 net377 vssd1 vssd1 vccd1 vccd1 _00513_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_488 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09706__S net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13056_ clknet_leaf_114_clk _00648_ net964 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[17\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_10268_ net1649 net251 net385 vssd1 vssd1 vccd1 vccd1 _00446_ sky130_fd_sc_hd__mux2_1
XANTENNA__12418__RESET_B net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12007_ _05865_ _05866_ _05870_ net126 _05869_ vssd1 vssd1 vccd1 vccd1 _05890_ sky130_fd_sc_hd__a41o_1
XFILLER_0_84_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_206_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10199_ net263 net2118 net393 vssd1 vssd1 vccd1 vccd1 _00379_ sky130_fd_sc_hd__mux2_1
XFILLER_0_206_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11256__B _05130_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_163_2888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_200_3439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12909_ clknet_leaf_41_clk _00501_ net1057 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[12\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10587__S net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_201_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_196_3387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06430_ top.DUT.register\[1\]\[30\] net445 net509 top.DUT.register\[4\]\[30\] _01568_
+ vssd1 vssd1 vccd1 vccd1 _01569_ sky130_fd_sc_hd__a221o_1
XFILLER_0_158_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_174_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_376 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06361_ net896 _01473_ vssd1 vssd1 vccd1 vccd1 _01500_ sky130_fd_sc_hd__and2_2
XFILLER_0_44_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_139_590 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08100_ net325 net315 vssd1 vssd1 vccd1 vccd1 _03239_ sky130_fd_sc_hd__nand2_1
X_09080_ top.a1.instruction\[7\] top.a1.instruction\[8\] vssd1 vssd1 vccd1 vccd1 _04155_
+ sky130_fd_sc_hd__and2_2
XFILLER_0_16_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07454__A2 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06292_ net882 net815 net813 top.lcd.currentState\[1\] net1084 vssd1 vssd1 vccd1
+ vccd1 _01330_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_79_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08031_ net319 net315 vssd1 vssd1 vccd1 vccd1 _03170_ sky130_fd_sc_hd__nor2_2
XPHY_EDGE_ROW_204_Right_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09396__B _02025_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold802 top.DUT.register\[22\]\[17\] vssd1 vssd1 vccd1 vccd1 net1918 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold813 top.DUT.register\[21\]\[20\] vssd1 vssd1 vccd1 vccd1 net1929 sky130_fd_sc_hd__dlygate4sd3_1
Xhold824 top.DUT.register\[9\]\[19\] vssd1 vssd1 vccd1 vccd1 net1940 sky130_fd_sc_hd__dlygate4sd3_1
Xhold835 top.DUT.register\[18\]\[5\] vssd1 vssd1 vccd1 vccd1 net1951 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09600__B1 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold846 top.DUT.register\[22\]\[20\] vssd1 vssd1 vccd1 vccd1 net1962 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_1828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold857 top.DUT.register\[7\]\[21\] vssd1 vssd1 vccd1 vccd1 net1973 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08954__A2 net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09982_ net265 net1752 net623 vssd1 vssd1 vccd1 vccd1 _00187_ sky130_fd_sc_hd__mux2_1
Xhold868 top.DUT.register\[9\]\[1\] vssd1 vssd1 vccd1 vccd1 net1984 sky130_fd_sc_hd__dlygate4sd3_1
Xhold879 top.a1.row1\[111\] vssd1 vssd1 vccd1 vccd1 net1995 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07484__X _02623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08933_ net281 _03529_ vssd1 vssd1 vccd1 vccd1 _04041_ sky130_fd_sc_hd__nor2_2
XFILLER_0_110_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07925__A _02453_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08864_ _01745_ _03974_ vssd1 vssd1 vccd1 vccd1 _03975_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout1005_A net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07815_ top.DUT.register\[10\]\[0\] net770 net750 top.DUT.register\[26\]\[0\] vssd1
+ vssd1 vccd1 vccd1 _02954_ sky130_fd_sc_hd__a22o_1
X_08795_ _03909_ vssd1 vssd1 vccd1 vccd1 _03910_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout465_A net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07746_ top.DUT.register\[13\]\[3\] net465 net538 top.DUT.register\[19\]\[3\] vssd1
+ vssd1 vccd1 vccd1 _02885_ sky130_fd_sc_hd__a22o_1
XFILLER_0_211_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09131__A2 net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07660__A _02798_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10497__S net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07677_ top.DUT.register\[7\]\[4\] net660 net772 top.DUT.register\[10\]\[4\] vssd1
+ vssd1 vccd1 vccd1 _02816_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout632_A _04714_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09416_ _04472_ _04473_ vssd1 vssd1 vccd1 vccd1 _04474_ sky130_fd_sc_hd__nand2_1
X_06628_ top.DUT.register\[5\]\[27\] net654 net638 top.DUT.register\[6\]\[27\] _01766_
+ vssd1 vssd1 vccd1 vccd1 _01767_ sky130_fd_sc_hd__a221o_1
XFILLER_0_164_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_36_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07693__A2 net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10029__A1 net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09347_ net136 _04395_ _04408_ net899 vssd1 vssd1 vccd1 vccd1 _04409_ sky130_fd_sc_hd__o211ai_1
X_06559_ net808 _01697_ net438 vssd1 vssd1 vccd1 vccd1 _01698_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout420_X net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_1957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_1968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout518_X net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_240 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07659__X _02798_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_700 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09278_ net136 _04328_ _04343_ vssd1 vssd1 vccd1 vccd1 _04344_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07445__A2 net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08642__B2 net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08229_ _03364_ _03365_ net311 vssd1 vssd1 vccd1 vccd1 _03366_ sky130_fd_sc_hd__mux2_1
XANTENNA__06653__B1 net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_232 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_2456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_539 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11240_ top.lcd.nextState\[3\] net878 vssd1 vssd1 vccd1 vccd1 _05133_ sky130_fd_sc_hd__nor2_1
XANTENNA__09874__X _04885_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12681__CLK clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06405__B1 net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12514__Q top.pc\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_630 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11171_ top.a1.halfData\[5\] _01415_ _01414_ top.a1.hexop\[3\] vssd1 vssd1 vccd1
+ vccd1 _05095_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_113_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_652 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10122_ net231 net2156 net607 vssd1 vssd1 vccd1 vccd1 _00322_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12511__RESET_B net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10053_ top.DUT.register\[5\]\[6\] net241 net615 vssd1 vssd1 vccd1 vccd1 _00255_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_180_3144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08002__Y _03141_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input26_A DAT_I[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08937__Y _04045_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13812_ net72 vssd1 vssd1 vccd1 vccd1 net109 sky130_fd_sc_hd__clkbuf_1
XANTENNA__06738__X _01877_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_203_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_199_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_786 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13743_ clknet_leaf_100_clk _01314_ vssd1 vssd1 vccd1 vccd1 top.lcd.cnt_20ms\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_10955_ _00016_ _01416_ vssd1 vssd1 vccd1 vccd1 _04998_ sky130_fd_sc_hd__nand2_1
XFILLER_0_97_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_211_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10200__S net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07684__A2 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13674_ clknet_leaf_92_clk _01250_ net998 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_10886_ net148 net2064 net596 vssd1 vssd1 vccd1 vccd1 _01047_ sky130_fd_sc_hd__mux2_1
XANTENNA__06892__B1 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12625_ clknet_leaf_112_clk _00217_ net988 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[4\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_14_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12556_ clknet_leaf_63_clk _00148_ net1090 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[1\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07436__A2 net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06473__X _01612_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11507_ _05388_ _05389_ vssd1 vssd1 vccd1 vccd1 _05390_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_13_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12487_ clknet_leaf_75_clk _00008_ net1077 vssd1 vssd1 vccd1 vccd1 top.a1.hexop\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_151_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold109 top.a1.data\[9\] vssd1 vssd1 vccd1 vccd1 net1225 sky130_fd_sc_hd__dlygate4sd3_1
X_11438_ _05286_ _05320_ vssd1 vssd1 vccd1 vccd1 _05321_ sky130_fd_sc_hd__nand2_1
XFILLER_0_123_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10870__S net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11369_ _05249_ _05250_ top.a1.dataIn\[19\] vssd1 vssd1 vccd1 vccd1 _05252_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09944__B _04712_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_210_3590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13108_ clknet_leaf_55_clk _00700_ net1031 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[19\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_165_2917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_165_2928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13039_ clknet_leaf_32_clk _00631_ net1024 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[16\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_119_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09897__B1 net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_198_3416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07600_ top.DUT.register\[28\]\[6\] net766 net710 top.DUT.register\[11\]\[6\] _02735_
+ vssd1 vssd1 vccd1 vccd1 _02739_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_105_2024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08580_ _03693_ _03698_ _03704_ vssd1 vssd1 vccd1 vccd1 _03705_ sky130_fd_sc_hd__or3b_2
XFILLER_0_178_438 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07531_ top.DUT.register\[7\]\[7\] net515 _02669_ vssd1 vssd1 vccd1 vccd1 _02670_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_49_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07462_ _02594_ _02597_ _02599_ _02600_ vssd1 vssd1 vccd1 vccd1 _02601_ sky130_fd_sc_hd__or4_1
XANTENNA__10110__S net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07675__A2 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09201_ net136 _04270_ vssd1 vssd1 vccd1 vccd1 _04271_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_33_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06413_ net684 _01523_ _01531_ vssd1 vssd1 vccd1 vccd1 _01552_ sky130_fd_sc_hd__and3_2
XANTENNA__06883__B1 net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07393_ top.DUT.register\[30\]\[9\] net579 net575 top.DUT.register\[22\]\[9\] vssd1
+ vssd1 vccd1 vccd1 _02532_ sky130_fd_sc_hd__a22o_1
XFILLER_0_72_631 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09132_ _01406_ _04051_ _04206_ vssd1 vssd1 vccd1 vccd1 _00082_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_8_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06344_ top.a1.instruction\[13\] top.a1.instruction\[14\] vssd1 vssd1 vccd1 vccd1
+ _01486_ sky130_fd_sc_hd__nand2_1
XFILLER_0_56_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06824__A _01940_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_506 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06635__B1 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09063_ _03410_ _03483_ _03501_ _03539_ vssd1 vssd1 vccd1 vccd1 _04138_ sky130_fd_sc_hd__or4b_1
X_06275_ top.lcd.cnt_500hz\[9\] top.lcd.cnt_500hz\[10\] vssd1 vssd1 vccd1 vccd1 _01438_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_114_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08014_ net894 _03148_ _02337_ _01477_ vssd1 vssd1 vccd1 vccd1 _03153_ sky130_fd_sc_hd__o211a_1
Xhold610 top.DUT.register\[12\]\[14\] vssd1 vssd1 vccd1 vccd1 net1726 sky130_fd_sc_hd__dlygate4sd3_1
Xhold621 top.DUT.register\[27\]\[24\] vssd1 vssd1 vccd1 vccd1 net1737 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_116_2186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12184__A1 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold632 top.DUT.register\[28\]\[29\] vssd1 vssd1 vccd1 vccd1 net1748 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_71 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold643 top.DUT.register\[26\]\[24\] vssd1 vssd1 vccd1 vccd1 net1759 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10780__S net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold654 top.DUT.register\[29\]\[6\] vssd1 vssd1 vccd1 vccd1 net1770 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold665 top.DUT.register\[31\]\[27\] vssd1 vssd1 vccd1 vccd1 net1781 sky130_fd_sc_hd__dlygate4sd3_1
Xhold676 top.DUT.register\[30\]\[18\] vssd1 vssd1 vccd1 vccd1 net1792 sky130_fd_sc_hd__dlygate4sd3_1
Xhold687 top.DUT.register\[3\]\[6\] vssd1 vssd1 vccd1 vccd1 net1803 sky130_fd_sc_hd__dlygate4sd3_1
Xhold698 top.DUT.register\[10\]\[15\] vssd1 vssd1 vccd1 vccd1 net1814 sky130_fd_sc_hd__dlygate4sd3_1
X_09965_ net1727 net202 net630 vssd1 vssd1 vccd1 vccd1 _00173_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout582_A _01514_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08916_ net436 _04020_ _04021_ _03259_ _04024_ vssd1 vssd1 vccd1 vccd1 _04025_ sky130_fd_sc_hd__a221o_1
XFILLER_0_176_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09896_ _04150_ _04901_ _04902_ _04904_ vssd1 vssd1 vccd1 vccd1 _04905_ sky130_fd_sc_hd__a31o_1
XANTENNA__09870__A top.pc\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08847_ net279 _03797_ _03958_ net282 vssd1 vssd1 vccd1 vccd1 _03959_ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout370_X net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout847_A net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout468_X net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08778_ _02134_ _02220_ _03892_ _02135_ vssd1 vssd1 vccd1 vccd1 _03893_ sky130_fd_sc_hd__a211o_1
X_07729_ _02863_ _02865_ _02867_ vssd1 vssd1 vccd1 vccd1 _02868_ sky130_fd_sc_hd__or3_1
XFILLER_0_192_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout635_X net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10020__S net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10740_ net2055 net211 net418 vssd1 vssd1 vccd1 vccd1 _00901_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_45_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_430 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06874__B1 net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10671_ net1583 net232 net338 vssd1 vssd1 vccd1 vccd1 _00834_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_11_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12410_ clknet_leaf_108_clk top.ru.next_FetchedInstr\[22\] net975 vssd1 vssd1 vccd1
+ vccd1 top.a1.instruction\[22\] sky130_fd_sc_hd__dfrtp_4
X_13390_ clknet_leaf_41_clk _00982_ net1057 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[27\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08615__A1 net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07418__A2 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_180_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_180_647 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_210 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12341_ top.pad.button_control.r_counter\[15\] top.pad.button_control.r_counter\[14\]
+ _06134_ vssd1 vssd1 vccd1 vccd1 _06137_ sky130_fd_sc_hd__and3_1
XANTENNA__06626__B1 net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12272_ top.lcd.cnt_500hz\[5\] top.lcd.cnt_500hz\[4\] top.lcd.cnt_500hz\[6\] _01436_
+ vssd1 vssd1 vccd1 vccd1 _06094_ sky130_fd_sc_hd__and4_1
XFILLER_0_133_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08918__A2 net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11223_ net1302 net472 vssd1 vssd1 vccd1 vccd1 _01263_ sky130_fd_sc_hd__nand2b_1
XANTENNA__10690__S net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07565__A _02703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11154_ _05002_ _05082_ vssd1 vssd1 vccd1 vccd1 _05084_ sky130_fd_sc_hd__nor2_1
XANTENNA__08013__X _03152_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10105_ net1391 net170 net611 vssd1 vssd1 vccd1 vccd1 _00306_ sky130_fd_sc_hd__mux2_1
X_11085_ net62 net864 vssd1 vssd1 vccd1 vccd1 _05048_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_147_2647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_147_2658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10036_ net2095 net182 net622 vssd1 vssd1 vccd1 vccd1 _00239_ sky130_fd_sc_hd__mux2_1
XANTENNA__11150__A2 net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08396__A net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_160_2847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06468__X _01607_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06909__A _02026_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11987_ _05839_ _05867_ vssd1 vssd1 vccd1 vccd1 _05870_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_85_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13726_ clknet_leaf_90_clk _01297_ net1002 vssd1 vssd1 vccd1 vccd1 top.a1.row2\[15\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_193_3335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10938_ net1336 net203 net591 vssd1 vssd1 vccd1 vccd1 _01099_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_193_3346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_430 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10865__S net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13657_ clknet_leaf_93_clk _00015_ net994 vssd1 vssd1 vccd1 vccd1 wb.curr_state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_10869_ net208 net2240 net596 vssd1 vssd1 vccd1 vccd1 _01030_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_30_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07409__A2 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12608_ clknet_leaf_114_clk _00200_ net964 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[3\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_13588_ clknet_leaf_89_clk net1189 net1002 vssd1 vssd1 vccd1 vccd1 net79 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06617__B1 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12539_ clknet_leaf_124_clk _00131_ net923 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[1\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_30_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07290__B1 net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07042__B1 net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout419 net421 vssd1 vssd1 vccd1 vccd1 net419 sky130_fd_sc_hd__clkbuf_8
XANTENNA__10105__S net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09750_ top.pc\[12\] _04352_ vssd1 vssd1 vccd1 vccd1 _04773_ sky130_fd_sc_hd__nand2_1
X_06962_ _02094_ _02096_ _02098_ _02100_ vssd1 vssd1 vccd1 vccd1 _02101_ sky130_fd_sc_hd__or4_1
XANTENNA__13639__RESET_B net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08701_ net290 _03209_ _03215_ vssd1 vssd1 vccd1 vccd1 _03820_ sky130_fd_sc_hd__and3_1
X_09681_ net795 _04715_ vssd1 vssd1 vccd1 vccd1 _04717_ sky130_fd_sc_hd__or2_1
X_06893_ top.DUT.register\[12\]\[18\] net740 net716 top.DUT.register\[27\]\[18\] vssd1
+ vssd1 vccd1 vccd1 _02032_ sky130_fd_sc_hd__a22o_1
X_08632_ _03331_ _03333_ net320 vssd1 vssd1 vccd1 vccd1 _03754_ sky130_fd_sc_hd__o21a_1
XFILLER_0_179_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07922__B _02522_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13292__RESET_B net1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07896__A2 net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08563_ _03601_ _03687_ net309 vssd1 vssd1 vccd1 vccd1 _03688_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_583 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07514_ net807 _02652_ net437 vssd1 vssd1 vccd1 vccd1 _02653_ sky130_fd_sc_hd__o21a_1
XFILLER_0_49_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08494_ _02880_ _03408_ _03538_ vssd1 vssd1 vccd1 vccd1 _03622_ sky130_fd_sc_hd__o21a_1
XANTENNA__07648__A2 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06856__B1 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07445_ top.DUT.register\[9\]\[15\] net467 net465 top.DUT.register\[13\]\[15\] _02583_
+ vssd1 vssd1 vccd1 vccd1 _02584_ sky130_fd_sc_hd__a221o_1
XFILLER_0_9_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10775__S net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout330_A net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09849__B _01584_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1072_A net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout428_A net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_236 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_379 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_118_2215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07376_ top.DUT.register\[30\]\[8\] net759 _02503_ _02514_ vssd1 vssd1 vccd1 vccd1
+ _02515_ sky130_fd_sc_hd__a211o_1
XFILLER_0_147_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09115_ _03000_ _03040_ vssd1 vssd1 vccd1 vccd1 _04190_ sky130_fd_sc_hd__nor2_1
XANTENNA__06608__B1 net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06327_ net896 _01389_ _01472_ vssd1 vssd1 vccd1 vccd1 _01474_ sky130_fd_sc_hd__nor3_2
XFILLER_0_32_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_40_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09046_ net284 _03498_ _03737_ _04041_ _03258_ vssd1 vssd1 vccd1 vccd1 _04121_ sky130_fd_sc_hd__a2111oi_1
XANTENNA__07281__B1 net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_2404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06258_ net2314 net853 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedData\[19\] sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_131_2415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07820__A2 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout797_A _05082_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold440 top.DUT.register\[14\]\[12\] vssd1 vssd1 vccd1 vccd1 net1556 sky130_fd_sc_hd__dlygate4sd3_1
X_06189_ _00009_ top.a1.nextHex\[7\] vssd1 vssd1 vccd1 vccd1 top.a1.nextHex\[2\] sky130_fd_sc_hd__or2_1
Xhold451 top.DUT.register\[8\]\[28\] vssd1 vssd1 vccd1 vccd1 net1567 sky130_fd_sc_hd__dlygate4sd3_1
Xhold462 top.DUT.register\[23\]\[13\] vssd1 vssd1 vccd1 vccd1 net1578 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07033__B1 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold473 top.DUT.register\[6\]\[17\] vssd1 vssd1 vccd1 vccd1 net1589 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07385__A _02497_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold484 top.DUT.register\[30\]\[15\] vssd1 vssd1 vccd1 vccd1 net1600 sky130_fd_sc_hd__dlygate4sd3_1
Xhold495 top.ramaddr\[16\] vssd1 vssd1 vccd1 vccd1 net1611 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout964_A net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout585_X net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout920 net921 vssd1 vssd1 vccd1 vccd1 net920 sky130_fd_sc_hd__clkbuf_2
XANTENNA__06387__A2 net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout931 net935 vssd1 vssd1 vccd1 vccd1 net931 sky130_fd_sc_hd__buf_2
Xfanout942 net943 vssd1 vssd1 vccd1 vccd1 net942 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10015__S net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09948_ net1594 net262 net629 vssd1 vssd1 vccd1 vccd1 _00156_ sky130_fd_sc_hd__mux2_1
Xfanout953 net956 vssd1 vssd1 vccd1 vccd1 net953 sky130_fd_sc_hd__clkbuf_4
Xfanout964 net965 vssd1 vssd1 vccd1 vccd1 net964 sky130_fd_sc_hd__clkbuf_4
Xfanout975 net977 vssd1 vssd1 vccd1 vccd1 net975 sky130_fd_sc_hd__clkbuf_4
Xfanout986 net987 vssd1 vssd1 vccd1 vccd1 net986 sky130_fd_sc_hd__buf_2
XFILLER_0_99_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_129_2377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout997 net1000 vssd1 vssd1 vccd1 vccd1 net997 sky130_fd_sc_hd__clkbuf_2
X_09879_ _04887_ _04888_ vssd1 vssd1 vccd1 vccd1 _04889_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout752_X net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_2388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1140 top.DUT.register\[21\]\[19\] vssd1 vssd1 vccd1 vccd1 net2256 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1151 top.pad.keyCode\[7\] vssd1 vssd1 vccd1 vccd1 net2267 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1162 top.pad.keyCode\[2\] vssd1 vssd1 vccd1 vccd1 net2278 sky130_fd_sc_hd__dlygate4sd3_1
X_11910_ _05759_ _05784_ vssd1 vssd1 vccd1 vccd1 _05793_ sky130_fd_sc_hd__or2_1
XFILLER_0_197_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1173 top.ramaddr\[14\] vssd1 vssd1 vccd1 vccd1 net2289 sky130_fd_sc_hd__dlygate4sd3_1
X_12890_ clknet_leaf_0_clk _00482_ net916 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[12\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07887__A2 net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_187_Left_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1184 top.DUT.register\[22\]\[7\] vssd1 vssd1 vccd1 vccd1 net2300 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1195 top.ramaddr\[14\] vssd1 vssd1 vccd1 vccd1 net2311 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10891__A1 net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11841_ net130 _05718_ _05703_ vssd1 vssd1 vccd1 vccd1 _05724_ sky130_fd_sc_hd__a21boi_1
XTAP_TAPCELL_ROW_142_2577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06448__B _01584_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08836__A1 net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11772_ _05644_ _05652_ _05637_ vssd1 vssd1 vccd1 vccd1 _05655_ sky130_fd_sc_hd__a21o_2
XFILLER_0_200_559 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06847__B1 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10723_ net2011 net160 net336 vssd1 vssd1 vccd1 vccd1 _00884_ sky130_fd_sc_hd__mux2_1
XFILLER_0_184_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13511_ clknet_leaf_9_clk _01103_ net945 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[31\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_586 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_175_3065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10685__S net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_175_3076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10654_ net171 net1920 net343 vssd1 vssd1 vccd1 vccd1 _00818_ sky130_fd_sc_hd__mux2_1
X_13442_ clknet_leaf_10_clk _01034_ net950 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[29\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_165_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13373_ clknet_leaf_127_clk _00965_ net920 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[27\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_10585_ net1818 net180 net353 vssd1 vssd1 vccd1 vccd1 _00751_ sky130_fd_sc_hd__mux2_1
Xclkload18 clknet_leaf_125_clk vssd1 vssd1 vccd1 vccd1 clkload18/Y sky130_fd_sc_hd__clkinv_2
Xclkload29 clknet_leaf_116_clk vssd1 vssd1 vccd1 vccd1 clkload29/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_106_563 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12324_ _06126_ net790 _06125_ vssd1 vssd1 vccd1 vccd1 _01360_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_58_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07272__B1 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12255_ _06084_ net979 _06083_ vssd1 vssd1 vccd1 vccd1 _01327_ sky130_fd_sc_hd__and3b_1
XANTENNA__06911__B _02007_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07024__B1 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11206_ _05109_ net1248 net471 vssd1 vssd1 vccd1 vccd1 _01253_ sky130_fd_sc_hd__mux2_1
X_12186_ top.a1.row2\[41\] net847 net797 _05719_ vssd1 vssd1 vccd1 vccd1 _01294_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_71_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11137_ net60 net868 vssd1 vssd1 vccd1 vccd1 _05074_ sky130_fd_sc_hd__and2_1
XFILLER_0_207_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11068_ net83 net870 net834 net1154 vssd1 vssd1 vccd1 vccd1 _01179_ sky130_fd_sc_hd__a22o_1
XFILLER_0_207_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08838__B _03950_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_500 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10019_ net1900 net253 net619 vssd1 vssd1 vccd1 vccd1 _00222_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07878__A2 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_69_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06550__A2 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_203_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08827__B2 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_715 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06838__B1 net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13709_ clknet_leaf_94_clk _01280_ net985 vssd1 vssd1 vccd1 vccd1 top.a1.row2\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_82_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_439 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07230_ top.DUT.register\[26\]\[10\] net750 net714 top.DUT.register\[27\]\[10\] vssd1
+ vssd1 vccd1 vccd1 _02369_ sky130_fd_sc_hd__a22o_1
XANTENNA__06374__A top.a1.instruction\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_647 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07161_ top.DUT.register\[16\]\[11\] net734 net635 top.DUT.register\[6\]\[11\] vssd1
+ vssd1 vccd1 vccd1 _02300_ sky130_fd_sc_hd__a22o_1
XANTENNA__08055__A2 _03122_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_171_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_656 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07263__B1 net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07092_ top.DUT.register\[28\]\[16\] net556 net515 top.DUT.register\[7\]\[16\] _02230_
+ vssd1 vssd1 vccd1 vccd1 _02231_ sky130_fd_sc_hd__a221o_1
XANTENNA__07802__A2 net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_2134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_2145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08669__A_N _02047_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout205 net206 vssd1 vssd1 vccd1 vccd1 net205 sky130_fd_sc_hd__buf_2
Xfanout216 net218 vssd1 vssd1 vccd1 vccd1 net216 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout227 net228 vssd1 vssd1 vccd1 vccd1 net227 sky130_fd_sc_hd__clkbuf_2
X_09802_ _04806_ _04807_ _04808_ vssd1 vssd1 vccd1 vccd1 _04820_ sky130_fd_sc_hd__o21ba_1
Xfanout238 _04757_ vssd1 vssd1 vccd1 vccd1 net238 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout249 _05439_ vssd1 vssd1 vccd1 vccd1 net249 sky130_fd_sc_hd__clkbuf_2
X_07994_ _03125_ _03127_ _03131_ _03132_ vssd1 vssd1 vccd1 vccd1 _03133_ sky130_fd_sc_hd__or4_1
X_06945_ top.DUT.register\[5\]\[21\] net654 net733 top.DUT.register\[14\]\[21\] _02083_
+ vssd1 vssd1 vccd1 vccd1 _02084_ sky130_fd_sc_hd__a221o_1
X_09733_ _03594_ net403 net488 _04759_ vssd1 vssd1 vccd1 vccd1 _04760_ sky130_fd_sc_hd__o211a_4
XFILLER_0_207_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout378_A net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06876_ top.DUT.register\[16\]\[18\] net544 net445 top.DUT.register\[1\]\[18\] _02014_
+ vssd1 vssd1 vccd1 vccd1 _02015_ sky130_fd_sc_hd__a221o_1
XANTENNA__07869__A2 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09664_ top.a1.halfData\[3\] _01471_ _04702_ net1086 vssd1 vssd1 vccd1 vccd1 _00118_
+ sky130_fd_sc_hd__o211a_1
X_08615_ net429 net427 _03737_ vssd1 vssd1 vccd1 vccd1 _03738_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_2_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09595_ net812 _04632_ _04641_ vssd1 vssd1 vccd1 vccd1 _04642_ sky130_fd_sc_hd__o21ai_1
XANTENNA__06541__A2 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06268__B net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout545_A net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08546_ net320 _03671_ _03670_ vssd1 vssd1 vccd1 vccd1 _03672_ sky130_fd_sc_hd__a21o_1
XANTENNA__08764__A net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06829__B1 net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08477_ net319 _03605_ vssd1 vssd1 vccd1 vccd1 _03606_ sky130_fd_sc_hd__or2_2
XANTENNA_fanout712_A net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09491__A1 _01887_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout333_X net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07428_ _02547_ _02566_ net825 vssd1 vssd1 vccd1 vccd1 _02567_ sky130_fd_sc_hd__mux2_2
XFILLER_0_147_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_21_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout500_X net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07359_ _02497_ vssd1 vssd1 vccd1 vccd1 _02498_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_21_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07254__B1 net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10370_ net1482 net235 net374 vssd1 vssd1 vccd1 vccd1 _00545_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_149_Right_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09029_ _04098_ _04099_ _04100_ _04103_ vssd1 vssd1 vccd1 vccd1 _04104_ sky130_fd_sc_hd__or4_1
XFILLER_0_130_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12040_ _05899_ _05910_ _05921_ vssd1 vssd1 vccd1 vccd1 _05923_ sky130_fd_sc_hd__a21bo_1
XANTENNA__09882__X _04892_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold270 top.DUT.register\[28\]\[17\] vssd1 vssd1 vccd1 vccd1 net1386 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08004__A _03122_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold281 top.DUT.register\[24\]\[31\] vssd1 vssd1 vccd1 vccd1 net1397 sky130_fd_sc_hd__dlygate4sd3_1
Xhold292 top.DUT.register\[18\]\[7\] vssd1 vssd1 vccd1 vccd1 net1408 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout967_X net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout750 _01621_ vssd1 vssd1 vccd1 vccd1 net750 sky130_fd_sc_hd__clkbuf_8
Xfanout761 _01617_ vssd1 vssd1 vccd1 vccd1 net761 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_144_2606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout772 _01614_ vssd1 vssd1 vccd1 vccd1 net772 sky130_fd_sc_hd__buf_6
XPHY_EDGE_ROW_195_Left_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout783 net784 vssd1 vssd1 vccd1 vccd1 net783 sky130_fd_sc_hd__buf_2
Xfanout794 _01581_ vssd1 vssd1 vccd1 vccd1 net794 sky130_fd_sc_hd__buf_2
XFILLER_0_99_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08506__B1 _03626_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08658__B net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12942_ clknet_leaf_41_clk _00534_ net1057 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[13\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_177_3105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12873_ clknet_leaf_50_clk _00465_ net1061 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[11\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06532__A2 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11824_ _05706_ vssd1 vssd1 vccd1 vccd1 _05707_ sky130_fd_sc_hd__inv_2
XFILLER_0_68_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11755_ _05623_ _05629_ vssd1 vssd1 vccd1 vccd1 _05638_ sky130_fd_sc_hd__and2_1
X_10706_ net1313 net228 net334 vssd1 vssd1 vccd1 vccd1 _00867_ sky130_fd_sc_hd__mux2_1
XFILLER_0_193_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11686_ _05568_ vssd1 vssd1 vccd1 vccd1 _05569_ sky130_fd_sc_hd__inv_2
XFILLER_0_125_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_155_2768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13425_ clknet_leaf_111_clk _01017_ net988 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[29\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_114_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10637_ net237 net1776 net343 vssd1 vssd1 vccd1 vccd1 _00801_ sky130_fd_sc_hd__mux2_1
Xclkload107 clknet_leaf_64_clk vssd1 vssd1 vccd1 vccd1 clkload107/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_141_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_319 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13356_ clknet_leaf_63_clk _00948_ net1091 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[26\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06481__X _01620_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11041__B2 top.ramload\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10568_ net1519 net252 net350 vssd1 vssd1 vccd1 vccd1 _00734_ sky130_fd_sc_hd__mux2_1
XANTENNA__09785__A2 net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_116_Right_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_178_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06599__A2 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12307_ _06114_ _06115_ net790 vssd1 vssd1 vccd1 vccd1 _01354_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_188_3267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13287_ clknet_leaf_8_clk _00879_ net947 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[24\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_10499_ net1841 net261 net358 vssd1 vssd1 vccd1 vccd1 _00668_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09792__X _04811_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12238_ top.lcd.cnt_20ms\[10\] top.lcd.cnt_20ms\[9\] _06070_ vssd1 vssd1 vccd1 vccd1
+ _06074_ sky130_fd_sc_hd__and3_1
X_12169_ net1299 net846 net796 _06042_ vssd1 vssd1 vccd1 vccd1 _01277_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_207_3551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08201__X _03339_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06771__A2 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput5 DAT_I[12] vssd1 vssd1 vccd1 vccd1 net5 sky130_fd_sc_hd__clkbuf_1
X_06730_ top.DUT.register\[12\]\[25\] net738 net702 top.DUT.register\[3\]\[25\] vssd1
+ vssd1 vccd1 vccd1 _01869_ sky130_fd_sc_hd__a22o_1
XFILLER_0_204_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06661_ top.DUT.register\[15\]\[26\] net682 net678 top.DUT.register\[31\]\[26\] vssd1
+ vssd1 vccd1 vccd1 _01800_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_84_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06523__A2 net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_503 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08400_ net275 _03524_ _03531_ _02830_ _03526_ vssd1 vssd1 vccd1 vccd1 _03532_ sky130_fd_sc_hd__a221o_1
X_09380_ _01930_ _01939_ _04438_ vssd1 vssd1 vccd1 vccd1 _04440_ sky130_fd_sc_hd__o21ai_1
X_06592_ top.DUT.register\[4\]\[28\] net670 net781 top.DUT.register\[25\]\[28\] _01729_
+ vssd1 vssd1 vccd1 vccd1 _01731_ sky130_fd_sc_hd__a221o_1
X_08331_ _03283_ _03297_ net312 vssd1 vssd1 vccd1 vccd1 _03465_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_98 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_191_528 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06287__A1 top.lcd.nextState\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08262_ _03397_ vssd1 vssd1 vccd1 vccd1 _03398_ sky130_fd_sc_hd__inv_2
XFILLER_0_46_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07213_ _02334_ _02351_ vssd1 vssd1 vccd1 vccd1 _02352_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_117_658 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08193_ _02995_ net276 _03288_ vssd1 vssd1 vccd1 vccd1 _03331_ sky130_fd_sc_hd__or3_1
XANTENNA_fanout126_A _05879_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07236__B1 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07144_ top.DUT.register\[17\]\[11\] net459 net455 top.DUT.register\[25\]\[11\] vssd1
+ vssd1 vccd1 vccd1 _02283_ sky130_fd_sc_hd__a22o_1
XFILLER_0_72_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07075_ top.DUT.register\[8\]\[22\] net640 net755 top.DUT.register\[1\]\[22\] _02211_
+ vssd1 vssd1 vccd1 vccd1 _02214_ sky130_fd_sc_hd__a221o_1
XFILLER_0_112_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout283_X net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout662_A _01606_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07977_ top.DUT.register\[2\]\[31\] net561 net528 top.DUT.register\[26\]\[31\] vssd1
+ vssd1 vccd1 vccd1 _03116_ sky130_fd_sc_hd__a22o_1
XFILLER_0_199_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06762__A2 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08478__B _03606_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09716_ net2195 net241 net631 vssd1 vssd1 vccd1 vccd1 _00127_ sky130_fd_sc_hd__mux2_1
X_06928_ top.DUT.register\[9\]\[21\] net469 net514 top.DUT.register\[24\]\[21\] _02066_
+ vssd1 vssd1 vccd1 vccd1 _02067_ sky130_fd_sc_hd__a221o_1
XFILLER_0_184_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09700__A2 net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout450_X net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09647_ top.pad.keyCode\[0\] top.pad.keyCode\[2\] top.pad.keyCode\[3\] top.pad.keyCode\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04689_ sky130_fd_sc_hd__or4b_1
X_06859_ top.DUT.register\[7\]\[19\] net661 net641 top.DUT.register\[8\]\[19\] _01997_
+ vssd1 vssd1 vccd1 vccd1 _01998_ sky130_fd_sc_hd__a221o_1
XANTENNA__08765__Y _03881_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout927_A net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout548_X net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06514__A2 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_195_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_322 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09578_ _04622_ _04623_ _04625_ _04619_ net134 vssd1 vssd1 vccd1 vccd1 _04626_ sky130_fd_sc_hd__o32a_1
XFILLER_0_167_547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08529_ net434 _03653_ _03655_ net427 vssd1 vssd1 vccd1 vccd1 _03656_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA_fanout715_X net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09464__A1 net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_194_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10529__A _04712_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_1999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_172_3024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11540_ top.a1.dataIn\[15\] _05328_ _05361_ vssd1 vssd1 vccd1 vccd1 _05423_ sky130_fd_sc_hd__or3_1
XFILLER_0_203_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11271__B2 top.a1.row1\[58\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xwire414 _02002_ vssd1 vssd1 vccd1 vccd1 net414 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_108_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11471_ _05351_ _05353_ vssd1 vssd1 vccd1 vccd1 _05354_ sky130_fd_sc_hd__nor2_1
XFILLER_0_92_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07227__B1 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13210_ clknet_leaf_1_clk _00802_ net916 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[22\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_10422_ net1543 net168 _04982_ vssd1 vssd1 vccd1 vccd1 _00594_ sky130_fd_sc_hd__mux2_1
XFILLER_0_116_680 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_2498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10353_ net1390 net174 net378 vssd1 vssd1 vccd1 vccd1 _00529_ sky130_fd_sc_hd__mux2_1
X_13141_ clknet_leaf_30_clk _00733_ net1020 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[20\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_150_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06461__B top.a1.instruction\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13072_ clknet_leaf_27_clk _00664_ net1010 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[17\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_150_2698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10284_ top.DUT.register\[11\]\[21\] net195 net387 vssd1 vssd1 vccd1 vccd1 _00462_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12023_ _05884_ _05905_ vssd1 vssd1 vccd1 vccd1 _05906_ sky130_fd_sc_hd__xnor2_2
XTAP_TAPCELL_ROW_183_3186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_183_3197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07950__A1 _01887_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06753__A2 net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout580 _01514_ vssd1 vssd1 vccd1 vccd1 net580 sky130_fd_sc_hd__buf_2
Xfanout591 _04971_ vssd1 vssd1 vccd1 vccd1 net591 sky130_fd_sc_hd__clkbuf_8
XANTENNA__10203__S net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07860__X _02999_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_650 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12925_ clknet_leaf_3_clk _00517_ net919 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[13\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06505__A2 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_202_3470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_202_3481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12856_ clknet_leaf_128_clk _00448_ net911 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[11\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_157_2808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11807_ _05646_ _05678_ _05681_ _05685_ _05689_ vssd1 vssd1 vccd1 vccd1 _05690_ sky130_fd_sc_hd__a41o_2
XFILLER_0_201_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12787_ clknet_leaf_124_clk _00379_ net926 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[9\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_113_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07466__B1 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11738_ _05620_ vssd1 vssd1 vccd1 vccd1 _05621_ sky130_fd_sc_hd__inv_2
XANTENNA__11261__C _05148_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10873__S net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_181_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11669_ _05546_ _05551_ vssd1 vssd1 vccd1 vccd1 _05552_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_98_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_291 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_431 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13408_ clknet_leaf_79_clk _01000_ net1072 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[28\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_113_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08966__B1 _02218_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_486 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13339_ clknet_leaf_124_clk _00931_ net925 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[26\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13065__RESET_B net1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11317__A2 _05148_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_168_2959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07900_ _03032_ _03034_ _03036_ _03038_ vssd1 vssd1 vccd1 vccd1 _03039_ sky130_fd_sc_hd__or4_4
X_08880_ net884 top.pc\[28\] net695 _03990_ vssd1 vssd1 vccd1 vccd1 _03991_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_4_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_208_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07831_ top.DUT.register\[7\]\[0\] net659 net639 top.DUT.register\[8\]\[0\] _02969_
+ vssd1 vssd1 vccd1 vccd1 _02970_ sky130_fd_sc_hd__a221o_1
XANTENNA__06744__A2 net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10113__S net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07762_ top.a1.instruction\[22\] _01507_ net793 net893 _02900_ vssd1 vssd1 vccd1
+ vccd1 _02901_ sky130_fd_sc_hd__a221o_1
XFILLER_0_79_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_108_2066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09143__B1 _04216_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09501_ _04551_ _04552_ vssd1 vssd1 vccd1 vccd1 _04553_ sky130_fd_sc_hd__and2_1
X_06713_ _01847_ _01849_ _01851_ vssd1 vssd1 vccd1 vccd1 _01852_ sky130_fd_sc_hd__or3_1
X_07693_ top.DUT.register\[28\]\[4\] net557 net544 top.DUT.register\[16\]\[4\] _02831_
+ vssd1 vssd1 vccd1 vccd1 _02832_ sky130_fd_sc_hd__a221o_1
XFILLER_0_189_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09694__A1 top.pc\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06644_ _01773_ _01782_ vssd1 vssd1 vccd1 vccd1 _01783_ sky130_fd_sc_hd__nor2_1
X_09432_ _04469_ _04473_ vssd1 vssd1 vccd1 vccd1 _04489_ sky130_fd_sc_hd__nand2_1
XANTENNA__06386__X _01525_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_154_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_2255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_121_2266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06575_ top.DUT.register\[2\]\[28\] net562 net505 top.DUT.register\[27\]\[28\] vssd1
+ vssd1 vccd1 vccd1 _01714_ sky130_fd_sc_hd__a22o_1
X_09363_ _04401_ _04404_ _04405_ vssd1 vssd1 vccd1 vccd1 _04424_ sky130_fd_sc_hd__o21ai_2
XANTENNA__13721__Q top.a1.row2\[35\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout243_A _04745_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08314_ _03225_ _03233_ vssd1 vssd1 vccd1 vccd1 _03449_ sky130_fd_sc_hd__and2_1
XFILLER_0_19_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07457__B1 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09294_ net136 _04345_ _04358_ net897 vssd1 vssd1 vccd1 vccd1 _04359_ sky130_fd_sc_hd__o211ai_1
XANTENNA_10 _05147_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08245_ _02946_ _03185_ vssd1 vssd1 vccd1 vccd1 _03382_ sky130_fd_sc_hd__nor2_1
XFILLER_0_28_792 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10783__S net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout410_A net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09857__B _04543_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_291 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout508_A _01565_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07658__A _02796_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08176_ _03306_ _03313_ net312 vssd1 vssd1 vccd1 vccd1 _03314_ sky130_fd_sc_hd__mux2_1
X_07127_ _02263_ _02265_ vssd1 vssd1 vccd1 vccd1 _02266_ sky130_fd_sc_hd__or2_2
XANTENNA_clkbuf_leaf_63_clk_A clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1038_X net1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07058_ _02190_ _02192_ _02194_ _02196_ vssd1 vssd1 vccd1 vccd1 _02197_ sky130_fd_sc_hd__or4_2
XANTENNA__11308__A2 _05136_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout498_X net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_78_clk_A clknet_4_12__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout665_X net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07932__A1 _02623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12788__RESET_B net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_121_clk_A clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10023__S net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10971_ top.a1.dataInTemp\[2\] net785 vssd1 vssd1 vccd1 vccd1 _05012_ sky130_fd_sc_hd__or2_1
XFILLER_0_97_434 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout832_X net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08495__Y _03623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_136 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12710_ clknet_leaf_38_clk _00302_ net1053 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[6\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11643__A top.a1.dataIn\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07696__B1 net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13690_ clknet_leaf_71_clk _00002_ vssd1 vssd1 vccd1 vccd1 top.lcd.nextState\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__06737__A _01853_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07160__A2 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12641_ clknet_leaf_15_clk _00233_ net961 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[4\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_155_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_139_2527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_139_2538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_16_clk_A clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07448__B1 net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12572_ clknet_leaf_130_clk _00164_ net909 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[2\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11523_ _05403_ _05405_ _05400_ vssd1 vssd1 vccd1 vccd1 _05406_ sky130_fd_sc_hd__a21o_1
XANTENNA__10693__S net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08660__A2 net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_152_2727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11454_ _05303_ _05304_ _05324_ _05287_ _05299_ vssd1 vssd1 vccd1 vccd1 _05337_ sky130_fd_sc_hd__a221o_1
XFILLER_0_123_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10405_ net1441 net237 net369 vssd1 vssd1 vccd1 vccd1 _00577_ sky130_fd_sc_hd__mux2_1
X_11385_ _05249_ _05250_ _05236_ vssd1 vssd1 vccd1 vccd1 _05268_ sky130_fd_sc_hd__a21oi_2
XANTENNA__09070__C1 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_672 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_185_3215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07855__X _02994_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13124_ clknet_leaf_36_clk _00716_ net1049 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[19\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_185_3226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10336_ net2023 net245 net377 vssd1 vssd1 vccd1 vccd1 _00512_ sky130_fd_sc_hd__mux2_1
XANTENNA__07620__B1 net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06974__A2 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11818__A top.a1.dataIn\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10267_ net1385 net258 net387 vssd1 vssd1 vccd1 vccd1 _00445_ sky130_fd_sc_hd__mux2_1
X_13055_ clknet_leaf_24_clk _00647_ net1013 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[17\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08970__A2_N net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08399__A _03530_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_175_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12006_ _05865_ _05866_ net126 vssd1 vssd1 vccd1 vccd1 _05889_ sky130_fd_sc_hd__and3_1
X_10198_ net267 net1984 net394 vssd1 vssd1 vccd1 vccd1 _00378_ sky130_fd_sc_hd__mux2_1
XANTENNA__11180__B1 net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_204_3510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06726__A2 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_205_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11256__C _05148_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_205_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_163_2889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10868__S net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09676__A1 top.a1.instruction\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08479__A2 net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12908_ clknet_leaf_47_clk _00500_ net1069 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[12\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08884__C1 net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06647__A _01764_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_186_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_158_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07151__A2 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_196_3388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13541__Q top.ramload\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12839_ clknet_leaf_6_clk _00431_ net937 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[10\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_174_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06366__B net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_17_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06360_ top.ru.state\[2\] net887 _00011_ net873 vssd1 vssd1 vccd1 vccd1 _01499_ sky130_fd_sc_hd__a211o_1
XANTENNA__07439__B1 net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06291_ _01331_ vssd1 vssd1 vccd1 vccd1 _01450_ sky130_fd_sc_hd__inv_2
XFILLER_0_142_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08030_ _03160_ _03167_ vssd1 vssd1 vccd1 vccd1 _03169_ sky130_fd_sc_hd__or2_2
XFILLER_0_141_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput30 DAT_I[6] vssd1 vssd1 vccd1 vccd1 net30 sky130_fd_sc_hd__buf_1
XANTENNA__09396__C _04453_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold803 top.DUT.register\[10\]\[21\] vssd1 vssd1 vccd1 vccd1 net1919 sky130_fd_sc_hd__dlygate4sd3_1
Xhold814 top.DUT.register\[10\]\[20\] vssd1 vssd1 vccd1 vccd1 net1930 sky130_fd_sc_hd__dlygate4sd3_1
Xhold825 top.DUT.register\[13\]\[10\] vssd1 vssd1 vccd1 vccd1 net1941 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10108__S net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold836 top.DUT.register\[16\]\[14\] vssd1 vssd1 vccd1 vccd1 net1952 sky130_fd_sc_hd__dlygate4sd3_1
Xhold847 top.DUT.register\[14\]\[4\] vssd1 vssd1 vccd1 vccd1 net1963 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07765__X _02904_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_1829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold858 top.DUT.register\[19\]\[20\] vssd1 vssd1 vccd1 vccd1 net1974 sky130_fd_sc_hd__dlygate4sd3_1
Xhold869 top.DUT.register\[31\]\[9\] vssd1 vssd1 vccd1 vccd1 net1985 sky130_fd_sc_hd__dlygate4sd3_1
X_09981_ net269 net2013 net624 vssd1 vssd1 vccd1 vccd1 _00186_ sky130_fd_sc_hd__mux2_1
XANTENNA__06965__A2 net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08932_ _03143_ net492 _04039_ vssd1 vssd1 vccd1 vccd1 _04040_ sky130_fd_sc_hd__o21ai_1
XANTENNA__10191__X _04971_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08863_ _01786_ _03973_ vssd1 vssd1 vccd1 vccd1 _03974_ sky130_fd_sc_hd__nor2_1
XANTENNA__08102__A _02590_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout193_A _04850_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06717__A2 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07814_ _02952_ vssd1 vssd1 vccd1 vccd1 _02953_ sky130_fd_sc_hd__inv_2
XANTENNA__08596__X _03720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08794_ _03897_ _03906_ _03908_ vssd1 vssd1 vccd1 vccd1 _03909_ sky130_fd_sc_hd__or3_2
XANTENNA__07941__A _02242_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07390__A2 net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07745_ top.DUT.register\[4\]\[3\] net510 net441 top.DUT.register\[5\]\[3\] _02883_
+ vssd1 vssd1 vccd1 vccd1 _02884_ sky130_fd_sc_hd__a221o_1
XANTENNA__10778__S net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout458_A _01553_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_9_Left_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09131__A3 net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07676_ top.DUT.register\[24\]\[4\] net646 net763 top.DUT.register\[9\]\[4\] _02810_
+ vssd1 vssd1 vccd1 vccd1 _02815_ sky130_fd_sc_hd__a221o_1
XANTENNA__07142__A2 net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09415_ _01983_ _04471_ vssd1 vssd1 vccd1 vccd1 _04473_ sky130_fd_sc_hd__or2_1
X_06627_ top.DUT.register\[24\]\[27\] net646 net725 top.DUT.register\[29\]\[27\] vssd1
+ vssd1 vccd1 vccd1 _01766_ sky130_fd_sc_hd__a22o_1
XANTENNA__09419__A1 net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_181_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_36_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout625_A net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06558_ _01683_ _01688_ _01696_ vssd1 vssd1 vccd1 vccd1 _01697_ sky130_fd_sc_hd__nor3_2
XFILLER_0_191_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09346_ net132 _04400_ _04407_ net810 vssd1 vssd1 vccd1 vccd1 _04408_ sky130_fd_sc_hd__o22a_1
XANTENNA__06844__X _01983_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_1958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10012__A_N top.a1.instruction\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_192_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06489_ net788 _01611_ _01618_ vssd1 vssd1 vccd1 vccd1 _01628_ sky130_fd_sc_hd__and3_4
X_09277_ net132 _04333_ _04341_ _04342_ net897 vssd1 vssd1 vccd1 vccd1 _04343_ sky130_fd_sc_hd__o221a_1
XFILLER_0_90_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_43_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_43_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08228_ _03211_ _03216_ net292 vssd1 vssd1 vccd1 vccd1 _03365_ sky130_fd_sc_hd__mux2_1
XANTENNA__07850__B1 net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout994_A net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_134_2457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08159_ _03296_ vssd1 vssd1 vccd1 vccd1 _03297_ sky130_fd_sc_hd__inv_2
XANTENNA__10018__S net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07602__B1 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11170_ top.a1.row1\[60\] _05094_ _05085_ vssd1 vssd1 vccd1 vccd1 _01232_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_787 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10121_ net235 net1538 net608 vssd1 vssd1 vccd1 vccd1 _00321_ sky130_fd_sc_hd__mux2_1
XANTENNA__06956__A2 net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10052_ net1668 net251 net615 vssd1 vssd1 vccd1 vccd1 _00254_ sky130_fd_sc_hd__mux2_1
XANTENNA__06708__A2 net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_180_3145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13811_ net72 vssd1 vssd1 vccd1 vccd1 net108 sky130_fd_sc_hd__clkbuf_1
XANTENNA__10688__S net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input19_A DAT_I[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13742_ clknet_leaf_100_clk _01313_ vssd1 vssd1 vccd1 vccd1 top.lcd.cnt_20ms\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_10954_ net904 _01409_ _01416_ _04996_ vssd1 vssd1 vccd1 vccd1 _04997_ sky130_fd_sc_hd__or4b_1
XFILLER_0_58_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07133__A2 net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13673_ clknet_leaf_90_clk _01249_ net999 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_10885_ net154 top.DUT.register\[29\]\[29\] net597 vssd1 vssd1 vccd1 vccd1 _01046_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_168_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12624_ clknet_leaf_28_clk _00216_ net1010 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[3\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08618__C1 _03740_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12555_ clknet_leaf_46_clk _00147_ net1065 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[1\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_183_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_170_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_170_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_274 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11506_ _05346_ _05348_ _05357_ vssd1 vssd1 vccd1 vccd1 _05389_ sky130_fd_sc_hd__and3_1
XANTENNA__07841__B1 net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12486_ clknet_leaf_46_clk _00081_ net1090 vssd1 vssd1 vccd1 vccd1 top.ramstore\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_34_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12354__D net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11437_ _05277_ _05284_ _05281_ vssd1 vssd1 vccd1 vccd1 _05320_ sky130_fd_sc_hd__a21o_1
XFILLER_0_80_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11368_ _05249_ _05250_ vssd1 vssd1 vccd1 vccd1 _05251_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_210_3591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06947__A2 net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13107_ clknet_leaf_123_clk _00699_ net926 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[19\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10319_ net176 net1924 net382 vssd1 vssd1 vccd1 vccd1 _00496_ sky130_fd_sc_hd__mux2_1
X_11299_ net1191 net813 _05187_ net1078 vssd1 vssd1 vccd1 vccd1 _01268_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_165_2918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13038_ clknet_leaf_41_clk _00630_ net1057 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[16\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_178_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07372__A2 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_198_3417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13131__CLK clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07761__A top.a1.instruction\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_406 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10598__S net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_2014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06580__B1 net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_2025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_89_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07530_ top.DUT.register\[15\]\[7\] net679 net675 top.DUT.register\[31\]\[7\] vssd1
+ vssd1 vccd1 vccd1 _02669_ sky130_fd_sc_hd__a22o_1
XFILLER_0_49_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07461_ top.DUT.register\[8\]\[15\] net640 net719 top.DUT.register\[19\]\[15\] _02592_
+ vssd1 vssd1 vccd1 vccd1 _02600_ sky130_fd_sc_hd__a221o_1
XFILLER_0_48_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_201_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06412_ top.DUT.register\[26\]\[30\] net528 _01549_ vssd1 vssd1 vccd1 vccd1 _01551_
+ sky130_fd_sc_hd__a21o_1
X_09200_ _04268_ _04269_ vssd1 vssd1 vccd1 vccd1 _04270_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_33_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07392_ top.DUT.register\[9\]\[9\] net467 net524 top.DUT.register\[11\]\[9\] _02530_
+ vssd1 vssd1 vccd1 vccd1 _02531_ sky130_fd_sc_hd__a221o_1
XFILLER_0_57_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06343_ top.a1.instruction\[13\] net893 vssd1 vssd1 vccd1 vccd1 _01485_ sky130_fd_sc_hd__and2_2
X_09131_ top.pc\[2\] net827 net411 _04203_ _04205_ vssd1 vssd1 vccd1 vccd1 _04206_
+ sky130_fd_sc_hd__a311o_1
XFILLER_0_174_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10186__X _04966_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08624__A2 net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_98 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09062_ _03561_ _03589_ _03623_ _03655_ vssd1 vssd1 vccd1 vccd1 _04137_ sky130_fd_sc_hd__or4_1
X_06274_ _01436_ vssd1 vssd1 vccd1 vccd1 _01437_ sky130_fd_sc_hd__inv_2
X_08013_ _02351_ _03150_ _01500_ vssd1 vssd1 vccd1 vccd1 _03152_ sky130_fd_sc_hd__o21a_2
XFILLER_0_8_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold600 top.DUT.register\[31\]\[21\] vssd1 vssd1 vccd1 vccd1 net1716 sky130_fd_sc_hd__dlygate4sd3_1
Xhold611 top.DUT.register\[2\]\[20\] vssd1 vssd1 vccd1 vccd1 net1727 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_116_2187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold622 top.DUT.register\[13\]\[8\] vssd1 vssd1 vccd1 vccd1 net1738 sky130_fd_sc_hd__dlygate4sd3_1
Xhold633 top.DUT.register\[23\]\[26\] vssd1 vssd1 vccd1 vccd1 net1749 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07936__A _01983_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold644 top.ramaddr\[29\] vssd1 vssd1 vccd1 vccd1 net1760 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_83 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold655 top.DUT.register\[6\]\[13\] vssd1 vssd1 vccd1 vccd1 net1771 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06399__B1 net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06938__A2 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold666 top.DUT.register\[18\]\[23\] vssd1 vssd1 vccd1 vccd1 net1782 sky130_fd_sc_hd__dlygate4sd3_1
Xhold677 top.ramload\[0\] vssd1 vssd1 vccd1 vccd1 net1793 sky130_fd_sc_hd__dlygate4sd3_1
Xhold688 top.DUT.register\[25\]\[1\] vssd1 vssd1 vccd1 vccd1 net1804 sky130_fd_sc_hd__dlygate4sd3_1
X_09964_ net2121 net185 net629 vssd1 vssd1 vccd1 vccd1 _00172_ sky130_fd_sc_hd__mux2_1
Xhold699 top.DUT.register\[18\]\[10\] vssd1 vssd1 vccd1 vccd1 net1815 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08915_ net284 net429 _03498_ _04023_ vssd1 vssd1 vccd1 vccd1 _04024_ sky130_fd_sc_hd__a31o_1
X_09895_ top.a1.instruction\[27\] net486 net402 top.a1.dataIn\[27\] net398 vssd1 vssd1
+ vccd1 vccd1 _04904_ sky130_fd_sc_hd__a221o_2
XANTENNA_fanout575_A net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08846_ _03876_ _03957_ net313 vssd1 vssd1 vccd1 vccd1 _03958_ sky130_fd_sc_hd__mux2_1
XANTENNA__09870__B _04560_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07899__B1 net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08767__A net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08777_ _02136_ _02222_ _03851_ vssd1 vssd1 vccd1 vccd1 _03892_ sky130_fd_sc_hd__nor3b_1
XANTENNA_fanout742_A _01623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06558__Y _01697_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06571__B1 net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout363_X net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10301__S net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07728_ top.DUT.register\[4\]\[3\] net669 net665 top.DUT.register\[20\]\[3\] _02866_
+ vssd1 vssd1 vccd1 vccd1 _02867_ sky130_fd_sc_hd__a221o_1
XANTENNA__09731__A1_N net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07115__A2 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_177_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout530_X net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07659_ _02777_ _02797_ net825 vssd1 vssd1 vccd1 vccd1 _02798_ sky130_fd_sc_hd__mux2_2
XTAP_TAPCELL_ROW_45_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout628_X net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10670_ net2008 net235 net339 vssd1 vssd1 vccd1 vccd1 _00833_ sky130_fd_sc_hd__mux2_1
XFILLER_0_192_442 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07610__S net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09329_ _04389_ _04391_ vssd1 vssd1 vccd1 vccd1 _04392_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_192_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08615__A2 net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09812__A1 _02679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09885__X _04895_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12340_ top.pad.button_control.r_counter\[14\] _06134_ top.pad.button_control.r_counter\[15\]
+ vssd1 vssd1 vccd1 vccd1 _06136_ sky130_fd_sc_hd__a21o_1
XFILLER_0_180_659 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09110__B _03000_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_211_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07823__B1 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12525__Q top.a1.halfData\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12271_ top.lcd.cnt_500hz\[5\] top.lcd.cnt_500hz\[4\] _01436_ top.lcd.cnt_500hz\[6\]
+ vssd1 vssd1 vccd1 vccd1 _06093_ sky130_fd_sc_hd__a31o_1
XANTENNA__08379__A1 net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08379__B2 _03334_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11222_ top.a1.state\[1\] _05084_ net472 net1146 vssd1 vssd1 vccd1 vccd1 _01262_
+ sky130_fd_sc_hd__a22o_1
X_11153_ _04658_ net850 vssd1 vssd1 vccd1 vccd1 _05083_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_56_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10104_ net1773 net175 net614 vssd1 vssd1 vccd1 vccd1 _00305_ sky130_fd_sc_hd__mux2_1
XANTENNA__11087__B net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11084_ net906 net2018 net861 _05047_ vssd1 vssd1 vccd1 vccd1 _01193_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_147_2648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10035_ net1412 net194 net621 vssd1 vssd1 vccd1 vccd1 _00238_ sky130_fd_sc_hd__mux2_1
XANTENNA__08000__B1 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07354__A2 net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_203_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_19_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_160_2848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10211__S net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_187_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11986_ _05828_ _05868_ vssd1 vssd1 vccd1 vccd1 _05869_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07106__A2 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13725_ clknet_leaf_95_clk _01296_ net986 vssd1 vssd1 vccd1 vccd1 top.a1.row2\[43\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10937_ net1534 net215 net593 vssd1 vssd1 vccd1 vccd1 _01098_ sky130_fd_sc_hd__mux2_1
XFILLER_0_196_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_193_3336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_193_3347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06484__X _01623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13656_ clknet_leaf_94_clk _00014_ net994 vssd1 vssd1 vccd1 vccd1 wb.curr_state\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_85_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_183_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10868_ net213 net1805 net594 vssd1 vssd1 vccd1 vccd1 _01029_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12607_ clknet_leaf_24_clk _00199_ net1015 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[3\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_155_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13587_ clknet_leaf_46_clk net1144 net1066 vssd1 vssd1 vccd1 vccd1 net78 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10799_ net245 top.DUT.register\[27\]\[7\] net598 vssd1 vssd1 vccd1 vccd1 _00960_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__09795__X _04814_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12538_ clknet_leaf_2_clk _00130_ net916 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[1\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_124_542 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_79 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10881__S net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07290__A1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12469_ clknet_leaf_47_clk _00064_ net1066 vssd1 vssd1 vccd1 vccd1 top.ramstore\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_151_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06931__Y _02070_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08204__X _03342_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11278__A _05121_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07593__A2 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06961_ top.DUT.register\[2\]\[23\] net561 net460 top.DUT.register\[17\]\[23\] _02099_
+ vssd1 vssd1 vccd1 vccd1 _02100_ sky130_fd_sc_hd__a221o_1
XANTENNA__12402__RESET_B net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_207_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08700_ net296 _03453_ net325 vssd1 vssd1 vccd1 vccd1 _03819_ sky130_fd_sc_hd__a21o_1
X_09680_ net795 _04715_ vssd1 vssd1 vccd1 vccd1 _04716_ sky130_fd_sc_hd__nor2_2
X_06892_ top.DUT.register\[23\]\[18\] net673 net658 top.DUT.register\[21\]\[18\] _02030_
+ vssd1 vssd1 vccd1 vccd1 _02031_ sky130_fd_sc_hd__a221o_1
XANTENNA__07345__A2 net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08631_ net428 _03750_ _03751_ _03752_ vssd1 vssd1 vccd1 vccd1 _03753_ sky130_fd_sc_hd__a211o_1
XANTENNA__06553__B1 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08562_ _03648_ _03686_ net290 vssd1 vssd1 vccd1 vccd1 _03687_ sky130_fd_sc_hd__mux2_1
XANTENNA__10121__S net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07513_ _02644_ _02651_ vssd1 vssd1 vccd1 vccd1 _02652_ sky130_fd_sc_hd__nor2_4
XFILLER_0_193_206 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08493_ net286 _03395_ _03405_ net275 vssd1 vssd1 vccd1 vccd1 _03621_ sky130_fd_sc_hd__a22o_1
XFILLER_0_159_472 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout156_A _04916_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11741__A top.a1.dataIn\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07444_ top.DUT.register\[22\]\[15\] net578 net560 top.DUT.register\[2\]\[15\] vssd1
+ vssd1 vccd1 vccd1 _02583_ sky130_fd_sc_hd__a22o_1
XFILLER_0_18_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_204 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_99_Left_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10628__Y _04992_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_174_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09211__A _01505_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07375_ top.DUT.register\[5\]\[8\] net652 net765 top.DUT.register\[9\]\[8\] _02511_
+ vssd1 vssd1 vccd1 vccd1 _02514_ sky130_fd_sc_hd__a221o_1
XFILLER_0_91_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_118_2216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout323_A net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09114_ net827 net411 _04188_ net806 vssd1 vssd1 vccd1 vccd1 _04189_ sky130_fd_sc_hd__a22o_1
XFILLER_0_161_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06326_ top.a1.instruction\[6\] _01472_ vssd1 vssd1 vccd1 vccd1 _01473_ sky130_fd_sc_hd__nor2_2
XFILLER_0_17_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_161_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09045_ _03204_ _03328_ _03370_ net281 vssd1 vssd1 vccd1 vccd1 _04120_ sky130_fd_sc_hd__a31o_1
X_06257_ net1706 net852 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedData\[18\] sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_131_2405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10791__S net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_2416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold430 top.DUT.register\[2\]\[8\] vssd1 vssd1 vccd1 vccd1 net1546 sky130_fd_sc_hd__dlygate4sd3_1
X_06188_ _01425_ net1650 _01419_ vssd1 vssd1 vccd1 vccd1 top.a1.nextHex\[1\] sky130_fd_sc_hd__mux2_1
Xhold441 top.DUT.register\[10\]\[14\] vssd1 vssd1 vccd1 vccd1 net1557 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout692_A _04050_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold452 top.DUT.register\[12\]\[4\] vssd1 vssd1 vccd1 vccd1 net1568 sky130_fd_sc_hd__dlygate4sd3_1
Xhold463 top.DUT.register\[25\]\[28\] vssd1 vssd1 vccd1 vccd1 net1579 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_187_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold474 top.DUT.register\[28\]\[19\] vssd1 vssd1 vccd1 vccd1 net1590 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07385__B _02522_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1020_X net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold485 top.DUT.register\[26\]\[1\] vssd1 vssd1 vccd1 vccd1 net1601 sky130_fd_sc_hd__dlygate4sd3_1
Xhold496 top.DUT.register\[8\]\[10\] vssd1 vssd1 vccd1 vccd1 net1612 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout910 net935 vssd1 vssd1 vccd1 vccd1 net910 sky130_fd_sc_hd__clkbuf_4
Xfanout921 net922 vssd1 vssd1 vccd1 vccd1 net921 sky130_fd_sc_hd__clkbuf_2
Xfanout932 net934 vssd1 vssd1 vccd1 vccd1 net932 sky130_fd_sc_hd__clkbuf_4
X_09947_ net2061 net265 net627 vssd1 vssd1 vccd1 vccd1 _00155_ sky130_fd_sc_hd__mux2_1
Xfanout943 net967 vssd1 vssd1 vccd1 vccd1 net943 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout480_X net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout954 net956 vssd1 vssd1 vccd1 vccd1 net954 sky130_fd_sc_hd__clkbuf_2
XANTENNA__06792__B1 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout578_X net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout965 net966 vssd1 vssd1 vccd1 vccd1 net965 sky130_fd_sc_hd__buf_2
Xfanout976 net977 vssd1 vssd1 vccd1 vccd1 net976 sky130_fd_sc_hd__clkbuf_4
Xfanout987 net1007 vssd1 vssd1 vccd1 vccd1 net987 sky130_fd_sc_hd__buf_2
X_09878_ top.pc\[26\] _04577_ vssd1 vssd1 vccd1 vccd1 _04888_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_129_2378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08497__A net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout998 net1000 vssd1 vssd1 vccd1 vccd1 net998 sky130_fd_sc_hd__clkbuf_4
Xhold1130 top.DUT.register\[4\]\[31\] vssd1 vssd1 vccd1 vccd1 net2246 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1141 top.ramload\[7\] vssd1 vssd1 vccd1 vccd1 net2257 sky130_fd_sc_hd__dlygate4sd3_1
X_08829_ _01832_ net433 net501 _01831_ _03883_ vssd1 vssd1 vccd1 vccd1 _03942_ sky130_fd_sc_hd__a221o_1
Xhold1152 top.pad.count\[1\] vssd1 vssd1 vccd1 vccd1 net2268 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1163 top.DUT.register\[28\]\[18\] vssd1 vssd1 vccd1 vccd1 net2279 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06544__B1 net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout745_X net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1174 top.DUT.register\[1\]\[31\] vssd1 vssd1 vccd1 vccd1 net2290 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1185 top.DUT.register\[5\]\[29\] vssd1 vssd1 vccd1 vccd1 net2301 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_197_523 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1196 top.ramload\[13\] vssd1 vssd1 vccd1 vccd1 net2312 sky130_fd_sc_hd__dlygate4sd3_1
X_11840_ _05695_ _05720_ vssd1 vssd1 vccd1 vccd1 _05723_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10031__S net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_142_2578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11771_ _05644_ _05652_ vssd1 vssd1 vccd1 vccd1 _05654_ sky130_fd_sc_hd__nand2_1
XFILLER_0_184_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13510_ clknet_leaf_38_clk _01102_ net1054 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[31\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_10722_ net1741 net167 net336 vssd1 vssd1 vccd1 vccd1 _00883_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_175_3066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_175_3077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08049__B1 net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13441_ clknet_leaf_16_clk _01033_ net962 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[29\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_10653_ net173 net1671 net344 vssd1 vssd1 vccd1 vccd1 _00817_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13372_ clknet_leaf_0_clk _00964_ net909 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[27\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_63_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10584_ net1523 net192 net352 vssd1 vssd1 vccd1 vccd1 _00750_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkload19 clknet_leaf_126_clk vssd1 vssd1 vccd1 vccd1 clkload19/Y sky130_fd_sc_hd__clkinv_8
X_12323_ top.pad.button_control.r_counter\[8\] top.pad.button_control.r_counter\[7\]
+ _06122_ vssd1 vssd1 vccd1 vccd1 _06126_ sky130_fd_sc_hd__and3_1
XFILLER_0_2_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_575 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_692 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12913__RESET_B net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12254_ top.lcd.cnt_20ms\[16\] top.lcd.cnt_20ms\[15\] _06080_ vssd1 vssd1 vccd1 vccd1
+ _06084_ sky130_fd_sc_hd__and3_1
XANTENNA__06911__C _02049_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11205_ net845 _05019_ _05030_ vssd1 vssd1 vccd1 vccd1 _05109_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_71_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12185_ top.a1.row2\[40\] net847 net797 _05752_ vssd1 vssd1 vccd1 vccd1 _01293_ sky130_fd_sc_hd__a22o_1
XANTENNA__10206__S net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07575__A2 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11136_ net907 net1317 net862 _05073_ vssd1 vssd1 vccd1 vccd1 _01219_ sky130_fd_sc_hd__a31o_1
XANTENNA__06783__B1 net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_207_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11067_ net82 net871 net835 net1134 vssd1 vssd1 vccd1 vccd1 _01178_ sky130_fd_sc_hd__a22o_1
XANTENNA__07327__A2 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10018_ net2239 net255 net621 vssd1 vssd1 vccd1 vccd1 _00221_ sky130_fd_sc_hd__mux2_1
XFILLER_0_188_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06535__B1 net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_203_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_370 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09730__S net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_206 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10876__S net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11969_ _05755_ _05851_ vssd1 vssd1 vccd1 vccd1 _05852_ sky130_fd_sc_hd__xnor2_1
XANTENNA__13019__RESET_B net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13708_ clknet_leaf_95_clk _01279_ net985 vssd1 vssd1 vccd1 vccd1 top.a1.row2\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_74_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_82_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11280__B top.lcd.nextState\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13639_ clknet_leaf_84_clk _01225_ net1000 vssd1 vssd1 vccd1 vccd1 top.pc\[0\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__06374__B top.a1.instruction\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_210_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_805 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07160_ top.DUT.register\[28\]\[11\] net766 net726 top.DUT.register\[18\]\[11\] vssd1
+ vssd1 vccd1 vccd1 _02299_ sky130_fd_sc_hd__a22o_1
XFILLER_0_41_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_659 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_164 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_171_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07091_ top.DUT.register\[20\]\[16\] net564 net550 top.DUT.register\[18\]\[16\] vssd1
+ vssd1 vccd1 vccd1 _02230_ sky130_fd_sc_hd__a22o_1
XFILLER_0_152_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_113_2135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06390__A top.a1.instruction\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_2146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_787 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10116__S net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout206 _04823_ vssd1 vssd1 vccd1 vccd1 net206 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08763__A1 _03534_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07566__A2 net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout217 net218 vssd1 vssd1 vccd1 vccd1 net217 sky130_fd_sc_hd__buf_2
X_09801_ _04817_ _04818_ vssd1 vssd1 vccd1 vccd1 _04819_ sky130_fd_sc_hd__nand2_1
XANTENNA__08763__B2 net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout228 net230 vssd1 vssd1 vccd1 vccd1 net228 sky130_fd_sc_hd__buf_2
X_07993_ top.DUT.register\[6\]\[31\] net637 net713 top.DUT.register\[11\]\[31\] _03123_
+ vssd1 vssd1 vccd1 vccd1 _03132_ sky130_fd_sc_hd__a221o_1
XANTENNA__06774__B1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09732_ top.pc\[9\] net799 _04754_ _04758_ vssd1 vssd1 vccd1 vccd1 _04759_ sky130_fd_sc_hd__a211o_1
X_06944_ top.DUT.register\[15\]\[21\] net709 net701 top.DUT.register\[31\]\[21\] vssd1
+ vssd1 vccd1 vccd1 _02083_ sky130_fd_sc_hd__a22o_1
XFILLER_0_157_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06389__X _01528_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07318__A2 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_207_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_198_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11114__A3 net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09206__A _02678_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09663_ _04676_ _04686_ _04700_ _04701_ vssd1 vssd1 vccd1 vccd1 _04702_ sky130_fd_sc_hd__or4b_1
XANTENNA__08110__A _02286_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06526__B1 net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06875_ top.DUT.register\[3\]\[18\] net553 net462 top.DUT.register\[17\]\[18\] vssd1
+ vssd1 vccd1 vccd1 _02014_ sky130_fd_sc_hd__a22o_1
XANTENNA__13724__Q top.a1.row2\[42\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08614_ net325 _03223_ vssd1 vssd1 vccd1 vccd1 _03737_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_2_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09594_ net138 _04635_ _04640_ net133 net902 vssd1 vssd1 vccd1 vccd1 _04641_ sky130_fd_sc_hd__o221a_1
XFILLER_0_49_201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08545_ net333 _03333_ _03480_ net297 vssd1 vssd1 vccd1 vccd1 _03671_ sky130_fd_sc_hd__a22o_1
XFILLER_0_167_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10786__S net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_128_clk clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_128_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout440_A _01566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout538_A _01541_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08476_ _03381_ _03604_ net296 vssd1 vssd1 vccd1 vccd1 _03605_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09491__A2 _01896_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07427_ _02558_ _02565_ vssd1 vssd1 vccd1 vccd1 _02566_ sky130_fd_sc_hd__nor2_2
XANTENNA__09228__C1 net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout705_A _01642_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout326_X net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09876__A _03950_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07358_ _02487_ _02496_ vssd1 vssd1 vccd1 vccd1 _02497_ sky130_fd_sc_hd__nor2_4
XTAP_TAPCELL_ROW_21_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06309_ _01464_ _01461_ _01332_ vssd1 vssd1 vccd1 vccd1 _01465_ sky130_fd_sc_hd__mux2_1
XANTENNA__12567__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08451__B1 _03187_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07289_ _02421_ _02427_ vssd1 vssd1 vccd1 vccd1 _02428_ sky130_fd_sc_hd__nor2_2
XFILLER_0_143_692 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09028_ _01700_ _01744_ _04101_ _04102_ vssd1 vssd1 vccd1 vccd1 _04103_ sky130_fd_sc_hd__or4_1
XFILLER_0_142_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10026__S net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold260 top.DUT.register\[31\]\[1\] vssd1 vssd1 vccd1 vccd1 net1376 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09400__C1 net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold271 top.DUT.register\[31\]\[14\] vssd1 vssd1 vccd1 vccd1 net1387 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08004__B _03142_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold282 top.DUT.register\[14\]\[5\] vssd1 vssd1 vccd1 vccd1 net1398 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07557__A2 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold293 top.DUT.register\[19\]\[0\] vssd1 vssd1 vccd1 vccd1 net1409 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_53_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08498__Y _03626_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06765__B1 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout740 net741 vssd1 vssd1 vccd1 vccd1 net740 sky130_fd_sc_hd__buf_4
XANTENNA__08939__B _04045_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout751 _01621_ vssd1 vssd1 vccd1 vccd1 net751 sky130_fd_sc_hd__buf_2
Xfanout762 net765 vssd1 vssd1 vccd1 vccd1 net762 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_144_2607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout773 _01614_ vssd1 vssd1 vccd1 vccd1 net773 sky130_fd_sc_hd__buf_4
XANTENNA__07309__A2 net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout784 _05000_ vssd1 vssd1 vccd1 vccd1 net784 sky130_fd_sc_hd__clkbuf_2
Xfanout795 _01489_ vssd1 vssd1 vccd1 vccd1 net795 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09116__A _02952_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09703__B1 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08506__B2 net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12941_ clknet_leaf_42_clk _00533_ net1057 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[13\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06517__B1 net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12872_ clknet_leaf_26_clk _00464_ net1008 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[11\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_177_3106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11823_ _05671_ _05691_ vssd1 vssd1 vccd1 vccd1 _05706_ sky130_fd_sc_hd__xor2_4
XFILLER_0_96_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_119_clk clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_119_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__10696__S net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08809__A2 net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11754_ _05632_ _05636_ vssd1 vssd1 vccd1 vccd1 _05637_ sky130_fd_sc_hd__nand2_1
X_10705_ net2151 net232 net334 vssd1 vssd1 vccd1 vccd1 _00866_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_64_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08690__B1 _02047_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11685_ _05534_ _05563_ vssd1 vssd1 vccd1 vccd1 _05568_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_153_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13424_ clknet_leaf_23_clk _01016_ net1018 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[28\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_153_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10636_ net247 net2300 net342 vssd1 vssd1 vccd1 vccd1 _00800_ sky130_fd_sc_hd__mux2_1
XFILLER_0_180_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_155_2769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload108 clknet_leaf_60_clk vssd1 vssd1 vccd1 vccd1 clkload108/Y sky130_fd_sc_hd__inv_12
XFILLER_0_63_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13355_ clknet_leaf_46_clk _00947_ net1065 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[26\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_10567_ net1435 net256 net352 vssd1 vssd1 vccd1 vccd1 _00733_ sky130_fd_sc_hd__mux2_1
XFILLER_0_140_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12306_ top.pad.button_control.r_counter\[0\] top.pad.button_control.r_counter\[1\]
+ top.pad.button_control.r_counter\[2\] vssd1 vssd1 vccd1 vccd1 _06115_ sky130_fd_sc_hd__a21o_1
XANTENNA__07796__A2 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13286_ clknet_leaf_40_clk _00878_ net1046 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[24\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_188_3268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10498_ net1723 net265 net357 vssd1 vssd1 vccd1 vccd1 _00667_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12237_ top.lcd.cnt_20ms\[9\] top.lcd.cnt_20ms\[8\] _06069_ top.lcd.cnt_20ms\[10\]
+ vssd1 vssd1 vccd1 vccd1 _06073_ sky130_fd_sc_hd__a31o_1
XANTENNA__07548__A2 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12168_ net1271 net848 net797 _06048_ vssd1 vssd1 vccd1 vccd1 _01276_ sky130_fd_sc_hd__a22o_1
XANTENNA__06756__B1 net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_194_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11119_ net50 net868 vssd1 vssd1 vccd1 vccd1 _05065_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_207_3552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12099_ _05972_ _05978_ vssd1 vssd1 vccd1 vccd1 _05982_ sky130_fd_sc_hd__xnor2_2
Xinput6 DAT_I[13] vssd1 vssd1 vccd1 vccd1 net6 sky130_fd_sc_hd__clkbuf_1
XANTENNA__06508__B1 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06660_ _01792_ _01794_ _01796_ _01798_ vssd1 vssd1 vccd1 vccd1 _01799_ sky130_fd_sc_hd__or4_1
XFILLER_0_78_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_84_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08865__A net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07181__B1 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07720__A2 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06591_ top.DUT.register\[15\]\[28\] net709 net701 top.DUT.register\[31\]\[28\] vssd1
+ vssd1 vccd1 vccd1 _01730_ sky130_fd_sc_hd__a22o_1
XFILLER_0_176_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08330_ _03276_ _03313_ net304 vssd1 vssd1 vccd1 vccd1 _03464_ sky130_fd_sc_hd__mux2_1
XANTENNA__11265__C1 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08261_ net293 _03282_ _03396_ vssd1 vssd1 vccd1 vccd1 _03397_ sky130_fd_sc_hd__o21ai_1
XANTENNA__06287__A2 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_172_721 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09833__B1_N _04847_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12835__RESET_B net1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07212_ net894 net893 _02333_ vssd1 vssd1 vccd1 vccd1 _02351_ sky130_fd_sc_hd__o21a_1
XFILLER_0_172_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_99_1930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08192_ net321 _03329_ _03299_ vssd1 vssd1 vccd1 vccd1 _03330_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_42_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07143_ top.DUT.register\[24\]\[11\] net511 net443 top.DUT.register\[1\]\[11\] _02281_
+ vssd1 vssd1 vccd1 vccd1 _02282_ sky130_fd_sc_hd__a221o_1
XFILLER_0_125_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10240__A0 net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07787__A2 net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07074_ top.DUT.register\[23\]\[22\] net672 net652 top.DUT.register\[5\]\[22\] _02212_
+ vssd1 vssd1 vccd1 vccd1 _02213_ sky130_fd_sc_hd__a221o_1
XFILLER_0_140_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08105__A _02409_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07944__A _02070_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11674__A1_N top.a1.dataIn\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout390_A net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06747__B1 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout488_A net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07976_ top.DUT.register\[23\]\[31\] net573 net449 top.DUT.register\[21\]\[31\] _03114_
+ vssd1 vssd1 vccd1 vccd1 _03115_ sky130_fd_sc_hd__a221o_1
X_09715_ _03514_ net403 net488 _04744_ vssd1 vssd1 vccd1 vccd1 _04745_ sky130_fd_sc_hd__o211a_4
X_06927_ top.DUT.register\[12\]\[21\] net534 net529 top.DUT.register\[26\]\[21\] vssd1
+ vssd1 vccd1 vccd1 _02066_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_126_2337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout655_A _01609_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09161__A1 net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09646_ _04680_ _04684_ vssd1 vssd1 vccd1 vccd1 _04688_ sky130_fd_sc_hd__nor2_1
X_06858_ top.DUT.register\[25\]\[19\] net781 net637 top.DUT.register\[6\]\[19\] vssd1
+ vssd1 vccd1 vccd1 _01997_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_27_Left_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07172__B1 net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_182_Right_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09577_ _04606_ _04609_ _04621_ net812 vssd1 vssd1 vccd1 vccd1 _04625_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_26_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout443_X net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06789_ top.DUT.register\[30\]\[17\] net580 net571 top.DUT.register\[23\]\[17\] vssd1
+ vssd1 vccd1 vccd1 _01928_ sky130_fd_sc_hd__a22o_1
XFILLER_0_194_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08528_ net317 _03654_ _03643_ vssd1 vssd1 vccd1 vccd1 _03655_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_167_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_194_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_172_3025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08459_ _03584_ _03586_ _03588_ vssd1 vssd1 vccd1 vccd1 _03589_ sky130_fd_sc_hd__or3_1
XFILLER_0_175_570 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout610_X net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_14_Right_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout708_X net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwire415 net416 vssd1 vssd1 vccd1 vccd1 net415 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_46_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11470_ _05287_ _05319_ _05352_ _05313_ vssd1 vssd1 vccd1 vccd1 _05353_ sky130_fd_sc_hd__o22a_1
XFILLER_0_18_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_4_6__f_clk_A clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12505__RESET_B net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10421_ net1430 net174 net370 vssd1 vssd1 vccd1 vccd1 _00593_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_137_2499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_36_Left_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07778__A2 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13140_ clknet_leaf_79_clk _00732_ net1073 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[20\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_10352_ net2029 net176 net379 vssd1 vssd1 vccd1 vccd1 _00528_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13071_ clknet_leaf_41_clk _00663_ net1045 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[17\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_10283_ net1905 net202 net387 vssd1 vssd1 vccd1 vccd1 _00461_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_150_2699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12022_ _05904_ _05886_ vssd1 vssd1 vccd1 vccd1 _05905_ sky130_fd_sc_hd__and2b_1
XPHY_EDGE_ROW_23_Right_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_183_3187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_183_3198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout570 _01525_ vssd1 vssd1 vccd1 vccd1 net570 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07950__A2 _01896_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout581 _01514_ vssd1 vssd1 vccd1 vccd1 net581 sky130_fd_sc_hd__clkbuf_8
Xfanout592 _04971_ vssd1 vssd1 vccd1 vccd1 net592 sky130_fd_sc_hd__buf_4
XANTENNA__11095__B net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_45_Left_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_205_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12924_ clknet_leaf_130_clk _00516_ net910 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[13\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08685__A _02007_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06757__X _01896_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_198_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07702__A2 net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_202_3471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_202_3482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12855_ clknet_leaf_2_clk _00447_ net918 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[11\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_66_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_185_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11806_ _05681_ _05688_ _05686_ _05655_ vssd1 vssd1 vccd1 vccd1 _05689_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_84_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_32_Right_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12786_ clknet_leaf_24_clk _00378_ net1012 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[9\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_28_226 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11737_ _05603_ _05617_ _05619_ vssd1 vssd1 vccd1 vccd1 _05620_ sky130_fd_sc_hd__a21bo_2
XFILLER_0_139_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_207 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11668_ _05542_ _05549_ vssd1 vssd1 vccd1 vccd1 _05551_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_54_Left_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_181_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13407_ clknet_leaf_24_clk _00999_ net1013 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[28\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08415__B1 _03532_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11014__A2 net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10619_ net179 net1545 net347 vssd1 vssd1 vccd1 vccd1 _00784_ sky130_fd_sc_hd__mux2_1
X_11599_ net234 _05476_ _05470_ vssd1 vssd1 vccd1 vccd1 _05482_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_3_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07769__A2 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08966__B2 _04049_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13338_ clknet_leaf_1_clk _00930_ net917 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[26\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_498 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06977__B1 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_94_1860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13269_ clknet_leaf_31_clk _00861_ net1023 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[24\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_209_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_41_Right_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06729__B1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_208_232 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07830_ top.DUT.register\[22\]\[0\] net647 net746 top.DUT.register\[17\]\[0\] vssd1
+ vssd1 vccd1 vccd1 _02969_ sky130_fd_sc_hd__a22o_1
XFILLER_0_208_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_63_Left_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07761_ top.a1.instruction\[9\] _01474_ vssd1 vssd1 vccd1 vccd1 _02900_ sky130_fd_sc_hd__and2_1
X_09500_ _04537_ _04538_ _04539_ vssd1 vssd1 vccd1 vccd1 _04552_ sky130_fd_sc_hd__o21a_1
XANTENNA__09143__A1 _02857_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06712_ top.DUT.register\[21\]\[25\] net447 net443 top.DUT.register\[1\]\[25\] _01850_
+ vssd1 vssd1 vccd1 vccd1 _01851_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_108_2067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07692_ top.DUT.register\[22\]\[4\] net577 net509 top.DUT.register\[4\]\[4\] vssd1
+ vssd1 vccd1 vccd1 _02831_ sky130_fd_sc_hd__a22o_1
XFILLER_0_189_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09694__A2 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11292__Y _05182_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09431_ _02155_ _04487_ vssd1 vssd1 vccd1 vccd1 _04488_ sky130_fd_sc_hd__xor2_1
X_06643_ top.DUT.register\[10\]\[27\] net773 _01774_ _01775_ _01781_ vssd1 vssd1 vccd1
+ vccd1 _01782_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_63_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_50_Right_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06901__B1 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_121_2256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09362_ _04421_ _04422_ vssd1 vssd1 vccd1 vccd1 _04423_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_121_2267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06574_ top.DUT.register\[20\]\[28\] net565 _01712_ vssd1 vssd1 vccd1 vccd1 _01713_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_136_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08313_ _02851_ net432 net500 _02850_ _03447_ vssd1 vssd1 vccd1 vccd1 _03448_ sky130_fd_sc_hd__a221o_1
XFILLER_0_191_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09293_ net132 _04350_ _04357_ net810 vssd1 vssd1 vccd1 vccd1 _04358_ sky130_fd_sc_hd__o22a_1
XFILLER_0_145_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_11 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_72_Left_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout236_A _04757_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08244_ net306 _03380_ vssd1 vssd1 vccd1 vccd1 _03381_ sky130_fd_sc_hd__or2_1
XFILLER_0_170_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_106 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08175_ _03309_ _03312_ net289 vssd1 vssd1 vccd1 vccd1 _03313_ sky130_fd_sc_hd__mux2_1
XANTENNA__06680__A2 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout403_A net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08957__B2 net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07126_ _02264_ vssd1 vssd1 vccd1 vccd1 _02265_ sky130_fd_sc_hd__inv_2
XANTENNA__06968__B1 net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07057_ top.DUT.register\[28\]\[22\] net558 net540 top.DUT.register\[8\]\[22\] _02195_
+ vssd1 vssd1 vccd1 vccd1 _02196_ sky130_fd_sc_hd__a221o_1
XFILLER_0_140_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13804__RESET_B net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08709__A1 net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_334 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08709__B2 _03342_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout393_X net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_81_Left_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout772_A _01614_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10304__S net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07393__B1 net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07932__A2 _02632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07959_ _01702_ _03097_ vssd1 vssd1 vccd1 vccd1 _03098_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout560_X net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout658_X net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_202_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10970_ top.a1.halfData\[2\] net784 vssd1 vssd1 vccd1 vccd1 _05011_ sky130_fd_sc_hd__or2_1
XANTENNA__07145__B1 net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09629_ _04672_ _04673_ top.a1.state\[0\] _04670_ vssd1 vssd1 vccd1 vccd1 _00112_
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA_fanout825_X net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_107 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12757__RESET_B net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12640_ clknet_leaf_55_clk _00232_ net1030 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[4\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_183_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_182_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_155_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12528__Q top.pc\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_139_2528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12571_ clknet_leaf_119_clk _00163_ net930 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[2\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11244__A2 _05132_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_50_clk clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_50_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_61_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11522_ _05389_ _05404_ vssd1 vssd1 vccd1 vccd1 _05405_ sky130_fd_sc_hd__or2_1
XFILLER_0_108_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07999__A2 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_404 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_152_2728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11453_ _05287_ net278 _05299_ vssd1 vssd1 vccd1 vccd1 _05336_ sky130_fd_sc_hd__a21oi_1
X_10404_ net246 net2141 _04984_ vssd1 vssd1 vccd1 vccd1 _00576_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11384_ _05260_ _05265_ vssd1 vssd1 vccd1 vccd1 _05267_ sky130_fd_sc_hd__nand2_1
XANTENNA__06959__B1 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_185_3216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13123_ clknet_leaf_53_clk _00715_ net1038 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[19\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_185_3227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10335_ top.DUT.register\[13\]\[6\] net241 net377 vssd1 vssd1 vccd1 vccd1 _00511_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_684 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13054_ clknet_leaf_18_clk _00646_ net1027 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[17\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_10266_ net1547 net262 net388 vssd1 vssd1 vccd1 vccd1 _00444_ sky130_fd_sc_hd__mux2_1
X_12005_ _05873_ net126 _05877_ vssd1 vssd1 vccd1 vccd1 _05888_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10214__S net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10197_ net145 net2083 net393 vssd1 vssd1 vccd1 vccd1 _00377_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_204_3500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_204_3511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07136__B1 net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09676__A2 top.a1.instruction\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12907_ clknet_leaf_47_clk _00499_ net1067 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[12\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_186_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12838_ clknet_leaf_33_clk _00430_ net1046 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[10\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_196_3389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_518 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10884__S net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12769_ clknet_leaf_16_clk _00361_ net964 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[8\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_173_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_41_clk clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_41_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_123_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06290_ net879 net815 net813 net2306 net1084 vssd1 vssd1 vccd1 vccd1 _01331_ sky130_fd_sc_hd__o221a_2
XANTENNA__09677__C top.a1.instruction\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_787 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput20 DAT_I[26] vssd1 vssd1 vccd1 vccd1 net20 sky130_fd_sc_hd__clkbuf_1
XANTENNA__06662__A2 net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10185__A top.a1.instruction\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput31 DAT_I[7] vssd1 vssd1 vccd1 vccd1 net31 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06382__B top.a1.instruction\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold804 top.DUT.register\[22\]\[25\] vssd1 vssd1 vccd1 vccd1 net1920 sky130_fd_sc_hd__dlygate4sd3_1
Xhold815 top.DUT.register\[22\]\[11\] vssd1 vssd1 vccd1 vccd1 net1931 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold826 top.DUT.register\[26\]\[13\] vssd1 vssd1 vccd1 vccd1 net1942 sky130_fd_sc_hd__dlygate4sd3_1
Xhold837 top.DUT.register\[22\]\[4\] vssd1 vssd1 vccd1 vccd1 net1953 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_92_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold848 top.DUT.register\[2\]\[27\] vssd1 vssd1 vccd1 vccd1 net1964 sky130_fd_sc_hd__dlygate4sd3_1
X_09980_ net2058 net144 _04951_ vssd1 vssd1 vccd1 vccd1 _00185_ sky130_fd_sc_hd__mux2_1
Xhold859 top.DUT.register\[7\]\[16\] vssd1 vssd1 vccd1 vccd1 net1975 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07494__A _02623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08931_ _03122_ _03142_ _03187_ _03739_ _03185_ vssd1 vssd1 vccd1 vccd1 _04039_ sky130_fd_sc_hd__o311a_1
XFILLER_0_149_87 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08862_ _01833_ _03935_ _03972_ vssd1 vssd1 vccd1 vccd1 _03973_ sky130_fd_sc_hd__o21a_1
XANTENNA__10124__S net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07375__B1 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07813_ _02501_ _02951_ _01577_ vssd1 vssd1 vccd1 vccd1 _02952_ sky130_fd_sc_hd__mux2_4
X_08793_ net435 _03902_ _03907_ net424 _03904_ vssd1 vssd1 vccd1 vccd1 _03908_ sky130_fd_sc_hd__a221o_1
XFILLER_0_28_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07744_ top.DUT.register\[2\]\[3\] net561 net513 top.DUT.register\[24\]\[3\] vssd1
+ vssd1 vccd1 vccd1 _02883_ sky130_fd_sc_hd__a22o_1
XFILLER_0_196_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_211_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_189_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13732__Q top.a1.dataInTemp\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07675_ top.DUT.register\[28\]\[4\] net768 net728 top.DUT.register\[18\]\[4\] _02812_
+ vssd1 vssd1 vccd1 vccd1 _02814_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout1095_A net1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09414_ _01983_ _04471_ vssd1 vssd1 vccd1 vccd1 _04472_ sky130_fd_sc_hd__nand2_1
X_06626_ top.DUT.register\[7\]\[27\] net661 net650 top.DUT.register\[22\]\[27\] vssd1
+ vssd1 vccd1 vccd1 _01765_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_36_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_191_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09345_ _04401_ _04406_ vssd1 vssd1 vccd1 vccd1 _04407_ sky130_fd_sc_hd__xor2_1
X_06557_ top.DUT.register\[20\]\[29\] net666 _01690_ _01692_ _01695_ vssd1 vssd1 vccd1
+ vccd1 _01696_ sky130_fd_sc_hd__a2111o_1
XANTENNA__10794__S net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout520_A net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_176_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09824__C1 _04839_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout618_A _04954_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_32_clk clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_32_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_35_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_101_1959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09276_ _04334_ _04338_ _04340_ net810 vssd1 vssd1 vccd1 vccd1 _04342_ sky130_fd_sc_hd__a31o_1
XANTENNA__08117__X _03256_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06488_ net787 _01607_ _01611_ vssd1 vssd1 vccd1 vccd1 _01627_ sky130_fd_sc_hd__and3_4
XTAP_TAPCELL_ROW_43_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10985__B2 top.a1.dataIn\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08227_ _03202_ _03208_ net291 vssd1 vssd1 vccd1 vccd1 _03364_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06653__A2 net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12187__B1 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout406_X net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_200_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_134_2458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08158_ _03292_ _03295_ net293 vssd1 vssd1 vccd1 vccd1 _03296_ sky130_fd_sc_hd__mux2_1
XFILLER_0_200_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10737__A1 _04760_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout987_A net1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07109_ top.DUT.register\[5\]\[16\] net652 net736 top.DUT.register\[16\]\[16\] vssd1
+ vssd1 vccd1 vccd1 _02248_ sky130_fd_sc_hd__a22o_1
XFILLER_0_132_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06405__A2 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08089_ net331 _03040_ vssd1 vssd1 vccd1 vccd1 _03228_ sky130_fd_sc_hd__nand2_1
XFILLER_0_30_276 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10120_ net246 top.DUT.register\[7\]\[7\] net607 vssd1 vssd1 vccd1 vccd1 _00320_
+ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout775_X net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_99_clk clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_99_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__10034__S net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10051_ net1796 net257 net617 vssd1 vssd1 vccd1 vccd1 _00253_ sky130_fd_sc_hd__mux2_1
XFILLER_0_209_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08787__X _03902_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07366__B1 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_180_3146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_199_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13810_ net72 vssd1 vssd1 vccd1 vccd1 net107 sky130_fd_sc_hd__clkbuf_1
XANTENNA__07118__B1 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_202_216 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13741_ clknet_leaf_100_clk _01312_ vssd1 vssd1 vccd1 vccd1 top.lcd.cnt_20ms\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__07669__A1 top.a1.instruction\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_119_Left_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10953_ top.a1.halfData\[5\] _01425_ vssd1 vssd1 vccd1 vccd1 _04996_ sky130_fd_sc_hd__nand2_1
XFILLER_0_202_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08866__B1 net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13672_ clknet_leaf_75_clk _01248_ net1081 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[109\]
+ sky130_fd_sc_hd__dfstp_1
X_10884_ net157 top.DUT.register\[29\]\[28\] net597 vssd1 vssd1 vccd1 vccd1 _01045_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_195_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_195_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12623_ clknet_leaf_22_clk _00215_ net1033 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[3\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08618__B1 net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06892__A2 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13083__CLK clknet_leaf_120_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09778__B _04420_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_23_clk clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_23_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_14_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12554_ clknet_leaf_116_clk _00146_ net958 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[1\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10976__A1 top.a1.halfData\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11505_ _05384_ _05387_ vssd1 vssd1 vccd1 vccd1 _05388_ sky130_fd_sc_hd__nand2_1
XFILLER_0_136_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12485_ clknet_leaf_64_clk _00080_ net1092 vssd1 vssd1 vccd1 vccd1 top.ramstore\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10209__S net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11436_ _05318_ vssd1 vssd1 vccd1 vccd1 _05319_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_128_Left_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09594__A1 net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09594__B2 net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11367_ top.a1.dataIn\[31\] _05218_ vssd1 vssd1 vccd1 vccd1 _05250_ sky130_fd_sc_hd__nand2_4
XANTENNA__12920__CLK clknet_leaf_128_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_74_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_210_3592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13106_ clknet_leaf_22_clk _00698_ net1023 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[19\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_10318_ net183 net1936 net384 vssd1 vssd1 vccd1 vccd1 _00495_ sky130_fd_sc_hd__mux2_1
X_11298_ _05182_ _05185_ _05186_ vssd1 vssd1 vccd1 vccd1 _05187_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_165_2919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09346__A1 net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13037_ clknet_leaf_42_clk _00629_ net1057 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[16\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09346__B2 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10249_ net185 net2216 net391 vssd1 vssd1 vccd1 vccd1 _00428_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10879__S net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08857__B _03968_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_198_3418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07109__B1 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_2015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_89_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12608__RESET_B net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_62_clk_A clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07460_ top.DUT.register\[26\]\[15\] net751 net635 top.DUT.register\[6\]\[15\] _02598_
+ vssd1 vssd1 vccd1 vccd1 _02599_ sky130_fd_sc_hd__a221o_1
XFILLER_0_186_462 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_159_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06411_ net684 _01512_ _01521_ vssd1 vssd1 vccd1 vccd1 _01550_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_33_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07391_ top.DUT.register\[2\]\[9\] net559 net546 top.DUT.register\[16\]\[9\] vssd1
+ vssd1 vccd1 vccd1 _02530_ sky130_fd_sc_hd__a22o_1
XANTENNA__06883__A2 net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_14_clk clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_14_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_84_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_151_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09130_ net889 net899 vssd1 vssd1 vccd1 vccd1 _04205_ sky130_fd_sc_hd__nand2_1
XFILLER_0_84_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06342_ _01389_ _01473_ vssd1 vssd1 vccd1 vccd1 _01484_ sky130_fd_sc_hd__nand2_1
XFILLER_0_56_173 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08084__S net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_77_clk_A clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09061_ _03791_ _04135_ _03854_ _03772_ vssd1 vssd1 vccd1 vccd1 _04136_ sky130_fd_sc_hd__or4b_1
XFILLER_0_60_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06635__A2 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10119__S net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06273_ top.lcd.cnt_500hz\[1\] top.lcd.cnt_500hz\[0\] top.lcd.cnt_500hz\[3\] top.lcd.cnt_500hz\[2\]
+ vssd1 vssd1 vccd1 vccd1 _01436_ sky130_fd_sc_hd__and4_1
XFILLER_0_127_595 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_120_clk_A clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08012_ _01392_ net893 _03148_ _01391_ vssd1 vssd1 vccd1 vccd1 _03151_ sky130_fd_sc_hd__a31o_2
XFILLER_0_130_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold601 top.DUT.register\[14\]\[28\] vssd1 vssd1 vccd1 vccd1 net1717 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold612 top.DUT.register\[12\]\[12\] vssd1 vssd1 vccd1 vccd1 net1728 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_116_2188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold623 top.DUT.register\[1\]\[24\] vssd1 vssd1 vccd1 vccd1 net1739 sky130_fd_sc_hd__dlygate4sd3_1
Xhold634 top.DUT.register\[20\]\[31\] vssd1 vssd1 vccd1 vccd1 net1750 sky130_fd_sc_hd__dlygate4sd3_1
Xhold645 top.DUT.register\[26\]\[10\] vssd1 vssd1 vccd1 vccd1 net1761 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold656 top.DUT.register\[12\]\[28\] vssd1 vssd1 vccd1 vccd1 net1772 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07596__B1 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_788 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold667 top.DUT.register\[29\]\[19\] vssd1 vssd1 vccd1 vccd1 net1783 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_95 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07428__S net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09963_ net2030 net204 net630 vssd1 vssd1 vccd1 vccd1 _00171_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_4_Right_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold678 top.DUT.register\[8\]\[23\] vssd1 vssd1 vccd1 vccd1 net1794 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08113__A _02544_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold689 top.DUT.register\[29\]\[12\] vssd1 vssd1 vccd1 vccd1 net1805 sky130_fd_sc_hd__dlygate4sd3_1
X_08914_ _01659_ net493 _03184_ _01658_ vssd1 vssd1 vccd1 vccd1 _04023_ sky130_fd_sc_hd__a2bb2o_1
X_09894_ net828 _04589_ vssd1 vssd1 vccd1 vccd1 _04903_ sky130_fd_sc_hd__nor2_1
XANTENNA_clkbuf_leaf_15_clk_A clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08845_ _03916_ _03956_ net287 vssd1 vssd1 vccd1 vccd1 _03957_ sky130_fd_sc_hd__mux2_1
XANTENNA__08400__X _03532_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10789__S net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout568_A _01525_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08776_ net1298 net830 net800 _03891_ vssd1 vssd1 vccd1 vccd1 _00041_ sky130_fd_sc_hd__a22o_1
X_07727_ top.DUT.register\[28\]\[3\] net767 net704 top.DUT.register\[3\]\[3\] vssd1
+ vssd1 vccd1 vccd1 _02866_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout735_A net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout356_X net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1098_X net1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07658_ _02796_ vssd1 vssd1 vccd1 vccd1 _02797_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_45_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_45_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06609_ top.DUT.register\[14\]\[27\] net586 net557 top.DUT.register\[28\]\[27\] vssd1
+ vssd1 vccd1 vccd1 _01748_ sky130_fd_sc_hd__a22o_1
XFILLER_0_177_484 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06874__A2 net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout523_X net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07589_ top.a1.instruction\[27\] net805 _02727_ vssd1 vssd1 vccd1 vccd1 _02728_ sky130_fd_sc_hd__a21oi_2
XANTENNA_fanout902_A net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09328_ _04372_ _04390_ vssd1 vssd1 vccd1 vccd1 _04391_ sky130_fd_sc_hd__and2_1
XFILLER_0_118_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_11_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11255__A_N top.lcd.nextState\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06626__A2 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09259_ net898 top.pc\[10\] _04325_ net889 vssd1 vssd1 vccd1 vccd1 _00090_ sky130_fd_sc_hd__o211a_1
XFILLER_0_7_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10029__S net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12270_ net686 _06092_ vssd1 vssd1 vccd1 vccd1 _01340_ sky130_fd_sc_hd__and2_1
XFILLER_0_90_496 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout892_X net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13137__RESET_B net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11221_ _05116_ net1201 net471 vssd1 vssd1 vccd1 vccd1 _01261_ sky130_fd_sc_hd__mux2_1
XANTENNA__09576__A1 net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11152_ _04657_ net848 vssd1 vssd1 vccd1 vccd1 _05082_ sky130_fd_sc_hd__nor2_2
XANTENNA__07051__A2 net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10103_ net1474 net179 net611 vssd1 vssd1 vccd1 vccd1 _00304_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11083_ net51 net867 vssd1 vssd1 vccd1 vccd1 _05047_ sky130_fd_sc_hd__and2_1
XANTENNA_input31_A DAT_I[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_147_2649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10034_ net2148 net201 net621 vssd1 vssd1 vccd1 vccd1 _00237_ sky130_fd_sc_hd__mux2_1
XANTENNA__10699__S net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_160_2849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11985_ _05847_ _05849_ _05840_ vssd1 vssd1 vccd1 vccd1 _05868_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_105_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_187_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13724_ clknet_leaf_95_clk _01295_ net986 vssd1 vssd1 vccd1 vccd1 top.a1.row2\[42\]
+ sky130_fd_sc_hd__dfrtp_1
X_10936_ net1658 net226 net591 vssd1 vssd1 vccd1 vccd1 _01097_ sky130_fd_sc_hd__mux2_1
XFILLER_0_168_451 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07511__B1 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_193_3337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_193_3348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10867_ net221 net1830 net594 vssd1 vssd1 vccd1 vccd1 _01028_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13655_ clknet_leaf_93_clk _00013_ net994 vssd1 vssd1 vccd1 vccd1 wb.curr_state\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_155_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_171_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12606_ clknet_leaf_52_clk _00198_ net1037 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[3\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_13586_ clknet_leaf_64_clk net1200 net1092 vssd1 vssd1 vccd1 vccd1 net77 sky130_fd_sc_hd__dfrtp_1
X_10798_ net242 net1747 net598 vssd1 vssd1 vccd1 vccd1 _00959_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06617__A2 net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12537_ clknet_leaf_13_clk _00129_ net942 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[1\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_152_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12468_ clknet_leaf_63_clk _00063_ net1092 vssd1 vssd1 vccd1 vccd1 top.ramstore\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07290__A2 _02428_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11419_ _05264_ _05300_ vssd1 vssd1 vccd1 vccd1 _05302_ sky130_fd_sc_hd__xnor2_2
X_12399_ clknet_leaf_104_clk top.ru.next_FetchedInstr\[11\] net972 vssd1 vssd1 vccd1
+ vccd1 top.a1.instruction\[11\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__07578__B1 net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07042__A2 net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_190_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06960_ top.DUT.register\[25\]\[23\] net458 net448 top.DUT.register\[21\]\[23\] vssd1
+ vssd1 vccd1 vccd1 _02099_ sky130_fd_sc_hd__a22o_1
XFILLER_0_39_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_3_clk clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_3_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__11126__A1 net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06891_ top.DUT.register\[15\]\[18\] net708 net700 top.DUT.register\[31\]\[18\] vssd1
+ vssd1 vccd1 vccd1 _02030_ sky130_fd_sc_hd__a22o_1
X_08630_ _01964_ net492 vssd1 vssd1 vccd1 vccd1 _03752_ sky130_fd_sc_hd__nor2_1
XFILLER_0_179_705 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10402__S net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08561_ _03240_ _03244_ vssd1 vssd1 vccd1 vccd1 _03686_ sky130_fd_sc_hd__and2_1
XFILLER_0_77_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07512_ _02646_ _02648_ _02650_ vssd1 vssd1 vccd1 vccd1 _02651_ sky130_fd_sc_hd__or3_1
XANTENNA__09699__A _04716_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08492_ _02310_ _03619_ vssd1 vssd1 vccd1 vccd1 _03620_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07502__B1 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_193_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_159_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07443_ top.DUT.register\[11\]\[15\] net524 _02581_ vssd1 vssd1 vccd1 vccd1 _02582_
+ sky130_fd_sc_hd__a21o_1
XANTENNA__06856__A2 net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout149_A _04938_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07374_ _02506_ _02509_ _02510_ _02512_ vssd1 vssd1 vccd1 vccd1 _02513_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_118_2217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09113_ _04184_ _04187_ vssd1 vssd1 vccd1 vccd1 _04188_ sky130_fd_sc_hd__xnor2_1
X_06325_ top.a1.instruction\[2\] top.a1.instruction\[3\] top.a1.instruction\[0\] top.a1.instruction\[1\]
+ vssd1 vssd1 vccd1 vccd1 _01472_ sky130_fd_sc_hd__or4bb_2
XFILLER_0_95_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06608__A2 net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout316_A _02880_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1058_A net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09044_ _04115_ _04118_ _04079_ _04112_ vssd1 vssd1 vccd1 vccd1 _04119_ sky130_fd_sc_hd__o211a_1
X_06256_ net1278 net852 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedData\[17\] sky130_fd_sc_hd__and2_1
XANTENNA__07281__A2 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_2406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_2417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold420 top.DUT.register\[2\]\[30\] vssd1 vssd1 vccd1 vccd1 net1536 sky130_fd_sc_hd__dlygate4sd3_1
X_06187_ net888 _01413_ vssd1 vssd1 vccd1 vccd1 _01425_ sky130_fd_sc_hd__nor2_1
Xhold431 top.DUT.register\[11\]\[3\] vssd1 vssd1 vccd1 vccd1 net1547 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07569__B1 net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold442 top.DUT.register\[28\]\[12\] vssd1 vssd1 vccd1 vccd1 net1558 sky130_fd_sc_hd__dlygate4sd3_1
Xhold453 top.DUT.register\[4\]\[8\] vssd1 vssd1 vccd1 vccd1 net1569 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07033__A2 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold464 top.DUT.register\[16\]\[9\] vssd1 vssd1 vccd1 vccd1 net1580 sky130_fd_sc_hd__dlygate4sd3_1
Xhold475 top.DUT.register\[18\]\[1\] vssd1 vssd1 vccd1 vccd1 net1591 sky130_fd_sc_hd__dlygate4sd3_1
Xhold486 top.DUT.register\[1\]\[16\] vssd1 vssd1 vccd1 vccd1 net1602 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12361__Q top.a1.dataIn\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout900 net903 vssd1 vssd1 vccd1 vccd1 net900 sky130_fd_sc_hd__clkbuf_4
Xfanout911 net913 vssd1 vssd1 vccd1 vccd1 net911 sky130_fd_sc_hd__clkbuf_4
Xhold497 top.DUT.register\[10\]\[17\] vssd1 vssd1 vccd1 vccd1 net1613 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout922 net935 vssd1 vssd1 vccd1 vccd1 net922 sky130_fd_sc_hd__clkbuf_2
X_09946_ net1526 net269 net629 vssd1 vssd1 vccd1 vccd1 _00154_ sky130_fd_sc_hd__mux2_1
Xfanout933 net934 vssd1 vssd1 vccd1 vccd1 net933 sky130_fd_sc_hd__clkbuf_4
Xfanout944 net952 vssd1 vssd1 vccd1 vccd1 net944 sky130_fd_sc_hd__clkbuf_4
Xfanout955 net956 vssd1 vssd1 vccd1 vccd1 net955 sky130_fd_sc_hd__clkbuf_4
Xfanout966 net967 vssd1 vssd1 vccd1 vccd1 net966 sky130_fd_sc_hd__clkbuf_2
Xfanout977 net1007 vssd1 vssd1 vccd1 vccd1 net977 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08130__X _03269_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout852_A net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout473_X net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1120 top.ramstore\[5\] vssd1 vssd1 vccd1 vccd1 net2236 sky130_fd_sc_hd__dlygate4sd3_1
X_09877_ top.pc\[26\] _04577_ vssd1 vssd1 vccd1 vccd1 _04887_ sky130_fd_sc_hd__and2_1
XANTENNA__08497__B _03427_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout988 net990 vssd1 vssd1 vccd1 vccd1 net988 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_129_2379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1131 top.DUT.register\[13\]\[30\] vssd1 vssd1 vccd1 vccd1 net2247 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout999 net1000 vssd1 vssd1 vccd1 vccd1 net999 sky130_fd_sc_hd__clkbuf_4
Xhold1142 top.DUT.register\[3\]\[5\] vssd1 vssd1 vccd1 vccd1 net2258 sky130_fd_sc_hd__dlygate4sd3_1
X_08828_ net274 _03775_ _03940_ vssd1 vssd1 vccd1 vccd1 _03941_ sky130_fd_sc_hd__a21o_1
Xhold1153 top.DUT.register\[8\]\[6\] vssd1 vssd1 vccd1 vccd1 net2269 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10312__S net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1164 top.DUT.register\[2\]\[21\] vssd1 vssd1 vccd1 vccd1 net2280 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07741__A0 _02857_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1175 top.DUT.register\[23\]\[10\] vssd1 vssd1 vccd1 vccd1 net2291 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_79_Right_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1186 top.a1.row2\[35\] vssd1 vssd1 vccd1 vccd1 net2302 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_197_535 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08759_ _03836_ _03874_ net287 vssd1 vssd1 vccd1 vccd1 _03875_ sky130_fd_sc_hd__mux2_1
Xhold1197 top.ramload\[10\] vssd1 vssd1 vccd1 vccd1 net2313 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout640_X net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout738_X net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_197_568 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_142_2579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11770_ _05606_ _05633_ vssd1 vssd1 vccd1 vccd1 _05653_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_178_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10721_ net1971 net168 net334 vssd1 vssd1 vccd1 vccd1 _00882_ sky130_fd_sc_hd__mux2_1
XANTENNA__06847__A2 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout905_X net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_175_3067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_175_3078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08049__A1 _03177_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13440_ clknet_leaf_113_clk _01032_ net992 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[29\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_192_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10652_ net177 net1968 net344 vssd1 vssd1 vccd1 vccd1 _00816_ sky130_fd_sc_hd__mux2_1
XFILLER_0_193_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09797__A1 _04453_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13371_ clknet_leaf_124_clk _00963_ net925 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[27\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09797__B2 top.a1.dataIn\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10583_ net1762 net200 net352 vssd1 vssd1 vccd1 vccd1 _00749_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12322_ top.pad.button_control.r_counter\[7\] top.pad.button_control.r_counter\[6\]
+ _06120_ top.pad.button_control.r_counter\[8\] vssd1 vssd1 vccd1 vccd1 _06125_ sky130_fd_sc_hd__a31o_1
XPHY_EDGE_ROW_88_Right_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07857__A _02974_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07272__A2 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12253_ top.lcd.cnt_20ms\[15\] top.lcd.cnt_20ms\[14\] _06079_ top.lcd.cnt_20ms\[16\]
+ vssd1 vssd1 vccd1 vccd1 _06083_ sky130_fd_sc_hd__a31o_1
X_11204_ _05108_ net1251 net471 vssd1 vssd1 vccd1 vccd1 _01252_ sky130_fd_sc_hd__mux2_1
XANTENNA__07024__A2 net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12184_ net797 _05758_ _05787_ net847 net2302 vssd1 vssd1 vccd1 vccd1 _01292_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_71_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11135_ net59 net869 vssd1 vssd1 vccd1 vccd1 _05073_ sky130_fd_sc_hd__and2_1
XFILLER_0_101_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_207_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11108__A1 net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_196_Right_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07980__B1 net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input34_X net34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11066_ net81 net870 net834 net1139 vssd1 vssd1 vccd1 vccd1 _01177_ sky130_fd_sc_hd__a22o_1
XFILLER_0_207_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_97_Right_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10017_ net2088 net260 net620 vssd1 vssd1 vccd1 vccd1 _00220_ sky130_fd_sc_hd__mux2_1
XANTENNA__10222__S net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07732__B1 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_86_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_382 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08288__A1 _03342_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08288__B2 net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_175_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11968_ _05847_ _05849_ vssd1 vssd1 vccd1 vccd1 _05851_ sky130_fd_sc_hd__and2_1
XFILLER_0_156_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13707_ clknet_leaf_96_clk _01278_ net985 vssd1 vssd1 vccd1 vccd1 top.a1.row2\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06838__A2 net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10919_ net1642 net141 net480 vssd1 vssd1 vccd1 vccd1 _01080_ sky130_fd_sc_hd__mux2_1
X_11899_ _05737_ _05764_ vssd1 vssd1 vccd1 vccd1 _05782_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_46_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07103__Y _02242_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11280__C _05148_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13638_ clknet_leaf_71_clk _01224_ vssd1 vssd1 vccd1 vccd1 top.lcd.nextState\[3\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_184_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_167 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10892__S net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_817 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13569_ clknet_leaf_104_clk _01156_ net972 vssd1 vssd1 vccd1 vccd1 top.ramload\[30\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_125_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07799__B1 net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_203_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_176 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_340 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08460__A1 net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07090_ top.DUT.register\[4\]\[16\] net508 net440 top.DUT.register\[5\]\[16\] _02228_
+ vssd1 vssd1 vccd1 vccd1 _02229_ sky130_fd_sc_hd__a221o_1
XANTENNA__07263__A2 net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06671__A _01809_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08215__X _03353_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08460__B2 net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10193__A net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_2136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_2147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06390__B top.a1.instruction\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08869__Y _03980_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09960__A1 net191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09800_ top.pc\[18\] _04453_ vssd1 vssd1 vccd1 vccd1 _04818_ sky130_fd_sc_hd__or2_1
Xfanout207 net210 vssd1 vssd1 vccd1 vccd1 net207 sky130_fd_sc_hd__clkbuf_2
Xfanout218 _04814_ vssd1 vssd1 vccd1 vccd1 net218 sky130_fd_sc_hd__clkbuf_2
Xfanout229 net230 vssd1 vssd1 vccd1 vccd1 net229 sky130_fd_sc_hd__buf_2
X_07992_ top.DUT.register\[20\]\[31\] net665 net645 top.DUT.register\[24\]\[31\] _03128_
+ vssd1 vssd1 vccd1 vccd1 _03131_ sky130_fd_sc_hd__a221o_1
XFILLER_0_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07971__B1 net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06943_ top.DUT.register\[2\]\[21\] net745 net725 top.DUT.register\[29\]\[21\] _02081_
+ vssd1 vssd1 vccd1 vccd1 _02082_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_163_Right_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09731_ net826 _04297_ _04752_ top.a1.dataIn\[9\] vssd1 vssd1 vccd1 vccd1 _04758_
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_207_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10132__S net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09662_ _04674_ _04681_ _04684_ _04678_ vssd1 vssd1 vccd1 vccd1 _04701_ sky130_fd_sc_hd__o22a_1
X_06874_ top.DUT.register\[30\]\[18\] net581 net449 top.DUT.register\[21\]\[18\] _02012_
+ vssd1 vssd1 vccd1 vccd1 _02013_ sky130_fd_sc_hd__a221o_1
XANTENNA__07723__B1 net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08613_ _03175_ _03534_ _03735_ vssd1 vssd1 vccd1 vccd1 _03736_ sky130_fd_sc_hd__o21ai_2
X_09593_ _04636_ _04639_ vssd1 vssd1 vccd1 vccd1 _04640_ sky130_fd_sc_hd__xor2_1
XANTENNA__11174__D _05082_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout266_A _04729_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08544_ net281 _03464_ _03468_ net275 vssd1 vssd1 vccd1 vccd1 _03670_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_49_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_210_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08475_ _03603_ vssd1 vssd1 vccd1 vccd1 _03604_ sky130_fd_sc_hd__inv_2
XANTENNA__06829__A2 net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_175_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout433_A _03184_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07426_ _02560_ _02562_ _02564_ vssd1 vssd1 vccd1 vccd1 _02565_ sky130_fd_sc_hd__or3_1
XFILLER_0_174_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13144__CLK clknet_leaf_128_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12356__Q top.a1.dataIn\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_603 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07357_ _02491_ _02493_ _02495_ vssd1 vssd1 vccd1 vccd1 _02496_ sky130_fd_sc_hd__or3_1
XFILLER_0_190_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout600_A net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09876__B _04716_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_190_766 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout319_X net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_636 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06308_ _01459_ _01463_ vssd1 vssd1 vccd1 vccd1 _01464_ sky130_fd_sc_hd__or2_1
XFILLER_0_131_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07254__A2 net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07288_ _02423_ _02425_ _02426_ vssd1 vssd1 vccd1 vccd1 _02427_ sky130_fd_sc_hd__or3_1
XANTENNA__08125__X _03264_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09027_ _01787_ _01832_ _01919_ _02005_ vssd1 vssd1 vccd1 vccd1 _04102_ sky130_fd_sc_hd__or4b_1
X_06239_ top.ramload\[0\] net855 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedData\[0\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_103_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10307__S net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold250 top.DUT.register\[8\]\[3\] vssd1 vssd1 vccd1 vccd1 net1366 sky130_fd_sc_hd__dlygate4sd3_1
Xhold261 top.DUT.register\[19\]\[28\] vssd1 vssd1 vccd1 vccd1 net1377 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold272 top.DUT.register\[18\]\[28\] vssd1 vssd1 vccd1 vccd1 net1388 sky130_fd_sc_hd__dlygate4sd3_1
Xhold283 top.DUT.register\[25\]\[27\] vssd1 vssd1 vccd1 vccd1 net1399 sky130_fd_sc_hd__dlygate4sd3_1
Xhold294 top.DUT.register\[24\]\[12\] vssd1 vssd1 vccd1 vccd1 net1410 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_53_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout730 _01627_ vssd1 vssd1 vccd1 vccd1 net730 sky130_fd_sc_hd__buf_4
XANTENNA__12364__RESET_B net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout741 _01624_ vssd1 vssd1 vccd1 vccd1 net741 sky130_fd_sc_hd__clkbuf_4
X_09929_ net828 _04635_ vssd1 vssd1 vccd1 vccd1 _04935_ sky130_fd_sc_hd__nor2_1
Xfanout752 _01621_ vssd1 vssd1 vccd1 vccd1 net752 sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_130_Right_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout763 net765 vssd1 vssd1 vccd1 vccd1 net763 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_144_2608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout855_X net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout774 net777 vssd1 vssd1 vccd1 vccd1 net774 sky130_fd_sc_hd__clkbuf_8
Xfanout785 _04999_ vssd1 vssd1 vccd1 vccd1 net785 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09703__A1 top.a1.dataIn\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08506__A2 net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout796 net797 vssd1 vssd1 vccd1 vccd1 net796 sky130_fd_sc_hd__buf_2
XFILLER_0_99_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10042__S net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12940_ clknet_leaf_60_clk _00532_ net1089 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[13\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09116__B _02994_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06517__A1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08969__A1_N net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12871_ clknet_leaf_6_clk _00463_ net938 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[11\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_177_3107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_29_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11822_ _05698_ _05703_ _05704_ vssd1 vssd1 vccd1 vccd1 _05705_ sky130_fd_sc_hd__a21boi_4
XTAP_TAPCELL_ROW_68_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11753_ _05608_ _05635_ vssd1 vssd1 vccd1 vccd1 _05636_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_68_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13650__Q top.a1.row1\[58\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10704_ net1626 net238 net337 vssd1 vssd1 vccd1 vccd1 _00865_ sky130_fd_sc_hd__mux2_1
XANTENNA__08690__A1 _01983_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11684_ _05557_ _05560_ _05562_ _05563_ _05564_ vssd1 vssd1 vccd1 vccd1 _05567_ sky130_fd_sc_hd__a2111o_1
X_10635_ net244 net2232 net342 vssd1 vssd1 vccd1 vccd1 _00799_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13423_ clknet_leaf_21_clk _01015_ net1033 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[28\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_181_755 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkload109 clknet_leaf_65_clk vssd1 vssd1 vccd1 vccd1 clkload109/Y sky130_fd_sc_hd__inv_6
XFILLER_0_23_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13354_ clknet_leaf_117_clk _00946_ net958 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[26\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_63_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10566_ net2133 net260 net351 vssd1 vssd1 vccd1 vccd1 _00732_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12305_ top.pad.button_control.r_counter\[0\] top.pad.button_control.r_counter\[2\]
+ top.pad.button_control.r_counter\[1\] vssd1 vssd1 vccd1 vccd1 _06114_ sky130_fd_sc_hd__and3_1
XFILLER_0_23_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10217__S net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13285_ clknet_leaf_34_clk _00877_ net1043 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[24\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_10497_ net1591 net270 net358 vssd1 vssd1 vccd1 vccd1 _00666_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_188_3269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12236_ net1240 _06070_ _06072_ vssd1 vssd1 vccd1 vccd1 _01320_ sky130_fd_sc_hd__a21oi_1
X_12167_ _06041_ _06047_ vssd1 vssd1 vccd1 vccd1 _06048_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_9_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11118_ net908 net2315 net863 _05064_ vssd1 vssd1 vccd1 vccd1 _01210_ sky130_fd_sc_hd__a31o_1
XANTENNA__09307__A _02399_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12098_ _05980_ vssd1 vssd1 vccd1 vccd1 _05981_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_207_3553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11049_ net1242 net872 net836 top.ramstore\[0\] vssd1 vssd1 vccd1 vccd1 _01160_ sky130_fd_sc_hd__a22o_1
XANTENNA__07705__B1 net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput7 DAT_I[14] vssd1 vssd1 vccd1 vccd1 net7 sky130_fd_sc_hd__clkbuf_1
XANTENNA__10887__S net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06590_ top.DUT.register\[1\]\[28\] net757 net720 top.DUT.register\[19\]\[28\] vssd1
+ vssd1 vccd1 vccd1 _01729_ sky130_fd_sc_hd__a22o_1
XFILLER_0_59_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13560__Q top.ramload\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08260_ net293 _03292_ vssd1 vssd1 vccd1 vccd1 _03396_ sky130_fd_sc_hd__nand2_1
XANTENNA__09977__A _04155_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08681__A1 _02007_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08681__B2 _03258_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07211_ _01486_ _02336_ vssd1 vssd1 vccd1 vccd1 _02350_ sky130_fd_sc_hd__or2_1
XANTENNA__11017__B1 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08191_ _03314_ _03328_ net316 vssd1 vssd1 vccd1 vccd1 _03329_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_99_1931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07142_ top.DUT.register\[3\]\[11\] net551 net447 top.DUT.register\[21\]\[11\] vssd1
+ vssd1 vccd1 vccd1 _02281_ sky130_fd_sc_hd__a22o_1
XANTENNA__08433__A1 _03263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07236__A2 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07073_ top.DUT.register\[9\]\[22\] net762 net743 top.DUT.register\[2\]\[22\] vssd1
+ vssd1 vccd1 vccd1 _02212_ sky130_fd_sc_hd__a22o_1
XFILLER_0_112_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_488 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10127__S net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07975_ top.DUT.register\[14\]\[31\] net585 net446 top.DUT.register\[1\]\[31\] vssd1
+ vssd1 vccd1 vccd1 _03114_ sky130_fd_sc_hd__a22o_1
XANTENNA__08121__A _03151_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout383_A net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09146__C1 _01393_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06926_ top.DUT.register\[3\]\[21\] net554 net461 top.DUT.register\[17\]\[21\] _02064_
+ vssd1 vssd1 vccd1 vccd1 _02065_ sky130_fd_sc_hd__a221o_1
X_09714_ net407 _04743_ vssd1 vssd1 vccd1 vccd1 _04744_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_126_2338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06857_ top.DUT.register\[14\]\[19\] net733 _01993_ _01995_ vssd1 vssd1 vccd1 vccd1
+ _01996_ sky130_fd_sc_hd__a211o_1
X_09645_ _04678_ _04681_ vssd1 vssd1 vccd1 vccd1 _04687_ sky130_fd_sc_hd__nor2_1
XANTENNA__10797__S net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_195_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout648_A _01612_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09576_ net138 _04613_ _04204_ vssd1 vssd1 vccd1 vccd1 _04624_ sky130_fd_sc_hd__o21a_1
X_06788_ top.DUT.register\[22\]\[17\] net575 net465 top.DUT.register\[13\]\[17\] _01926_
+ vssd1 vssd1 vccd1 vccd1 _01927_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_26_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08527_ net298 _03122_ _03371_ _03644_ vssd1 vssd1 vccd1 vccd1 _03654_ sky130_fd_sc_hd__o211a_1
XFILLER_0_65_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout436_X net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout815_A _01442_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_203_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08706__A2_N net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10529__C net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08458_ net298 _03587_ vssd1 vssd1 vccd1 vccd1 _03588_ sky130_fd_sc_hd__nor2_1
XFILLER_0_163_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09887__A _03968_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_172_3026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_582 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07409_ top.DUT.register\[15\]\[9\] net706 net698 top.DUT.register\[31\]\[9\] vssd1
+ vssd1 vccd1 vccd1 _02548_ sky130_fd_sc_hd__a22o_1
XANTENNA__06683__B1 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout603_X net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwire416 net417 vssd1 vssd1 vccd1 vccd1 net416 sky130_fd_sc_hd__clkbuf_2
X_08389_ _02752_ _03509_ _02751_ vssd1 vssd1 vccd1 vccd1 _03521_ sky130_fd_sc_hd__o21bai_1
XANTENNA__06582__Y _01721_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_580 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10420_ net1353 net178 net369 vssd1 vssd1 vccd1 vccd1 _00592_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_619 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07227__A2 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10351_ net1605 net182 net377 vssd1 vssd1 vccd1 vccd1 _00527_ sky130_fd_sc_hd__mux2_1
XANTENNA__10037__S net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09826__S net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13070_ clknet_leaf_39_clk _00662_ net1055 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[17\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_10282_ net1375 net187 net387 vssd1 vssd1 vccd1 vccd1 _00460_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_150_2689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12021_ _05893_ _05894_ _05895_ _05900_ _05903_ vssd1 vssd1 vccd1 vccd1 _05904_ sky130_fd_sc_hd__o41a_2
XANTENNA__08302__Y _03437_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08031__A net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_183_3188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout560 _01532_ vssd1 vssd1 vccd1 vccd1 net560 sky130_fd_sc_hd__buf_2
XFILLER_0_205_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout571 _01519_ vssd1 vssd1 vccd1 vccd1 net571 sky130_fd_sc_hd__clkbuf_8
Xfanout582 _01514_ vssd1 vssd1 vccd1 vccd1 net582 sky130_fd_sc_hd__clkbuf_4
Xfanout593 _04971_ vssd1 vssd1 vccd1 vccd1 net593 sky130_fd_sc_hd__buf_6
XANTENNA__09688__B1 net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09152__A2 _02904_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_100_Left_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12923_ clknet_leaf_124_clk _00515_ net923 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[13\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_186_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_201_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_202_3472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10500__S net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12854_ clknet_leaf_3_clk _00446_ net940 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[11\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_202_3483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_197_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11805_ _05684_ _05687_ vssd1 vssd1 vccd1 vccd1 _05688_ sky130_fd_sc_hd__nand2_1
X_12785_ clknet_leaf_113_clk _00377_ net991 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[9\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11736_ _05610_ _05616_ _05618_ _05613_ _05580_ vssd1 vssd1 vccd1 vccd1 _05619_ sky130_fd_sc_hd__o32a_1
XANTENNA__07466__A2 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06674__B1 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11667_ _01398_ _05549_ vssd1 vssd1 vccd1 vccd1 _05550_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_83_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_181_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13406_ clknet_leaf_18_clk _00998_ net1027 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[28\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_141_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08415__A1 net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10618_ net180 net2176 net347 vssd1 vssd1 vccd1 vccd1 _00783_ sky130_fd_sc_hd__mux2_1
XFILLER_0_113_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08415__B2 _03258_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11598_ net234 _05476_ _05462_ vssd1 vssd1 vccd1 vccd1 _05481_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_12_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08966__A2 net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10549_ net2244 net184 net355 vssd1 vssd1 vccd1 vccd1 _00716_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13337_ clknet_leaf_11_clk _00929_ net951 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[26\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_94_1850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_1861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13268_ clknet_4_12__leaf_clk _00860_ net1075 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[24\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_12219_ _06059_ _06062_ net980 vssd1 vssd1 vccd1 vccd1 _01313_ sky130_fd_sc_hd__o21a_1
X_13199_ clknet_leaf_22_clk _00791_ net1022 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[21\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_209_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_209_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_208_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_208_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07760_ _02889_ _02898_ vssd1 vssd1 vccd1 vccd1 _02899_ sky130_fd_sc_hd__nor2_4
X_06711_ top.DUT.register\[26\]\[25\] net530 net511 top.DUT.register\[24\]\[25\] vssd1
+ vssd1 vccd1 vccd1 _01850_ sky130_fd_sc_hd__a22o_1
XFILLER_0_79_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_108_2068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07691_ net824 _02808_ _02828_ vssd1 vssd1 vccd1 vccd1 _02830_ sky130_fd_sc_hd__o21ai_4
X_09430_ net820 _02330_ net422 vssd1 vssd1 vccd1 vccd1 _04487_ sky130_fd_sc_hd__o21bai_4
XFILLER_0_78_127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06642_ top.DUT.register\[8\]\[27\] net642 _01765_ _01778_ _01780_ vssd1 vssd1 vccd1
+ vccd1 _01781_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_149_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10410__S net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06396__A top.a1.instruction\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09361_ _02232_ _02241_ _04420_ vssd1 vssd1 vccd1 vccd1 _04422_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_121_2257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06573_ top.DUT.register\[15\]\[28\] net682 net678 top.DUT.register\[31\]\[28\] vssd1
+ vssd1 vccd1 vccd1 _01712_ sky130_fd_sc_hd__a22o_1
XFILLER_0_47_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_121_2268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08312_ _02852_ net492 vssd1 vssd1 vccd1 vccd1 _03447_ sky130_fd_sc_hd__nor2_1
X_09292_ _04355_ _04356_ vssd1 vssd1 vccd1 vccd1 _04357_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07457__A2 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06382__A_N top.a1.instruction\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08243_ _03172_ _03378_ net291 vssd1 vssd1 vccd1 vccd1 _03380_ sky130_fd_sc_hd__mux2_1
XANTENNA__06665__B1 net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_1990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_172_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout229_A net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08174_ _03310_ _03311_ vssd1 vssd1 vccd1 vccd1 _03312_ sky130_fd_sc_hd__nand2_1
XFILLER_0_172_574 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_118 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06417__B1 net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07125_ _02242_ _02261_ vssd1 vssd1 vccd1 vccd1 _02264_ sky130_fd_sc_hd__nand2_1
XFILLER_0_88_50 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07056_ top.DUT.register\[30\]\[22\] net580 net571 top.DUT.register\[23\]\[22\] vssd1
+ vssd1 vccd1 vccd1 _02195_ sky130_fd_sc_hd__a22o_1
XANTENNA__07090__B1 net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout598_A _04965_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09367__C1 net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09906__A1 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_346 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout386_X net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07958_ _01722_ _01742_ _03096_ vssd1 vssd1 vccd1 vccd1 _03097_ sky130_fd_sc_hd__a21oi_1
X_06909_ _02026_ _02046_ vssd1 vssd1 vccd1 vccd1 _02048_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout553_X net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07889_ top.DUT.register\[3\]\[1\] net553 net533 top.DUT.register\[12\]\[1\] vssd1
+ vssd1 vccd1 vccd1 _03028_ sky130_fd_sc_hd__a22o_1
X_09628_ _01410_ _04657_ _04661_ _04668_ vssd1 vssd1 vccd1 vccd1 _04673_ sky130_fd_sc_hd__a211o_1
XANTENNA__10320__S net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08893__A1 net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07696__A2 net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_194_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_3_7_0_clk_X clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09559_ _04606_ _04607_ vssd1 vssd1 vccd1 vccd1 _04608_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout720_X net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_182_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12570_ clknet_leaf_1_clk _00162_ net916 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[2\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_139_2529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07448__A2 net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_571 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_210 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06656__B1 net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11521_ _05348_ net273 _05346_ vssd1 vssd1 vccd1 vccd1 _05404_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_61_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11452_ _05329_ _05330_ _05334_ vssd1 vssd1 vccd1 vccd1 _05335_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_163_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_799 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_152_2729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10403_ net1584 net244 net369 vssd1 vssd1 vccd1 vccd1 _00575_ sky130_fd_sc_hd__mux2_1
X_11383_ _05260_ _05265_ vssd1 vssd1 vccd1 vccd1 _05266_ sky130_fd_sc_hd__and2_1
XFILLER_0_21_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10334_ net1384 net253 net377 vssd1 vssd1 vccd1 vccd1 _00510_ sky130_fd_sc_hd__mux2_1
X_13122_ clknet_leaf_9_clk _00714_ net948 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[19\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_185_3217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_185_3228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07620__A2 net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13053_ clknet_leaf_127_clk _00645_ net920 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[17\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_76_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_195 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10265_ top.DUT.register\[11\]\[2\] net263 net385 vssd1 vssd1 vccd1 vccd1 _00443_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_76_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12004_ _05873_ _05877_ net126 vssd1 vssd1 vccd1 vccd1 _05887_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_167_2950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10196_ _04959_ net399 vssd1 vssd1 vccd1 vccd1 _04976_ sky130_fd_sc_hd__nand2b_1
XANTENNA__08581__B1 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_204_3501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09514__A1_N net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_204_3512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_205_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout390 net392 vssd1 vssd1 vccd1 vccd1 net390 sky130_fd_sc_hd__buf_6
XFILLER_0_198_460 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12906_ clknet_leaf_120_clk _00498_ net933 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[12\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10230__S net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08884__A1 net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_622 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09847__B1_N _04859_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_185_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06895__B1 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_196_3379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12837_ clknet_leaf_33_clk _00429_ net1042 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[10\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_146_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08636__A1 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_186_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07439__A2 net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08636__B2 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12768_ clknet_leaf_114_clk _00360_ net963 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[8\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_16_208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11640__B1 top.a1.dataIn\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11719_ _05565_ _05595_ vssd1 vssd1 vccd1 vccd1 _05602_ sky130_fd_sc_hd__and2_1
X_12699_ clknet_leaf_124_clk _00291_ net924 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[6\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_154_563 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09046__D1 _03258_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput10 DAT_I[17] vssd1 vssd1 vccd1 vccd1 net10 sky130_fd_sc_hd__buf_1
XFILLER_0_126_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_799 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput21 DAT_I[27] vssd1 vssd1 vccd1 vccd1 net21 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_154_596 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput32 DAT_I[8] vssd1 vssd1 vccd1 vccd1 net32 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_235 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold805 top.DUT.register\[18\]\[31\] vssd1 vssd1 vccd1 vccd1 net1921 sky130_fd_sc_hd__dlygate4sd3_1
Xhold816 top.DUT.register\[23\]\[25\] vssd1 vssd1 vccd1 vccd1 net1932 sky130_fd_sc_hd__dlygate4sd3_1
Xhold827 top.DUT.register\[31\]\[4\] vssd1 vssd1 vccd1 vccd1 net1943 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07072__B1 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold838 top.DUT.register\[8\]\[14\] vssd1 vssd1 vccd1 vccd1 net1954 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold849 top.DUT.register\[29\]\[18\] vssd1 vssd1 vccd1 vccd1 net1965 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_150_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08930_ _04036_ _04037_ vssd1 vssd1 vccd1 vccd1 _04038_ sky130_fd_sc_hd__nand2_1
XFILLER_0_58_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07494__B _02632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10405__S net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08861_ _01788_ _01831_ vssd1 vssd1 vccd1 vccd1 _03972_ sky130_fd_sc_hd__nor2_1
X_07812_ _02949_ _02950_ net411 vssd1 vssd1 vccd1 vccd1 _02951_ sky130_fd_sc_hd__mux2_1
X_08792_ _01921_ _03088_ vssd1 vssd1 vccd1 vccd1 _03907_ sky130_fd_sc_hd__xnor2_1
X_07743_ top.DUT.register\[23\]\[3\] net573 net449 top.DUT.register\[21\]\[3\] _02881_
+ vssd1 vssd1 vccd1 vccd1 _02882_ sky130_fd_sc_hd__a221o_1
XFILLER_0_74_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_770 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout179_A _04868_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10140__S net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07674_ top.DUT.register\[23\]\[4\] net673 net753 top.DUT.register\[26\]\[4\] _02809_
+ vssd1 vssd1 vccd1 vccd1 _02813_ sky130_fd_sc_hd__a221o_1
XANTENNA__08875__A1 _03334_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08875__B2 net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09413_ net821 _02679_ net422 vssd1 vssd1 vccd1 vccd1 _04471_ sky130_fd_sc_hd__a21o_2
XFILLER_0_94_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06625_ _01754_ _01763_ vssd1 vssd1 vccd1 vccd1 _01764_ sky130_fd_sc_hd__nor2_4
XFILLER_0_149_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout346_A _04991_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1088_A net1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_491 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06556_ top.DUT.register\[9\]\[29\] net764 net701 top.DUT.register\[31\]\[29\] _01694_
+ vssd1 vssd1 vccd1 vccd1 _01695_ sky130_fd_sc_hd__a221o_1
XFILLER_0_177_699 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09344_ _04404_ _04405_ vssd1 vssd1 vccd1 vccd1 _04406_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_191_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_205_Left_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06638__B1 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09275_ _04338_ _04340_ _04334_ vssd1 vssd1 vccd1 vccd1 _04341_ sky130_fd_sc_hd__a21oi_1
X_06487_ _01604_ _01625_ vssd1 vssd1 vccd1 vccd1 _01626_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout134_X net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout513_A _01559_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08226_ net280 _03358_ _03362_ net285 vssd1 vssd1 vccd1 vccd1 _03363_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_7_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_43_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07850__A2 net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12187__A1 top.a1.row2\[42\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12364__Q top.a1.dataIn\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_200_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08157_ _03293_ _03294_ vssd1 vssd1 vccd1 vccd1 _03295_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_134_2459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07108_ top.DUT.register\[17\]\[16\] net747 net635 top.DUT.register\[6\]\[16\] vssd1
+ vssd1 vccd1 vccd1 _02247_ sky130_fd_sc_hd__a22o_1
XANTENNA__07063__B1 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08088_ net291 _03226_ vssd1 vssd1 vccd1 vccd1 _03227_ sky130_fd_sc_hd__nor2_1
XANTENNA__07602__A2 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07039_ _02155_ _02176_ vssd1 vssd1 vccd1 vccd1 _02178_ sky130_fd_sc_hd__nand2_1
XANTENNA__10315__S net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_288 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10050_ net1960 net262 net617 vssd1 vssd1 vccd1 vccd1 _00252_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout670_X net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout768_X net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_149_2680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07691__Y _02830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_180_3147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout935_X net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_162_2880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_202_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13740_ clknet_leaf_100_clk _01311_ vssd1 vssd1 vccd1 vccd1 top.lcd.cnt_20ms\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__10050__S net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10952_ top.a1.row1\[101\] _04668_ vssd1 vssd1 vccd1 vccd1 _01113_ sky130_fd_sc_hd__or2_1
XFILLER_0_58_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13671_ clknet_leaf_74_clk _01247_ net1078 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[108\]
+ sky130_fd_sc_hd__dfrtp_1
X_10883_ net161 top.DUT.register\[29\]\[27\] net597 vssd1 vssd1 vccd1 vccd1 _01044_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_155_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12622_ clknet_leaf_39_clk _00214_ net1053 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[3\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_182_102 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09815__B1 net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06629__B1 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_183_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_171_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12553_ clknet_leaf_53_clk _00145_ net1038 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[1\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_136_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_703 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11504_ _05315_ _05345_ vssd1 vssd1 vccd1 vccd1 _05387_ sky130_fd_sc_hd__or2_1
XFILLER_0_108_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_151_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12484_ clknet_leaf_64_clk _00079_ net1092 vssd1 vssd1 vccd1 vccd1 top.ramstore\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07841__A2 net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_550 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11435_ _05306_ _05314_ _05316_ _05317_ vssd1 vssd1 vccd1 vccd1 _05318_ sky130_fd_sc_hd__nor4_1
XFILLER_0_110_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07054__B1 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11366_ _05237_ _05245_ _05248_ vssd1 vssd1 vccd1 vccd1 _05249_ sky130_fd_sc_hd__a21bo_2
XTAP_TAPCELL_ROW_210_3593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10317_ net192 net1764 net383 vssd1 vssd1 vccd1 vccd1 _00494_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13105_ clknet_leaf_112_clk _00697_ net977 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[19\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10225__S net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11297_ top.a1.row1\[60\] _05136_ _05178_ top.a1.row1\[108\] _05184_ vssd1 vssd1
+ vccd1 vccd1 _05186_ sky130_fd_sc_hd__a221o_1
X_13036_ clknet_leaf_61_clk _00628_ net1089 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[16\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_10248_ net204 net2191 net391 vssd1 vssd1 vccd1 vccd1 _00427_ sky130_fd_sc_hd__mux2_1
XANTENNA__08554__B1 net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11845__A top.a1.dataIn\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10179_ _04713_ _04958_ vssd1 vssd1 vccd1 vccd1 _04959_ sky130_fd_sc_hd__nand2_1
XANTENNA__06498__X _01637_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09315__A top.pc\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_198_3419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06580__A2 net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_211 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_105_2016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_202_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06377__C top.a1.instruction\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_8__f_clk_X clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10895__S net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06410_ top.DUT.register\[15\]\[30\] net681 net677 top.DUT.register\[31\]\[30\] vssd1
+ vssd1 vccd1 vccd1 _01549_ sky130_fd_sc_hd__a22o_1
XFILLER_0_186_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_201_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07390_ top.DUT.register\[12\]\[9\] net531 net451 top.DUT.register\[29\]\[9\] _02528_
+ vssd1 vssd1 vccd1 vccd1 _02529_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_33_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06341_ net859 top.ru.next_dready vssd1 vssd1 vccd1 vccd1 _00005_ sky130_fd_sc_hd__or2_1
XFILLER_0_57_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09060_ _03672_ _03697_ _03719_ _03749_ vssd1 vssd1 vccd1 vccd1 _04135_ sky130_fd_sc_hd__or4b_1
XFILLER_0_161_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06272_ top.lcd.cnt_500hz\[1\] top.lcd.cnt_500hz\[0\] top.lcd.cnt_500hz\[2\] vssd1
+ vssd1 vccd1 vccd1 _01435_ sky130_fd_sc_hd__nand3_1
XFILLER_0_142_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07832__A2 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08011_ _03148_ _03149_ vssd1 vssd1 vccd1 vccd1 _03150_ sky130_fd_sc_hd__nor2_1
XFILLER_0_142_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_734 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold602 top.DUT.register\[29\]\[5\] vssd1 vssd1 vccd1 vccd1 net1718 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold613 top.DUT.register\[11\]\[29\] vssd1 vssd1 vccd1 vccd1 net1729 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07045__B1 net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_116_2189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold624 top.DUT.register\[28\]\[23\] vssd1 vssd1 vccd1 vccd1 net1740 sky130_fd_sc_hd__dlygate4sd3_1
Xhold635 top.DUT.register\[11\]\[0\] vssd1 vssd1 vccd1 vccd1 net1751 sky130_fd_sc_hd__dlygate4sd3_1
Xhold646 top.DUT.register\[20\]\[20\] vssd1 vssd1 vccd1 vccd1 net1762 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06399__A2 net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold657 top.DUT.register\[6\]\[24\] vssd1 vssd1 vccd1 vccd1 net1773 sky130_fd_sc_hd__dlygate4sd3_1
Xhold668 top.DUT.register\[22\]\[31\] vssd1 vssd1 vccd1 vccd1 net1784 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10135__S net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09962_ net1480 net215 net628 vssd1 vssd1 vccd1 vccd1 _00170_ sky130_fd_sc_hd__mux2_1
Xhold679 top.DUT.register\[10\]\[1\] vssd1 vssd1 vccd1 vccd1 net1795 sky130_fd_sc_hd__dlygate4sd3_1
X_08913_ _01659_ _03099_ vssd1 vssd1 vccd1 vccd1 _04022_ sky130_fd_sc_hd__xnor2_1
X_09893_ _04897_ _04900_ vssd1 vssd1 vccd1 vccd1 _04902_ sky130_fd_sc_hd__nand2_1
XFILLER_0_40_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout296_A net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08844_ _01764_ net301 _03318_ vssd1 vssd1 vccd1 vccd1 _03956_ sky130_fd_sc_hd__a21boi_1
XANTENNA__12350__S _00016_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07899__A2 net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08775_ net883 top.pc\[23\] net694 _03890_ vssd1 vssd1 vccd1 vccd1 _03891_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout463_A net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06571__A2 net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07016__Y _02155_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07726_ top.DUT.register\[19\]\[3\] net720 net700 top.DUT.register\[31\]\[3\] _02864_
+ vssd1 vssd1 vccd1 vccd1 _02865_ sky130_fd_sc_hd__a221o_1
XANTENNA__08848__A1 net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_192_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06859__B1 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12359__Q top.a1.dataIn\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_177_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout630_A _04948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07657_ _02789_ _02791_ _02793_ _02795_ vssd1 vssd1 vccd1 vccd1 _02796_ sky130_fd_sc_hd__or4_4
XFILLER_0_149_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout349_X net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout728_A _01628_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_154 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06608_ top.DUT.register\[19\]\[27\] net537 net453 top.DUT.register\[29\]\[27\] _01746_
+ vssd1 vssd1 vccd1 vccd1 _01747_ sky130_fd_sc_hd__a221o_1
X_07588_ _02679_ _02725_ net410 vssd1 vssd1 vccd1 vccd1 _02727_ sky130_fd_sc_hd__mux2_1
XFILLER_0_177_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06539_ _01668_ _01677_ vssd1 vssd1 vccd1 vccd1 _01678_ sky130_fd_sc_hd__nor2_4
X_09327_ _04368_ _04371_ vssd1 vssd1 vccd1 vccd1 _04390_ sky130_fd_sc_hd__nand2_1
XFILLER_0_48_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_11_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout516_X net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_180_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09258_ net136 _04312_ _04324_ vssd1 vssd1 vccd1 vccd1 _04325_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07823__A2 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08209_ net313 _03346_ _03321_ vssd1 vssd1 vccd1 vccd1 _03347_ sky130_fd_sc_hd__o21ai_1
X_09189_ _04258_ _04259_ net132 vssd1 vssd1 vccd1 vccd1 _04260_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_177_Right_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_160_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11220_ net845 _05103_ vssd1 vssd1 vccd1 vccd1 _05116_ sky130_fd_sc_hd__and2_1
XFILLER_0_120_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_160_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08304__A net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07587__A1 top.a1.instruction\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout885_X net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11151_ _01429_ _01432_ _05081_ net887 vssd1 vssd1 vccd1 vccd1 _01226_ sky130_fd_sc_hd__o22a_1
XANTENNA__10045__S net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10102_ net1323 net180 net611 vssd1 vssd1 vccd1 vccd1 _00303_ sky130_fd_sc_hd__mux2_1
X_11082_ net905 net1476 net860 _05046_ vssd1 vssd1 vccd1 vccd1 _01192_ sky130_fd_sc_hd__a31o_1
XFILLER_0_101_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10033_ net1361 net187 net621 vssd1 vssd1 vccd1 vccd1 _00236_ sky130_fd_sc_hd__mux2_1
XANTENNA__08000__A2 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09135__A net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input24_A DAT_I[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06478__B _01607_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_160_2839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11984_ _05831_ net127 _05847_ _05849_ vssd1 vssd1 vccd1 vccd1 _05867_ sky130_fd_sc_hd__a22oi_2
X_13723_ clknet_leaf_95_clk _01294_ net986 vssd1 vssd1 vccd1 vccd1 top.a1.row2\[41\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09789__B _04438_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10935_ net1337 net189 net593 vssd1 vssd1 vccd1 vccd1 _01096_ sky130_fd_sc_hd__mux2_1
XFILLER_0_168_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_614 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_193_3338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13654_ clknet_leaf_74_clk _01233_ net1078 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[63\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__08038__X _03177_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10866_ net227 top.DUT.register\[29\]\[10\] net594 vssd1 vssd1 vccd1 vccd1 _01027_
+ sky130_fd_sc_hd__mux2_1
X_12605_ clknet_leaf_119_clk _00197_ net953 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[3\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_66_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_155_146 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13585_ clknet_leaf_46_clk net1203 net1066 vssd1 vssd1 vccd1 vccd1 net76 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_171_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10797_ net254 net1883 net598 vssd1 vssd1 vccd1 vccd1 _00958_ sky130_fd_sc_hd__mux2_1
XFILLER_0_155_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07275__B1 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12536_ clknet_leaf_128_clk _00128_ net912 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[1\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12467_ clknet_leaf_46_clk _00062_ net1066 vssd1 vssd1 vccd1 vccd1 top.ramstore\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07027__B1 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_144_Right_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11418_ _05264_ _05300_ vssd1 vssd1 vccd1 vccd1 _05301_ sky130_fd_sc_hd__nor2_1
XFILLER_0_22_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12398_ clknet_leaf_104_clk top.ru.next_FetchedInstr\[10\] net973 vssd1 vssd1 vccd1
+ vccd1 top.a1.instruction\[10\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_111_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11349_ top.a1.dataIn\[24\] _05214_ _05219_ vssd1 vssd1 vccd1 vccd1 _05232_ sky130_fd_sc_hd__and3_1
XFILLER_0_183_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13019_ clknet_leaf_122_clk _00611_ net928 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[16\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_06890_ top.DUT.register\[9\]\[18\] net763 net744 top.DUT.register\[2\]\[18\] _02028_
+ vssd1 vssd1 vccd1 vccd1 _02029_ sky130_fd_sc_hd__a221o_1
XFILLER_0_206_320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13563__Q top.ramload\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06553__A2 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08560_ _02657_ _03684_ vssd1 vssd1 vccd1 vccd1 _03685_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_89_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07511_ top.DUT.register\[20\]\[14\] net665 net728 top.DUT.register\[18\]\[14\] _02649_
+ vssd1 vssd1 vccd1 vccd1 _02650_ sky130_fd_sc_hd__a221o_1
XFILLER_0_49_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08491_ _02388_ _03596_ _03066_ vssd1 vssd1 vccd1 vccd1 _03619_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_76_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07442_ top.DUT.register\[15\]\[15\] net680 net676 top.DUT.register\[31\]\[15\] vssd1
+ vssd1 vccd1 vccd1 _02581_ sky130_fd_sc_hd__a22o_1
XFILLER_0_147_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07373_ top.DUT.register\[18\]\[8\] net727 net636 top.DUT.register\[6\]\[8\] _02504_
+ vssd1 vssd1 vccd1 vccd1 _02512_ sky130_fd_sc_hd__a221o_1
XFILLER_0_17_314 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_2218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_628 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09112_ _04185_ _04186_ vssd1 vssd1 vccd1 vccd1 _04187_ sky130_fd_sc_hd__nor2_1
X_06324_ _01471_ vssd1 vssd1 vccd1 vccd1 top.edg2.button_i sky130_fd_sc_hd__inv_2
XANTENNA__07266__B1 net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09043_ _02267_ _02659_ _04116_ _04117_ vssd1 vssd1 vccd1 vccd1 _04118_ sky130_fd_sc_hd__or4b_1
X_06255_ net1178 net852 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedData\[16\] sky130_fd_sc_hd__and2_1
XFILLER_0_88_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_2407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_672 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07018__B1 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_2418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_111_Right_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold410 top.DUT.register\[2\]\[1\] vssd1 vssd1 vccd1 vccd1 net1526 sky130_fd_sc_hd__dlygate4sd3_1
X_06186_ net888 _01424_ _01422_ vssd1 vssd1 vccd1 vccd1 top.a1.nextHex\[0\] sky130_fd_sc_hd__mux2_1
Xhold421 top.ramaddr\[6\] vssd1 vssd1 vccd1 vccd1 net1537 sky130_fd_sc_hd__dlygate4sd3_1
Xhold432 top.DUT.register\[7\]\[27\] vssd1 vssd1 vccd1 vccd1 net1548 sky130_fd_sc_hd__dlygate4sd3_1
Xhold443 top.DUT.register\[2\]\[16\] vssd1 vssd1 vccd1 vccd1 net1559 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold454 top.DUT.register\[25\]\[21\] vssd1 vssd1 vccd1 vccd1 net1570 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold465 top.DUT.register\[25\]\[3\] vssd1 vssd1 vccd1 vccd1 net1581 sky130_fd_sc_hd__dlygate4sd3_1
Xhold476 top.DUT.register\[24\]\[21\] vssd1 vssd1 vccd1 vccd1 net1592 sky130_fd_sc_hd__dlygate4sd3_1
Xhold487 top.DUT.register\[1\]\[23\] vssd1 vssd1 vccd1 vccd1 net1603 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout901 net903 vssd1 vssd1 vccd1 vccd1 net901 sky130_fd_sc_hd__buf_2
Xhold498 top.DUT.register\[13\]\[13\] vssd1 vssd1 vccd1 vccd1 net1614 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout912 net913 vssd1 vssd1 vccd1 vccd1 net912 sky130_fd_sc_hd__clkbuf_4
X_09945_ net2059 net145 net627 vssd1 vssd1 vccd1 vccd1 _00153_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout923 net925 vssd1 vssd1 vccd1 vccd1 net923 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout580_A _01514_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_147_Left_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout934 net935 vssd1 vssd1 vccd1 vccd1 net934 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08518__B1 _03643_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout678_A _01548_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout945 net952 vssd1 vssd1 vccd1 vccd1 net945 sky130_fd_sc_hd__clkbuf_2
XANTENNA__06792__A2 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout956 net966 vssd1 vssd1 vccd1 vccd1 net956 sky130_fd_sc_hd__buf_2
Xfanout967 net1098 vssd1 vssd1 vccd1 vccd1 net967 sky130_fd_sc_hd__clkbuf_4
X_09876_ _03950_ _04716_ vssd1 vssd1 vccd1 vccd1 _04886_ sky130_fd_sc_hd__nand2_1
Xfanout978 net979 vssd1 vssd1 vccd1 vccd1 net978 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout1006_X net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1110 top.DUT.register\[18\]\[24\] vssd1 vssd1 vccd1 vccd1 net2226 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout989 net990 vssd1 vssd1 vccd1 vccd1 net989 sky130_fd_sc_hd__clkbuf_4
Xhold1121 top.DUT.register\[6\]\[3\] vssd1 vssd1 vccd1 vccd1 net2237 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1132 top.DUT.register\[6\]\[27\] vssd1 vssd1 vccd1 vccd1 net2248 sky130_fd_sc_hd__dlygate4sd3_1
X_08827_ net325 _03605_ _03939_ net285 vssd1 vssd1 vccd1 vccd1 _03940_ sky130_fd_sc_hd__a2bb2o_1
Xhold1143 top.pad.keyCode\[6\] vssd1 vssd1 vccd1 vccd1 net2259 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1154 top.DUT.register\[4\]\[26\] vssd1 vssd1 vccd1 vccd1 net2270 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout466_X net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06544__A2 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1165 top.DUT.register\[14\]\[0\] vssd1 vssd1 vccd1 vccd1 net2281 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07741__A1 _02878_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1176 top.DUT.register\[9\]\[29\] vssd1 vssd1 vccd1 vccd1 net2292 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1187 top.DUT.register\[12\]\[30\] vssd1 vssd1 vccd1 vccd1 net2303 sky130_fd_sc_hd__dlygate4sd3_1
X_08758_ _03301_ _03304_ vssd1 vssd1 vccd1 vccd1 _03874_ sky130_fd_sc_hd__nand2_1
Xhold1198 top.ramload\[19\] vssd1 vssd1 vccd1 vccd1 net2314 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_197_547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_142_2569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07709_ _02841_ _02843_ _02845_ _02847_ vssd1 vssd1 vccd1 vccd1 _02848_ sky130_fd_sc_hd__or4_2
XFILLER_0_178_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08689_ net1294 net830 net800 _03808_ vssd1 vssd1 vccd1 vccd1 _00037_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout633_X net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10720_ net1999 net172 net335 vssd1 vssd1 vccd1 vccd1 _00881_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_156_Left_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_175_3068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08049__A2 net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10651_ net180 net2003 net343 vssd1 vssd1 vccd1 vccd1 _00815_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_180_403 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07257__B1 net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10582_ net1659 net186 net352 vssd1 vssd1 vccd1 vccd1 _00748_ sky130_fd_sc_hd__mux2_1
X_13370_ clknet_leaf_1_clk _00962_ net917 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[27\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_146_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_306 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12321_ top.pad.button_control.r_counter\[7\] _06122_ _06124_ net790 vssd1 vssd1
+ vccd1 vccd1 _01359_ sky130_fd_sc_hd__o211a_1
XANTENNA__07857__B _02994_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_339 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08305__Y _03440_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07009__B1 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12252_ net1195 _06080_ _06082_ vssd1 vssd1 vccd1 vccd1 _01326_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_170_2990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11203_ net845 _05015_ _05027_ vssd1 vssd1 vccd1 vccd1 _05108_ sky130_fd_sc_hd__and3_1
X_12183_ top.a1.row2\[34\] net847 net797 _05819_ vssd1 vssd1 vccd1 vccd1 _01291_ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_61_clk_A clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_165_Left_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_71_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11134_ net907 net1923 net862 _05072_ vssd1 vssd1 vccd1 vccd1 _01218_ sky130_fd_sc_hd__a31o_1
XANTENNA__06783__A2 net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11065_ net80 net870 net834 net1205 vssd1 vssd1 vccd1 vccd1 _01176_ sky130_fd_sc_hd__a22o_1
XANTENNA__10503__S net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10016_ top.DUT.register\[4\]\[2\] net264 net619 vssd1 vssd1 vccd1 vccd1 _00219_
+ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_76_clk_A clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_204_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06535__A2 net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09612__A_N top.a1.halfData\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07812__S net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_174_Left_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11967_ _05849_ vssd1 vssd1 vccd1 vccd1 _05850_ sky130_fd_sc_hd__inv_2
XFILLER_0_98_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_169_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13706_ clknet_leaf_96_clk _01277_ net985 vssd1 vssd1 vccd1 vccd1 top.a1.row2\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_196_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07496__B1 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10918_ net1438 net148 net480 vssd1 vssd1 vccd1 vccd1 _01079_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11898_ _05710_ _05780_ vssd1 vssd1 vccd1 vccd1 _05781_ sky130_fd_sc_hd__xor2_2
X_13637_ clknet_leaf_95_clk net887 net987 vssd1 vssd1 vccd1 vccd1 wb.prev_BUSY_O sky130_fd_sc_hd__dfrtp_1
X_10849_ net1864 net170 net474 vssd1 vssd1 vccd1 vccd1 _01010_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_14_clk_A clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06952__A _02069_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_436 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13568_ clknet_leaf_105_clk _01155_ net972 vssd1 vssd1 vccd1 vccd1 top.ramload\[29\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_15_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13781__RESET_B net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12519_ clknet_leaf_77_clk _00111_ net1083 vssd1 vssd1 vccd1 vccd1 top.pc\[31\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_124_352 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13499_ clknet_leaf_124_clk _01091_ net925 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[31\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11289__B _05120_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_183_Left_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10193__B net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_2137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_113_2148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_558 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_29_clk_A clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07420__B1 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout208 net210 vssd1 vssd1 vccd1 vccd1 net208 sky130_fd_sc_hd__clkbuf_2
Xfanout219 net220 vssd1 vssd1 vccd1 vccd1 net219 sky130_fd_sc_hd__clkbuf_2
X_07991_ top.DUT.register\[12\]\[31\] net741 net704 top.DUT.register\[3\]\[31\] vssd1
+ vssd1 vccd1 vccd1 _03130_ sky130_fd_sc_hd__a22o_1
XANTENNA__06774__A2 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09730_ net2001 net235 net632 vssd1 vssd1 vccd1 vccd1 _00129_ sky130_fd_sc_hd__mux2_1
X_06942_ top.DUT.register\[7\]\[21\] net661 net764 top.DUT.register\[9\]\[21\] vssd1
+ vssd1 vccd1 vccd1 _02081_ sky130_fd_sc_hd__a22o_1
XANTENNA__10413__S net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_207_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09661_ _04674_ _04689_ _04677_ vssd1 vssd1 vccd1 vccd1 _04700_ sky130_fd_sc_hd__a21oi_1
X_06873_ top.DUT.register\[9\]\[18\] net468 net569 top.DUT.register\[6\]\[18\] vssd1
+ vssd1 vccd1 vccd1 _02012_ sky130_fd_sc_hd__a22o_1
XANTENNA__06526__A2 net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08612_ net279 _03554_ _03734_ net283 vssd1 vssd1 vccd1 vccd1 _03735_ sky130_fd_sc_hd__o22a_1
X_09592_ _04637_ _04638_ vssd1 vssd1 vccd1 vccd1 _04639_ sky130_fd_sc_hd__nand2_1
XFILLER_0_82_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08543_ net496 _03668_ vssd1 vssd1 vccd1 vccd1 _03669_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout161_A _04906_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_534 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_124_2299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout259_A net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07487__B1 net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08474_ net309 _03503_ _03602_ vssd1 vssd1 vccd1 vccd1 _03603_ sky130_fd_sc_hd__o21ai_1
XANTENNA__11283__B2 top.a1.row2\[43\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_175_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07425_ top.DUT.register\[4\]\[9\] net667 net635 top.DUT.register\[6\]\[9\] _02563_
+ vssd1 vssd1 vccd1 vccd1 _02564_ sky130_fd_sc_hd__a221o_1
XFILLER_0_190_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1070_A net1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout426_A net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07239__B1 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11035__B2 top.ramload\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07356_ top.DUT.register\[9\]\[8\] net467 net540 top.DUT.register\[8\]\[8\] _02494_
+ vssd1 vssd1 vccd1 vccd1 _02495_ sky130_fd_sc_hd__a221o_1
XFILLER_0_18_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_21_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_190_778 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06307_ _01451_ _01453_ vssd1 vssd1 vccd1 vccd1 _01463_ sky130_fd_sc_hd__nor2_1
X_07287_ top.DUT.register\[5\]\[13\] net653 net744 top.DUT.register\[2\]\[13\] _02410_
+ vssd1 vssd1 vccd1 vccd1 _02426_ sky130_fd_sc_hd__a221o_1
XFILLER_0_33_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_659 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09026_ _02134_ _02307_ _03177_ _03185_ vssd1 vssd1 vccd1 vccd1 _04101_ sky130_fd_sc_hd__or4_1
X_06238_ top.busy_o top.ru.state\[4\] vssd1 vssd1 vccd1 vccd1 _01433_ sky130_fd_sc_hd__and2b_1
XFILLER_0_20_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12372__Q top.a1.dataIn\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout795_A _01489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold240 top.DUT.register\[20\]\[30\] vssd1 vssd1 vccd1 vccd1 net1356 sky130_fd_sc_hd__dlygate4sd3_1
X_06169_ top.a1.halfData\[2\] top.a1.halfData\[1\] vssd1 vssd1 vccd1 vccd1 _01411_
+ sky130_fd_sc_hd__and2b_1
Xhold251 top.DUT.register\[24\]\[20\] vssd1 vssd1 vccd1 vccd1 net1367 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09400__A1 net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold262 top.a1.row2\[11\] vssd1 vssd1 vccd1 vccd1 net1378 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09400__B2 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold273 top.DUT.register\[1\]\[1\] vssd1 vssd1 vccd1 vccd1 net1389 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07411__B1 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold284 top.DUT.register\[12\]\[15\] vssd1 vssd1 vccd1 vccd1 net1400 sky130_fd_sc_hd__dlygate4sd3_1
Xhold295 top.DUT.register\[15\]\[31\] vssd1 vssd1 vccd1 vccd1 net1411 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout583_X net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout962_A net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06765__A2 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout720 _01635_ vssd1 vssd1 vccd1 vccd1 net720 sky130_fd_sc_hd__clkbuf_8
Xfanout731 _01627_ vssd1 vssd1 vccd1 vccd1 net731 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10323__S net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout742 _01623_ vssd1 vssd1 vccd1 vccd1 net742 sky130_fd_sc_hd__clkbuf_8
X_09928_ _04930_ _04933_ vssd1 vssd1 vccd1 vccd1 _04934_ sky130_fd_sc_hd__xor2_1
Xfanout753 _01621_ vssd1 vssd1 vccd1 vccd1 net753 sky130_fd_sc_hd__buf_4
Xfanout764 net765 vssd1 vssd1 vccd1 vccd1 net764 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_144_2609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout775 net777 vssd1 vssd1 vccd1 vccd1 net775 sky130_fd_sc_hd__clkbuf_8
Xfanout786 _04708_ vssd1 vssd1 vccd1 vccd1 net786 sky130_fd_sc_hd__buf_2
XANTENNA__09703__A2 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout750_X net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout797 _05082_ vssd1 vssd1 vccd1 vccd1 net797 sky130_fd_sc_hd__clkbuf_4
X_09859_ _04870_ _04869_ vssd1 vssd1 vccd1 vccd1 _04871_ sky130_fd_sc_hd__and2b_1
XFILLER_0_99_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06517__A2 _01655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout848_X net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12870_ clknet_leaf_38_clk _00462_ net1054 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[11\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_177_3108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11821_ _05693_ _05694_ _05691_ _05692_ vssd1 vssd1 vccd1 vccd1 _05704_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_1_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07478__B1 net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11752_ _05572_ _05634_ vssd1 vssd1 vccd1 vccd1 _05635_ sky130_fd_sc_hd__nor2_1
XANTENNA__11274__B2 top.a1.row2\[42\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_159_2830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09700__X _04733_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10703_ net1415 net247 net334 vssd1 vssd1 vccd1 vccd1 _00864_ sky130_fd_sc_hd__mux2_1
XFILLER_0_193_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11683_ _05562_ _05565_ _05561_ vssd1 vssd1 vccd1 vccd1 _05566_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_81_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_548 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13422_ clknet_leaf_40_clk _01014_ net1047 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[28\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_10634_ net251 net2107 net342 vssd1 vssd1 vccd1 vccd1 _00798_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_767 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13353_ clknet_leaf_52_clk _00945_ net1034 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[26\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10565_ top.DUT.register\[20\]\[2\] net263 net350 vssd1 vssd1 vccd1 vccd1 _00731_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12304_ top.pad.button_control.r_counter\[0\] net1265 _06113_ vssd1 vssd1 vccd1 vccd1
+ _01353_ sky130_fd_sc_hd__a21oi_1
X_13284_ clknet_leaf_40_clk _00876_ net1050 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[24\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_161_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10496_ net1365 net145 net357 vssd1 vssd1 vccd1 vccd1 _00665_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_188_3259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12235_ top.lcd.cnt_20ms\[9\] _06070_ net978 vssd1 vssd1 vccd1 vccd1 _06072_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07402__B1 net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12166_ _06035_ _06037_ _06040_ vssd1 vssd1 vccd1 vccd1 _06047_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_208_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07953__A1 _01854_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06756__A2 net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11117_ net49 net867 vssd1 vssd1 vccd1 vccd1 _05064_ sky130_fd_sc_hd__and2_1
XANTENNA__09307__B _02408_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10233__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12097_ _05971_ _05979_ vssd1 vssd1 vccd1 vccd1 _05980_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_207_3554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11048_ net72 net860 _01429_ vssd1 vssd1 vccd1 vccd1 _01159_ sky130_fd_sc_hd__o21a_1
XANTENNA__09026__C _03177_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput8 DAT_I[15] vssd1 vssd1 vccd1 vccd1 net8 sky130_fd_sc_hd__clkbuf_1
XANTENNA__06508__A2 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_311 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07181__A2 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12999_ clknet_leaf_12_clk _00591_ net938 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[15\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_203_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11265__A1 top.a1.row1\[57\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_146_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08130__A1 net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09977__B _04708_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08681__A2 net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07210_ _02342_ _02347_ _02348_ vssd1 vssd1 vccd1 vccd1 _02349_ sky130_fd_sc_hd__or3b_1
X_08190_ net313 _03327_ _03321_ vssd1 vssd1 vccd1 vccd1 _03328_ sky130_fd_sc_hd__o21a_1
XANTENNA__12214__B1 net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08226__X _03363_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_1932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07141_ top.DUT.register\[5\]\[11\] net439 net503 top.DUT.register\[27\]\[11\] _02279_
+ vssd1 vssd1 vccd1 vccd1 _02280_ sky130_fd_sc_hd__a221o_1
XFILLER_0_6_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_171_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_191_Left_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10408__S net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08433__A2 _03561_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07641__B1 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07072_ top.DUT.register\[13\]\[22\] net777 net715 top.DUT.register\[27\]\[22\] vssd1
+ vssd1 vccd1 vccd1 _02211_ sky130_fd_sc_hd__a22o_1
XFILLER_0_112_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_140_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08402__A net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06747__A2 net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12844__RESET_B net1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10143__S net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07974_ top.DUT.register\[25\]\[31\] net458 _03112_ vssd1 vssd1 vccd1 vccd1 _03113_
+ sky130_fd_sc_hd__a21o_1
X_09713_ top.a1.dataIn\[6\] net795 net799 top.pc\[6\] _04742_ vssd1 vssd1 vccd1 vccd1
+ _04743_ sky130_fd_sc_hd__a221o_1
X_06925_ top.DUT.register\[23\]\[21\] net574 net450 top.DUT.register\[21\]\[21\] vssd1
+ vssd1 vccd1 vccd1 _02064_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_126_2339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout376_A _04981_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_311 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09644_ _04677_ _04680_ _04685_ vssd1 vssd1 vccd1 vccd1 _04686_ sky130_fd_sc_hd__o21bai_1
X_06856_ top.DUT.register\[24\]\[19\] net645 net721 top.DUT.register\[19\]\[19\] _01994_
+ vssd1 vssd1 vccd1 vccd1 _01995_ sky130_fd_sc_hd__a221o_1
XANTENNA__13111__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07172__A2 net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09575_ _04606_ _04621_ vssd1 vssd1 vccd1 vccd1 _04623_ sky130_fd_sc_hd__nor2_1
XANTENNA__09449__A1 net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout543_A net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06787_ top.DUT.register\[2\]\[17\] net560 net547 top.DUT.register\[18\]\[17\] vssd1
+ vssd1 vccd1 vccd1 _01926_ sky130_fd_sc_hd__a22o_1
XFILLER_0_179_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_26_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08526_ net324 _03652_ vssd1 vssd1 vccd1 vccd1 _03653_ sky130_fd_sc_hd__nand2_1
XANTENNA__12367__Q top.a1.dataIn\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_203_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08457_ net317 net333 vssd1 vssd1 vccd1 vccd1 _03587_ sky130_fd_sc_hd__nand2_2
XANTENNA_fanout710_A _01638_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09887__B net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_172_3027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout808_A net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout429_X net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1073_X net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_175_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07408_ top.a1.instruction\[30\] net806 _02546_ vssd1 vssd1 vccd1 vccd1 _02547_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11008__B2 top.a1.dataIn\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xwire417 _01872_ vssd1 vssd1 vccd1 vccd1 net417 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_135_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08388_ _03055_ _03519_ vssd1 vssd1 vccd1 vccd1 _03520_ sky130_fd_sc_hd__xor2_1
XFILLER_0_92_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07339_ _02434_ _02476_ vssd1 vssd1 vccd1 vccd1 _02478_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_154_2760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10318__S net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10350_ net1720 net192 net378 vssd1 vssd1 vccd1 vccd1 _00526_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07632__B1 net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout798_X net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06986__A2 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09009_ net425 _03376_ _03414_ vssd1 vssd1 vccd1 vccd1 _04084_ sky130_fd_sc_hd__and3_1
X_10281_ net1630 net205 net387 vssd1 vssd1 vccd1 vccd1 _00459_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_3_3_0_clk_X clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12020_ _05902_ _05878_ _05857_ vssd1 vssd1 vccd1 vccd1 _05903_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout965_X net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10053__S net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08031__B net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_183_3189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout550 _01536_ vssd1 vssd1 vccd1 vccd1 net550 sky130_fd_sc_hd__clkbuf_8
Xfanout561 _01532_ vssd1 vssd1 vccd1 vccd1 net561 sky130_fd_sc_hd__clkbuf_8
Xfanout572 _01519_ vssd1 vssd1 vccd1 vccd1 net572 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12514__RESET_B net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout583 _01513_ vssd1 vssd1 vccd1 vccd1 net583 sky130_fd_sc_hd__clkbuf_8
XANTENNA__09688__A1 _03265_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout594 _04966_ vssd1 vssd1 vccd1 vccd1 net594 sky130_fd_sc_hd__clkbuf_8
X_12922_ clknet_leaf_5_clk _00514_ net936 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[13\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07699__B1 net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07163__A2 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12853_ clknet_leaf_31_clk _00445_ net1023 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[11\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_202_3473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_185_314 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11804_ _05654_ _05656_ _05680_ _05646_ vssd1 vssd1 vccd1 vccd1 _05687_ sky130_fd_sc_hd__a2bb2o_2
X_12784_ clknet_leaf_31_clk _00376_ net1018 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[8\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_11735_ _05609_ _05615_ vssd1 vssd1 vccd1 vccd1 _05618_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_113_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11666_ _05542_ _05548_ _05520_ vssd1 vssd1 vccd1 vccd1 _05549_ sky130_fd_sc_hd__a21o_2
XANTENNA__07871__B1 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08046__X _03185_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13405_ clknet_leaf_13_clk _00997_ net941 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[28\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_10617_ net194 net1638 net348 vssd1 vssd1 vccd1 vccd1 _00782_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10228__S net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11597_ _05443_ _05478_ vssd1 vssd1 vccd1 vccd1 _05480_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_141_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13336_ clknet_leaf_125_clk _00928_ net923 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[26\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07623__B1 net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10548_ net2260 net203 net356 vssd1 vssd1 vccd1 vccd1 _00715_ sky130_fd_sc_hd__mux2_1
Xclkbuf_4_5__f_clk clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_5__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_51_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06977__A2 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13267_ clknet_leaf_122_clk _00859_ net932 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[24\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_94_1851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10479_ net2128 net224 net362 vssd1 vssd1 vccd1 vccd1 _00649_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_94_1862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09759__A1_N net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12218_ _06051_ _06061_ vssd1 vssd1 vccd1 vccd1 _06062_ sky130_fd_sc_hd__nor2_1
XANTENNA__09318__A top.pc\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13198_ clknet_leaf_41_clk _00790_ net1045 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[21\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11183__B1 net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06729__A2 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12149_ _06014_ _06020_ _06025_ _06031_ vssd1 vssd1 vccd1 vccd1 _06032_ sky130_fd_sc_hd__o31ai_1
XANTENNA_max_cap606_A _04957_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10898__S net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06710_ top.DUT.register\[14\]\[25\] net583 net551 top.DUT.register\[3\]\[25\] _01848_
+ vssd1 vssd1 vccd1 vccd1 _01849_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_108_2069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07690_ net824 _02808_ _02828_ vssd1 vssd1 vccd1 vccd1 _02829_ sky130_fd_sc_hd__o21a_1
XANTENNA__08351__A1 net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07154__A2 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09053__A _03560_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_204_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_188_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06641_ top.DUT.register\[25\]\[27\] net781 _01779_ vssd1 vssd1 vccd1 vccd1 _01780_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_78_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13284__CLK clknet_leaf_40_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06901__A2 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09360_ _02232_ _02241_ _04420_ vssd1 vssd1 vccd1 vccd1 _04421_ sky130_fd_sc_hd__o21ai_1
X_06572_ _01704_ _01706_ _01708_ _01710_ vssd1 vssd1 vccd1 vccd1 _01711_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_121_2258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08311_ _02852_ _03445_ vssd1 vssd1 vccd1 vccd1 _03446_ sky130_fd_sc_hd__xor2_1
XFILLER_0_19_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09291_ _04334_ _04339_ _04338_ vssd1 vssd1 vccd1 vccd1 _04356_ sky130_fd_sc_hd__o21a_1
XFILLER_0_170_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08953__A1_N _02566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08242_ _03378_ vssd1 vssd1 vccd1 vccd1 _03379_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_103_1991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07862__B1 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_678 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08173_ _02026_ net327 vssd1 vssd1 vccd1 vccd1 _03311_ sky130_fd_sc_hd__nand2_1
XFILLER_0_27_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10138__S net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_172_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07795__X _02934_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07124_ _02242_ _02261_ vssd1 vssd1 vccd1 vccd1 _02263_ sky130_fd_sc_hd__nor2_1
XFILLER_0_125_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08968__A1_N _01916_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_2490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06968__A2 net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07055_ top.DUT.register\[25\]\[22\] net455 net451 top.DUT.register\[29\]\[22\] _02193_
+ vssd1 vssd1 vccd1 vccd1 _02194_ sky130_fd_sc_hd__a221o_1
XFILLER_0_88_62 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput120 net120 vssd1 vssd1 vccd1 vccd1 gpio_out[22] sky130_fd_sc_hd__buf_2
XFILLER_0_112_152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08132__A _02590_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout493_A _03339_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07917__A1 _02678_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_695 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_hold1141_A top.ramload\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07393__A2 net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07957_ _01785_ _03095_ _01745_ vssd1 vssd1 vccd1 vccd1 _03096_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout660_A net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout758_A _01617_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout379_X net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06908_ _02026_ _02046_ vssd1 vssd1 vccd1 vccd1 _02047_ sky130_fd_sc_hd__nor2_2
XANTENNA__10601__S net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07888_ top.DUT.register\[18\]\[1\] net548 net528 top.DUT.register\[26\]\[1\] _03026_
+ vssd1 vssd1 vccd1 vccd1 _03027_ sky130_fd_sc_hd__a221o_1
XANTENNA__07145__A2 net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09627_ _04164_ _04660_ _04665_ _04658_ _04670_ vssd1 vssd1 vccd1 vccd1 _04672_ sky130_fd_sc_hd__o221a_1
X_06839_ top.DUT.register\[23\]\[19\] net574 net534 top.DUT.register\[12\]\[19\] vssd1
+ vssd1 vccd1 vccd1 _01978_ sky130_fd_sc_hd__a22o_1
XFILLER_0_195_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout546_X net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout925_A net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09558_ _01722_ _04605_ vssd1 vssd1 vccd1 vccd1 _04607_ sky130_fd_sc_hd__or2_1
XFILLER_0_65_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12651__CLK clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08509_ _02310_ _03636_ vssd1 vssd1 vccd1 vccd1 _03637_ sky130_fd_sc_hd__xnor2_1
XANTENNA__08645__A2 net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09842__A1 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09489_ net134 _04541_ vssd1 vssd1 vccd1 vccd1 _04542_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout713_X net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_194_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_194_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11520_ _05396_ _05398_ _05374_ _05376_ _05378_ vssd1 vssd1 vccd1 vccd1 _05403_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_53_507 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07853__B1 net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_175_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11451_ _05332_ _05333_ _05296_ _05325_ vssd1 vssd1 vccd1 vccd1 _05334_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_152_2719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10048__S net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10402_ net1510 net251 net369 vssd1 vssd1 vccd1 vccd1 _00574_ sky130_fd_sc_hd__mux2_1
XANTENNA__07605__B1 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11382_ _05263_ _05264_ vssd1 vssd1 vccd1 vccd1 _05265_ sky130_fd_sc_hd__nor2_1
XFILLER_0_61_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06959__A2 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13121_ clknet_leaf_15_clk _00713_ net962 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[19\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10333_ net1734 net257 net378 vssd1 vssd1 vccd1 vccd1 _00509_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_185_3218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13052_ clknet_leaf_130_clk _00644_ net914 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[17\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_76_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10264_ net2224 net270 net388 vssd1 vssd1 vccd1 vccd1 _00442_ sky130_fd_sc_hd__mux2_1
XANTENNA__08042__A _03152_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12003_ _05883_ _05885_ vssd1 vssd1 vccd1 vccd1 _05886_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_167_2951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10195_ net418 _04974_ net598 _04970_ vssd1 vssd1 vccd1 vccd1 _04975_ sky130_fd_sc_hd__and4bb_1
XANTENNA__08581__A1 net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11180__A3 net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08581__B2 _03705_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_204_3502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_204_3513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06592__B1 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout380 _04980_ vssd1 vssd1 vccd1 vccd1 net380 sky130_fd_sc_hd__buf_4
Xclkbuf_4_13__f_clk clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_13__leaf_clk
+ sky130_fd_sc_hd__clkbuf_16
Xfanout391 net392 vssd1 vssd1 vccd1 vccd1 net391 sky130_fd_sc_hd__buf_4
XFILLER_0_108_49 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10511__S net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_205_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07136__A2 net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12905_ clknet_leaf_52_clk _00497_ net1035 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[12\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_198_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_201_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12836_ clknet_leaf_36_clk _00428_ net1049 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[10\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_186_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_174_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09294__C1 net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12767_ clknet_leaf_20_clk _00359_ net1028 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[8\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_139_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09833__A1 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11718_ _05596_ _05600_ vssd1 vssd1 vccd1 vccd1 _05601_ sky130_fd_sc_hd__or2_1
XANTENNA__07844__B1 net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12698_ clknet_leaf_1_clk _00290_ net917 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[6\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09046__C1 _04041_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11649_ _05501_ _05503_ _05506_ vssd1 vssd1 vccd1 vccd1 _05532_ sky130_fd_sc_hd__and3_1
Xinput11 DAT_I[18] vssd1 vssd1 vccd1 vccd1 net11 sky130_fd_sc_hd__buf_1
Xinput22 DAT_I[28] vssd1 vssd1 vccd1 vccd1 net22 sky130_fd_sc_hd__clkbuf_1
XANTENNA__10185__C net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput33 DAT_I[9] vssd1 vssd1 vccd1 vccd1 net33 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold806 top.DUT.register\[17\]\[14\] vssd1 vssd1 vccd1 vccd1 net1922 sky130_fd_sc_hd__dlygate4sd3_1
Xhold817 top.DUT.register\[12\]\[5\] vssd1 vssd1 vccd1 vccd1 net1933 sky130_fd_sc_hd__dlygate4sd3_1
Xhold828 top.DUT.register\[31\]\[29\] vssd1 vssd1 vccd1 vccd1 net1944 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13319_ clknet_leaf_4_clk _00911_ net938 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[25\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold839 top.DUT.register\[12\]\[2\] vssd1 vssd1 vccd1 vccd1 net1955 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13566__Q top.ramload\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_656 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12470__Q top.ramstore\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08860_ net1317 net831 net801 _03971_ vssd1 vssd1 vccd1 vccd1 _00045_ sky130_fd_sc_hd__a22o_1
XANTENNA__08887__A net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07375__A2 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07811_ net820 _02363_ vssd1 vssd1 vccd1 vccd1 _02950_ sky130_fd_sc_hd__and2_1
X_08791_ _03258_ _03260_ _03905_ vssd1 vssd1 vccd1 vccd1 _03906_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_165_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10421__S net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07742_ top.DUT.register\[12\]\[3\] net533 net458 top.DUT.register\[25\]\[3\] vssd1
+ vssd1 vccd1 vccd1 _02881_ sky130_fd_sc_hd__a22o_1
XFILLER_0_74_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08324__A1 net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08324__B2 _03263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_205_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07673_ top.DUT.register\[2\]\[4\] net744 net724 top.DUT.register\[29\]\[4\] vssd1
+ vssd1 vccd1 vccd1 _02812_ sky130_fd_sc_hd__a22o_1
X_09412_ net821 _01585_ vssd1 vssd1 vccd1 vccd1 _04470_ sky130_fd_sc_hd__nor2_1
X_06624_ _01758_ _01760_ _01762_ vssd1 vssd1 vccd1 vccd1 _01763_ sky130_fd_sc_hd__or3_4
XFILLER_0_137_509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09343_ _02580_ _02589_ _04403_ vssd1 vssd1 vccd1 vccd1 _04405_ sky130_fd_sc_hd__or3_1
X_06555_ top.DUT.register\[24\]\[29\] net645 net704 top.DUT.register\[3\]\[29\] _01693_
+ vssd1 vssd1 vccd1 vccd1 _01694_ sky130_fd_sc_hd__a221o_1
XANTENNA__12348__S _00016_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09824__A1 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_158_Right_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout339_A _04993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_16_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09274_ _02286_ _04337_ vssd1 vssd1 vccd1 vccd1 _04340_ sky130_fd_sc_hd__or2_1
X_06486_ top.a1.instruction\[22\] top.a1.instruction\[23\] net792 vssd1 vssd1 vccd1
+ vccd1 _01625_ sky130_fd_sc_hd__o21a_1
XFILLER_0_191_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08225_ net304 _03359_ _03360_ _03361_ vssd1 vssd1 vccd1 vccd1 _03362_ sky130_fd_sc_hd__a22o_1
XFILLER_0_133_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout506_A _01567_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12187__A2 net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08156_ _02723_ net331 vssd1 vssd1 vccd1 vccd1 _03294_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_134_2449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07107_ top.DUT.register\[7\]\[16\] net660 net763 top.DUT.register\[9\]\[16\] _02245_
+ vssd1 vssd1 vccd1 vccd1 _02246_ sky130_fd_sc_hd__a221o_1
XFILLER_0_132_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_160_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08087_ _03224_ _03225_ vssd1 vssd1 vccd1 vccd1 _03226_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07038_ _02155_ _02176_ vssd1 vssd1 vccd1 vccd1 _02177_ sky130_fd_sc_hd__nor2_1
XFILLER_0_140_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout496_X net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07366__A2 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input1_X net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_149_2681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_180_3148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08989_ _01699_ _01743_ vssd1 vssd1 vccd1 vccd1 _04064_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout663_X net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10331__S net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07118__A2 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_162_2870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_162_2881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10951_ net1892 net143 net591 vssd1 vssd1 vccd1 vccd1 _01112_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout928_X net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13670_ clknet_leaf_91_clk _01246_ net996 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[123\]
+ sky130_fd_sc_hd__dfrtp_1
X_10882_ net164 top.DUT.register\[29\]\[26\] net597 vssd1 vssd1 vccd1 vccd1 _01043_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_168_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_211_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12621_ clknet_leaf_45_clk _00213_ net1064 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[3\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_183_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08618__A2 _03185_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09815__A1 _03807_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_182_114 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_125_Right_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_14_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07826__B1 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12552_ clknet_leaf_7_clk _00144_ net946 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[1\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_182_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08037__A net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11503_ _05384_ _05385_ _05352_ vssd1 vssd1 vccd1 vccd1 _05386_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_124_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12483_ clknet_leaf_65_clk _00078_ net1094 vssd1 vssd1 vccd1 vccd1 top.ramstore\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12178__A2 net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11434_ _05263_ _05301_ vssd1 vssd1 vccd1 vccd1 _05317_ sky130_fd_sc_hd__xnor2_2
XTAP_TAPCELL_ROW_78_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06780__A _01897_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_100_clk clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_100_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__10506__S net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11365_ top.a1.dataIn\[30\] _05218_ _05247_ vssd1 vssd1 vccd1 vccd1 _05248_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_91_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13104_ clknet_leaf_29_clk _00696_ net1017 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[18\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_10316_ net201 net1889 net382 vssd1 vssd1 vccd1 vccd1 _00493_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_210_3594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11296_ net878 net881 top.a1.row2\[12\] _05118_ vssd1 vssd1 vccd1 vccd1 _05185_ sky130_fd_sc_hd__o211a_1
X_13035_ clknet_leaf_50_clk _00627_ net1059 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[16\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08003__B1 net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10247_ net216 net1613 net389 vssd1 vssd1 vccd1 vccd1 _00426_ sky130_fd_sc_hd__mux2_1
XANTENNA__08554__B2 _03673_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06565__B1 net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10178_ top.a1.instruction\[9\] _04711_ vssd1 vssd1 vccd1 vccd1 _04958_ sky130_fd_sc_hd__nor2_1
XFILLER_0_28_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_198_3409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10241__S net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08306__A1 net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07109__A2 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_2017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_223 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11310__B1 _05123_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_198_280 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_159_656 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12819_ clknet_leaf_124_clk _00411_ net928 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[10\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_13799_ clknet_leaf_68_clk _01368_ vssd1 vssd1 vccd1 vccd1 top.pad.button_control.r_counter\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_33_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_146_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06340_ top.lcd.cnt_500hz\[13\] _01483_ top.lcd.cnt_500hz\[14\] vssd1 vssd1 vccd1
+ vccd1 top.lcd.lcd_en sky130_fd_sc_hd__a21oi_1
XFILLER_0_139_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_1950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06271_ top.lcd.cnt_500hz\[1\] top.lcd.cnt_500hz\[0\] vssd1 vssd1 vccd1 vccd1 _01434_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_56_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08010_ _01391_ top.a1.instruction\[13\] net893 vssd1 vssd1 vccd1 vccd1 _03149_ sky130_fd_sc_hd__or3b_1
XFILLER_0_4_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold603 top.DUT.register\[29\]\[3\] vssd1 vssd1 vccd1 vccd1 net1719 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_116_2179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10416__S net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold614 top.DUT.register\[23\]\[1\] vssd1 vssd1 vccd1 vccd1 net1730 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold625 top.DUT.register\[24\]\[26\] vssd1 vssd1 vccd1 vccd1 net1741 sky130_fd_sc_hd__dlygate4sd3_1
Xhold636 top.DUT.register\[3\]\[2\] vssd1 vssd1 vccd1 vccd1 net1752 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07596__A2 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09990__A0 net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold647 top.DUT.register\[18\]\[13\] vssd1 vssd1 vccd1 vccd1 net1763 sky130_fd_sc_hd__dlygate4sd3_1
Xhold658 top.DUT.register\[7\]\[22\] vssd1 vssd1 vccd1 vccd1 net1774 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08793__B2 net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09961_ net1559 net223 net628 vssd1 vssd1 vccd1 vccd1 _00169_ sky130_fd_sc_hd__mux2_1
Xhold669 top.DUT.register\[24\]\[2\] vssd1 vssd1 vccd1 vccd1 net1785 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08912_ _03170_ _03499_ _03886_ vssd1 vssd1 vccd1 vccd1 _04021_ sky130_fd_sc_hd__a21bo_1
X_09892_ _04897_ _04900_ vssd1 vssd1 vccd1 vccd1 _04901_ sky130_fd_sc_hd__or2_1
XANTENNA__08545__A1 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08545__B2 net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_176_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09065__X _04140_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08843_ _01789_ _03954_ vssd1 vssd1 vccd1 vccd1 _03955_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_176_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06556__B1 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout289_A net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10151__S net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08774_ net424 _03889_ _03887_ _03873_ vssd1 vssd1 vccd1 vccd1 _03890_ sky130_fd_sc_hd__a211o_2
X_07725_ top.DUT.register\[25\]\[3\] net780 net736 top.DUT.register\[16\]\[3\] vssd1
+ vssd1 vccd1 vccd1 _02864_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_69_Left_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout456_A _01553_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07656_ top.DUT.register\[24\]\[5\] net643 net771 top.DUT.register\[10\]\[5\] _02794_
+ vssd1 vssd1 vccd1 vccd1 _02795_ sky130_fd_sc_hd__a221o_1
XFILLER_0_95_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07313__X _02452_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06607_ top.DUT.register\[30\]\[27\] net582 net509 top.DUT.register\[4\]\[27\] vssd1
+ vssd1 vccd1 vccd1 _01746_ sky130_fd_sc_hd__a22o_1
XFILLER_0_138_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout623_A net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07587_ top.a1.instruction\[18\] net794 _02725_ vssd1 vssd1 vccd1 vccd1 _02726_ sky130_fd_sc_hd__a21oi_1
X_09326_ _04387_ _04388_ vssd1 vssd1 vccd1 vccd1 _04389_ sky130_fd_sc_hd__nand2_1
X_06538_ _01672_ _01674_ _01676_ vssd1 vssd1 vccd1 vccd1 _01677_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_11_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09257_ net135 _04318_ _04323_ net810 net897 vssd1 vssd1 vccd1 vccd1 _04324_ sky130_fd_sc_hd__o221a_1
XFILLER_0_118_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08481__B1 _03598_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06469_ net787 _01602_ _01607_ vssd1 vssd1 vccd1 vccd1 _01608_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout411_X net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout509_X net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08208_ _03325_ _03345_ net276 vssd1 vssd1 vccd1 vccd1 _03346_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09188_ _04256_ _04257_ _04254_ vssd1 vssd1 vccd1 vccd1 _04259_ sky130_fd_sc_hd__o21ai_1
XPHY_EDGE_ROW_78_Left_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout992_A net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08139_ _02286_ net299 vssd1 vssd1 vccd1 vccd1 _03277_ sky130_fd_sc_hd__nand2_1
XANTENNA__10326__S net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11150_ wb.curr_state\[0\] net860 _01431_ vssd1 vssd1 vccd1 vccd1 _05081_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout780_X net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06795__B1 net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10101_ net1663 net194 net614 vssd1 vssd1 vccd1 vccd1 _00302_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_73_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11081_ net40 net864 vssd1 vssd1 vccd1 vccd1 _05046_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_164_2910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10032_ top.DUT.register\[4\]\[18\] net205 net620 vssd1 vssd1 vccd1 vccd1 _00235_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__09733__B1 net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06547__B1 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10061__S net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09703__X _04735_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input17_A DAT_I[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11983_ _05831_ _05858_ vssd1 vssd1 vccd1 vccd1 _05866_ sky130_fd_sc_hd__xnor2_1
X_13722_ clknet_leaf_98_clk _01293_ net986 vssd1 vssd1 vccd1 vccd1 top.a1.row2\[40\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_196_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10934_ net1387 net198 net591 vssd1 vssd1 vccd1 vccd1 _01095_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13345__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07511__A2 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09151__A net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_193_3339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_183_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13653_ clknet_leaf_74_clk _01232_ net1078 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[60\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_156_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10865_ net231 net1957 net594 vssd1 vssd1 vccd1 vccd1 _01026_ sky130_fd_sc_hd__mux2_1
X_12604_ clknet_leaf_0_clk _00196_ net915 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[3\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_156_659 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13584_ clknet_leaf_106_clk net1181 net970 vssd1 vssd1 vccd1 vccd1 net75 sky130_fd_sc_hd__dfrtp_1
X_10796_ net255 net1621 net600 vssd1 vssd1 vccd1 vccd1 _00957_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_155_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12535_ clknet_leaf_129_clk _00127_ net911 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[1\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_121_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_170_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12466_ clknet_leaf_106_clk _00061_ net970 vssd1 vssd1 vccd1 vccd1 top.ramstore\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_124_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11417_ _05260_ _05285_ vssd1 vssd1 vccd1 vccd1 _05300_ sky130_fd_sc_hd__nand2_1
XFILLER_0_50_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10236__S net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12397_ clknet_leaf_103_clk top.ru.next_FetchedInstr\[9\] net974 vssd1 vssd1 vccd1
+ vccd1 top.a1.instruction\[9\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__08989__X _04064_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07578__A2 net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08775__B2 _03890_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11348_ _05213_ _05218_ vssd1 vssd1 vccd1 vccd1 _05231_ sky130_fd_sc_hd__nor2_1
XANTENNA__06786__B1 net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11279_ net2255 net814 _05169_ net996 vssd1 vssd1 vccd1 vccd1 _01266_ sky130_fd_sc_hd__o211a_1
XANTENNA__08527__A1 net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13018_ clknet_leaf_5_clk _00610_ net936 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[16\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11126__A3 net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08230__A net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_176_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09613__X _04658_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07510_ top.DUT.register\[27\]\[14\] net715 net711 top.DUT.register\[11\]\[14\] vssd1
+ vssd1 vccd1 vccd1 _02649_ sky130_fd_sc_hd__a22o_1
X_08490_ net1895 net833 net803 _03618_ vssd1 vssd1 vccd1 vccd1 _00028_ sky130_fd_sc_hd__a22o_1
XANTENNA__07502__A2 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07441_ _02573_ _02575_ _02577_ _02579_ vssd1 vssd1 vccd1 vccd1 _02580_ sky130_fd_sc_hd__or4_4
XFILLER_0_187_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06710__B1 net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07372_ top.DUT.register\[16\]\[8\] net737 net699 top.DUT.register\[31\]\[8\] vssd1
+ vssd1 vccd1 vccd1 _02511_ sky130_fd_sc_hd__a22o_1
XFILLER_0_17_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09111_ top.pc\[2\] _02999_ vssd1 vssd1 vccd1 vccd1 _04186_ sky130_fd_sc_hd__nor2_1
X_06323_ top.pad.button_control.debounce_dly top.pad.button_control.debounce vssd1
+ vssd1 vccd1 vccd1 _01471_ sky130_fd_sc_hd__and2b_2
XFILLER_0_174_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_2219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_679 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09042_ _01701_ _01745_ _01921_ net495 vssd1 vssd1 vccd1 vccd1 _04117_ sky130_fd_sc_hd__and4_1
XFILLER_0_32_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06254_ net1204 net852 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedData\[15\] sky130_fd_sc_hd__and2_1
XFILLER_0_5_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_2408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_684 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10146__S net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold400 top.DUT.register\[19\]\[16\] vssd1 vssd1 vccd1 vccd1 net1516 sky130_fd_sc_hd__dlygate4sd3_1
Xhold411 top.DUT.register\[17\]\[11\] vssd1 vssd1 vccd1 vccd1 net1527 sky130_fd_sc_hd__dlygate4sd3_1
X_06185_ top.a1.hexop\[2\] top.a1.hexop\[3\] top.a1.hexop\[4\] _01420_ vssd1 vssd1
+ vccd1 vccd1 _01424_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout204_A net206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xmax_cap130 _05716_ vssd1 vssd1 vccd1 vccd1 net130 sky130_fd_sc_hd__clkbuf_2
Xhold422 top.DUT.register\[7\]\[8\] vssd1 vssd1 vccd1 vccd1 net1538 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07569__A2 net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold433 top.DUT.register\[5\]\[15\] vssd1 vssd1 vccd1 vccd1 net1549 sky130_fd_sc_hd__dlygate4sd3_1
Xhold444 top.DUT.register\[23\]\[27\] vssd1 vssd1 vccd1 vccd1 net1560 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap163 _05573_ vssd1 vssd1 vccd1 vccd1 net163 sky130_fd_sc_hd__clkbuf_1
Xhold455 top.DUT.register\[19\]\[3\] vssd1 vssd1 vccd1 vccd1 net1571 sky130_fd_sc_hd__dlygate4sd3_1
Xhold466 top.DUT.register\[8\]\[1\] vssd1 vssd1 vccd1 vccd1 net1582 sky130_fd_sc_hd__dlygate4sd3_1
Xhold477 top.DUT.register\[28\]\[5\] vssd1 vssd1 vccd1 vccd1 net1593 sky130_fd_sc_hd__dlygate4sd3_1
X_09944_ net690 _04712_ _04947_ vssd1 vssd1 vccd1 vccd1 _04948_ sky130_fd_sc_hd__and3_4
Xhold488 top.DUT.register\[6\]\[8\] vssd1 vssd1 vccd1 vccd1 net1604 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout902 net903 vssd1 vssd1 vccd1 vccd1 net902 sky130_fd_sc_hd__clkbuf_2
Xhold499 top.DUT.register\[3\]\[29\] vssd1 vssd1 vccd1 vccd1 net1615 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout913 net935 vssd1 vssd1 vccd1 vccd1 net913 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout924 net925 vssd1 vssd1 vccd1 vccd1 net924 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_55_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout935 net967 vssd1 vssd1 vccd1 vccd1 net935 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09715__B1 net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09236__A _02544_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout946 net952 vssd1 vssd1 vccd1 vccd1 net946 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08140__A _02453_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input9_A DAT_I[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09875_ net2017 net169 net631 vssd1 vssd1 vccd1 vccd1 _00146_ sky130_fd_sc_hd__mux2_1
Xfanout957 net958 vssd1 vssd1 vccd1 vccd1 net957 sky130_fd_sc_hd__clkbuf_4
Xhold1100 top.DUT.register\[10\]\[19\] vssd1 vssd1 vccd1 vccd1 net2216 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout968 net969 vssd1 vssd1 vccd1 vccd1 net968 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_209_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout573_A _01519_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1111 top.DUT.register\[12\]\[11\] vssd1 vssd1 vccd1 vccd1 net2227 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout979 net987 vssd1 vssd1 vccd1 vccd1 net979 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_146_2640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08826_ _03858_ _03938_ net308 vssd1 vssd1 vccd1 vccd1 _03939_ sky130_fd_sc_hd__mux2_1
Xhold1122 top.DUT.register\[24\]\[6\] vssd1 vssd1 vccd1 vccd1 net2238 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1133 top.DUT.register\[1\]\[21\] vssd1 vssd1 vccd1 vccd1 net2249 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1144 top.DUT.register\[19\]\[18\] vssd1 vssd1 vccd1 vccd1 net2260 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1155 top.DUT.register\[14\]\[6\] vssd1 vssd1 vccd1 vccd1 net2271 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13368__CLK clknet_leaf_128_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1166 top.DUT.register\[12\]\[26\] vssd1 vssd1 vccd1 vccd1 net2282 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_206_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08757_ net497 _03872_ vssd1 vssd1 vccd1 vccd1 _03873_ sky130_fd_sc_hd__nor2_1
Xhold1177 top.DUT.register\[30\]\[11\] vssd1 vssd1 vccd1 vccd1 net2293 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1188 top.DUT.register\[17\]\[26\] vssd1 vssd1 vccd1 vccd1 net2304 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout740_A net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout361_X net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1199 top.ramaddr\[18\] vssd1 vssd1 vccd1 vccd1 net2315 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout459_X net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07708_ top.DUT.register\[3\]\[4\] net553 net445 top.DUT.register\[1\]\[4\] _02846_
+ vssd1 vssd1 vccd1 vccd1 _02847_ sky130_fd_sc_hd__a221o_1
X_08688_ net883 top.pc\[19\] net694 _03807_ vssd1 vssd1 vccd1 vccd1 _03808_ sky130_fd_sc_hd__a22o_1
X_07639_ top.a1.instruction\[26\] net805 _02775_ _02776_ vssd1 vssd1 vccd1 vccd1 _02778_
+ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout626_X net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06701__B1 net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10650_ net195 net2040 net345 vssd1 vssd1 vccd1 vccd1 _00814_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_175_3069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09309_ _04371_ _04372_ vssd1 vssd1 vccd1 vccd1 _04373_ sky130_fd_sc_hd__nand2_1
XFILLER_0_91_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_24_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10581_ net1722 net205 net351 vssd1 vssd1 vccd1 vccd1 _00747_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12320_ top.pad.button_control.r_counter\[7\] _06122_ vssd1 vssd1 vccd1 vccd1 _06124_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_91_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_180_459 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12251_ net1195 _06080_ net979 vssd1 vssd1 vccd1 vccd1 _06082_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_106_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10056__S net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08034__B _03172_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_170_2991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11202_ _05107_ net1249 net471 vssd1 vssd1 vccd1 vccd1 _01251_ sky130_fd_sc_hd__mux2_1
XANTENNA__09845__S net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12182_ _05851_ _05083_ net847 net2263 vssd1 vssd1 vccd1 vccd1 _01290_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__06768__B1 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11133_ net58 net869 vssd1 vssd1 vccd1 vccd1 _05072_ sky130_fd_sc_hd__and2_1
XFILLER_0_101_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11108__A3 net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07980__A2 net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11064_ net1188 net864 net837 top.ramstore\[15\] vssd1 vssd1 vccd1 vccd1 _01175_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__08050__A _01722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10015_ net1280 net269 net620 vssd1 vssd1 vccd1 vccd1 _00218_ sky130_fd_sc_hd__mux2_1
XFILLER_0_204_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07732__A2 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06940__B1 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_86_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11966_ _05807_ _05848_ _05817_ vssd1 vssd1 vccd1 vccd1 _05849_ sky130_fd_sc_hd__o21ai_4
X_10917_ top.DUT.register\[30\]\[29\] net154 net481 vssd1 vssd1 vccd1 vccd1 _01078_
+ sky130_fd_sc_hd__mux2_1
X_13705_ clknet_leaf_96_clk _01276_ net984 vssd1 vssd1 vccd1 vccd1 top.a1.row2\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11897_ _05737_ _05764_ _05706_ _05736_ vssd1 vssd1 vccd1 vccd1 _05780_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_132_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_156_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13636_ clknet_leaf_75_clk _01223_ net1082 vssd1 vssd1 vccd1 vccd1 net64 sky130_fd_sc_hd__dfrtp_1
X_10848_ net2009 net173 net476 vssd1 vssd1 vccd1 vccd1 _01009_ sky130_fd_sc_hd__mux2_1
XFILLER_0_41_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13567_ clknet_leaf_104_clk _01154_ net972 vssd1 vssd1 vccd1 vccd1 top.ramload\[28\]
+ sky130_fd_sc_hd__dfrtp_2
X_10779_ net1413 net184 net484 vssd1 vssd1 vccd1 vccd1 _00940_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07799__A2 net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12518_ clknet_leaf_77_clk _00110_ net1083 vssd1 vssd1 vccd1 vccd1 top.pc\[30\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_42_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_152_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13498_ clknet_leaf_3_clk _01090_ net919 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[31\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_152_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12449_ clknet_leaf_75_clk _00045_ net1080 vssd1 vssd1 vccd1 vccd1 top.ramaddr\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11289__C _05128_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_2138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10193__C net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06759__B1 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout209 net210 vssd1 vssd1 vccd1 vccd1 net209 sky130_fd_sc_hd__clkbuf_2
X_07990_ top.DUT.register\[15\]\[31\] net708 net700 top.DUT.register\[31\]\[31\] vssd1
+ vssd1 vccd1 vccd1 _03129_ sky130_fd_sc_hd__a22o_1
XFILLER_0_5_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07971__A2 net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06941_ top.DUT.register\[13\]\[21\] net776 net704 top.DUT.register\[3\]\[21\] _02079_
+ vssd1 vssd1 vccd1 vccd1 _02080_ sky130_fd_sc_hd__a221o_1
XANTENNA__09173__A1 _02808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09660_ top.a1.halfData\[2\] _01471_ _04699_ net1086 vssd1 vssd1 vccd1 vccd1 _00117_
+ sky130_fd_sc_hd__o211a_1
X_06872_ top.DUT.register\[2\]\[18\] net561 net441 top.DUT.register\[5\]\[18\] _02010_
+ vssd1 vssd1 vccd1 vccd1 _02011_ sky130_fd_sc_hd__a221o_1
XFILLER_0_66_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07184__B1 net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_2370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08611_ net306 _03732_ _03733_ vssd1 vssd1 vccd1 vccd1 _03734_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07723__A2 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09591_ top.pc\[30\] _04620_ vssd1 vssd1 vccd1 vccd1 _04638_ sky130_fd_sc_hd__or2_1
XFILLER_0_206_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08542_ _02434_ _03667_ vssd1 vssd1 vccd1 vccd1 _03668_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_89_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08473_ net308 _03601_ vssd1 vssd1 vccd1 vccd1 _03602_ sky130_fd_sc_hd__nand2_1
XFILLER_0_159_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11283__A2 _05132_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07424_ top.DUT.register\[25\]\[9\] net778 net711 top.DUT.register\[11\]\[9\] vssd1
+ vssd1 vccd1 vccd1 _02563_ sky130_fd_sc_hd__a22o_1
XFILLER_0_9_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_175_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_174_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07355_ top.DUT.register\[18\]\[8\] net547 net504 top.DUT.register\[27\]\[8\] vssd1
+ vssd1 vccd1 vccd1 _02494_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout1063_A net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout419_A net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06306_ _01333_ _01329_ vssd1 vssd1 vccd1 vccd1 _01462_ sky130_fd_sc_hd__and2b_1
X_07286_ top.DUT.register\[14\]\[13\] net732 net704 top.DUT.register\[3\]\[13\] _02424_
+ vssd1 vssd1 vccd1 vccd1 _02425_ sky130_fd_sc_hd__a221o_1
XANTENNA__08135__A _02409_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06998__B1 net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09025_ _02178_ _02221_ _02611_ _02655_ vssd1 vssd1 vccd1 vccd1 _04100_ sky130_fd_sc_hd__or4_1
X_06237_ top.ramload\[31\] net858 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedInstr\[31\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_41_660 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_479 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold230 top.DUT.register\[17\]\[4\] vssd1 vssd1 vccd1 vccd1 net1346 sky130_fd_sc_hd__dlygate4sd3_1
Xhold241 top.DUT.register\[5\]\[0\] vssd1 vssd1 vccd1 vccd1 net1357 sky130_fd_sc_hd__dlygate4sd3_1
X_06168_ _01409_ vssd1 vssd1 vccd1 vccd1 _01410_ sky130_fd_sc_hd__inv_2
XFILLER_0_13_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold252 top.DUT.register\[6\]\[14\] vssd1 vssd1 vccd1 vccd1 net1368 sky130_fd_sc_hd__dlygate4sd3_1
Xhold263 top.ramaddr\[11\] vssd1 vssd1 vccd1 vccd1 net1379 sky130_fd_sc_hd__dlygate4sd3_1
Xhold274 top.DUT.register\[13\]\[24\] vssd1 vssd1 vccd1 vccd1 net1390 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold285 top.DUT.register\[28\]\[21\] vssd1 vssd1 vccd1 vccd1 net1401 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10604__S net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold296 top.DUT.register\[4\]\[21\] vssd1 vssd1 vccd1 vccd1 net1412 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout710 _01638_ vssd1 vssd1 vccd1 vccd1 net710 sky130_fd_sc_hd__clkbuf_8
Xfanout721 _01635_ vssd1 vssd1 vccd1 vccd1 net721 sky130_fd_sc_hd__buf_2
XANTENNA__13190__CLK clknet_leaf_40_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout732 _01627_ vssd1 vssd1 vccd1 vccd1 net732 sky130_fd_sc_hd__clkbuf_8
X_09927_ _04931_ _04932_ vssd1 vssd1 vccd1 vccd1 _04933_ sky130_fd_sc_hd__nor2_1
Xfanout743 _01623_ vssd1 vssd1 vccd1 vccd1 net743 sky130_fd_sc_hd__buf_2
Xfanout754 _01620_ vssd1 vssd1 vccd1 vccd1 net754 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout955_A net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout576_X net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout765 _01616_ vssd1 vssd1 vccd1 vccd1 net765 sky130_fd_sc_hd__buf_4
Xfanout776 net777 vssd1 vssd1 vccd1 vccd1 net776 sky130_fd_sc_hd__buf_4
Xfanout787 _01592_ vssd1 vssd1 vccd1 vccd1 net787 sky130_fd_sc_hd__buf_2
X_09858_ _04861_ _04862_ _04864_ vssd1 vssd1 vccd1 vccd1 _04870_ sky130_fd_sc_hd__o21ai_1
XANTENNA__06877__X _02016_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07175__B1 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout798 _04150_ vssd1 vssd1 vccd1 vccd1 net798 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08911__A1 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08809_ _01875_ net433 net501 _01876_ _03883_ vssd1 vssd1 vccd1 vccd1 _03923_ sky130_fd_sc_hd__a221o_1
X_09789_ top.pc\[17\] _04438_ vssd1 vssd1 vccd1 vccd1 _04808_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout743_X net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11820_ top.a1.dataIn\[6\] _05699_ _05700_ _05701_ vssd1 vssd1 vccd1 vccd1 _05703_
+ sky130_fd_sc_hd__a2bb2o_2
XTAP_TAPCELL_ROW_1_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_68_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11751_ _05603_ _05606_ _05619_ _05605_ vssd1 vssd1 vccd1 vccd1 _05634_ sky130_fd_sc_hd__o31a_1
XFILLER_0_138_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11274__A2 _05132_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_159_2831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_80_clk clknet_4_6__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_80_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_166_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10702_ net2238 net241 net334 vssd1 vssd1 vccd1 vccd1 _00863_ sky130_fd_sc_hd__mux2_1
XFILLER_0_166_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11682_ _05563_ _05564_ vssd1 vssd1 vccd1 vccd1 _05565_ sky130_fd_sc_hd__nor2_1
XFILLER_0_36_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13421_ clknet_leaf_51_clk _01013_ net1056 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[28\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_10633_ net256 net1953 net344 vssd1 vssd1 vccd1 vccd1 _00797_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_180_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_181_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13352_ clknet_leaf_25_clk _00944_ net1009 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[26\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_181_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10564_ net1525 net270 net351 vssd1 vssd1 vccd1 vccd1 _00730_ sky130_fd_sc_hd__mux2_1
XANTENNA__06989__B1 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12303_ top.pad.button_control.r_counter\[0\] net1265 net790 vssd1 vssd1 vccd1 vccd1
+ _06113_ sky130_fd_sc_hd__o21ai_1
XANTENNA__06491__C _01607_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13283_ clknet_leaf_58_clk _00875_ net1076 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[24\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_10495_ _04712_ _04947_ net400 vssd1 vssd1 vccd1 vccd1 _04987_ sky130_fd_sc_hd__and3_1
X_12234_ _06070_ _06071_ vssd1 vssd1 vccd1 vccd1 _01319_ sky130_fd_sc_hd__nor2_1
XFILLER_0_32_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08699__B _03441_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10514__S net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12165_ net2093 net846 net796 _06046_ vssd1 vssd1 vccd1 vccd1 _01275_ sky130_fd_sc_hd__a22o_1
XFILLER_0_102_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11116_ net905 net1708 net860 _05063_ vssd1 vssd1 vccd1 vccd1 _01209_ sky130_fd_sc_hd__a31o_1
X_12096_ top.a1.dataIn\[3\] _05948_ vssd1 vssd1 vccd1 vccd1 _05979_ sky130_fd_sc_hd__and2_1
XANTENNA__09307__C _04370_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_207_3544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_207_3555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11047_ net1133 net864 net837 vssd1 vssd1 vccd1 vccd1 _01158_ sky130_fd_sc_hd__a21o_1
XANTENNA__09026__D _03185_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07705__A2 net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput9 DAT_I[16] vssd1 vssd1 vccd1 vccd1 net9 sky130_fd_sc_hd__clkbuf_1
XANTENNA__06913__B1 net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_207_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_204_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12998_ clknet_leaf_38_clk _00590_ net1054 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[15\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_148_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07124__A _02242_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11265__A2 _05136_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11949_ _05796_ _05819_ vssd1 vssd1 vccd1 vccd1 _05832_ sky130_fd_sc_hd__and2_1
XANTENNA__09863__C1 _04874_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_71_clk clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_71_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_156_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_157_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_144_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11017__A2 net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13619_ clknet_leaf_72_clk _01206_ net1085 vssd1 vssd1 vccd1 vccd1 net45 sky130_fd_sc_hd__dfrtp_1
XANTENNA__10225__A0 net156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_99_1933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08969__B2 net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07140_ top.DUT.register\[9\]\[11\] net467 net507 top.DUT.register\[4\]\[11\] vssd1
+ vssd1 vccd1 vccd1 _02279_ sky130_fd_sc_hd__a22o_1
XFILLER_0_109_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_172_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13569__Q top.ramload\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07071_ top.DUT.register\[29\]\[22\] net722 net703 top.DUT.register\[3\]\[22\] vssd1
+ vssd1 vccd1 vccd1 _02210_ sky130_fd_sc_hd__a22o_1
XFILLER_0_180_790 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_695 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_140_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10424__S net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08402__B net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08553__A1_N net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07973_ top.DUT.register\[15\]\[31\] net681 net677 top.DUT.register\[31\]\[31\] vssd1
+ vssd1 vccd1 vccd1 _03112_ sky130_fd_sc_hd__a22o_1
XANTENNA__09146__A1 _01505_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09712_ net826 _04252_ vssd1 vssd1 vccd1 vccd1 _04742_ sky130_fd_sc_hd__nor2_1
X_06924_ top.DUT.register\[20\]\[21\] net565 net464 top.DUT.register\[13\]\[21\] _02062_
+ vssd1 vssd1 vccd1 vccd1 _02063_ sky130_fd_sc_hd__a221o_1
XANTENNA__07157__B1 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09643_ _04674_ _04684_ _01471_ vssd1 vssd1 vccd1 vccd1 _04685_ sky130_fd_sc_hd__o21ai_1
X_06855_ top.DUT.register\[30\]\[19\] net761 net748 top.DUT.register\[17\]\[19\] vssd1
+ vssd1 vccd1 vccd1 _01994_ sky130_fd_sc_hd__a22o_1
XFILLER_0_179_323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout369_A net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09574_ _04609_ _04621_ vssd1 vssd1 vccd1 vccd1 _04622_ sky130_fd_sc_hd__nor2_1
X_06786_ top.DUT.register\[8\]\[17\] net540 net440 top.DUT.register\[5\]\[17\] _01924_
+ vssd1 vssd1 vccd1 vccd1 _01925_ sky130_fd_sc_hd__a221o_1
X_08525_ _03453_ _03651_ net296 vssd1 vssd1 vccd1 vccd1 _03652_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_26_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout536_A _01541_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_62_clk clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_62_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_clkbuf_leaf_60_clk_A clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08456_ _03328_ _03534_ vssd1 vssd1 vccd1 vccd1 _03586_ sky130_fd_sc_hd__nor2_1
XFILLER_0_203_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_172_3028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07407_ _02359_ _02501_ _02545_ _01580_ vssd1 vssd1 vccd1 vccd1 _02546_ sky130_fd_sc_hd__o211a_1
XANTENNA__06683__A2 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08387_ _03516_ _03518_ vssd1 vssd1 vccd1 vccd1 _03519_ sky130_fd_sc_hd__and2_2
XANTENNA_fanout324_X net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout703_A _01642_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07338_ _02476_ vssd1 vssd1 vccd1 vccd1 _02477_ sky130_fd_sc_hd__inv_2
XFILLER_0_190_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_154_2750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_75_clk_A clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_154_2761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07269_ _02401_ _02403_ _02405_ _02407_ vssd1 vssd1 vccd1 vccd1 _02408_ sky130_fd_sc_hd__or4_4
X_09008_ _03928_ _04081_ vssd1 vssd1 vccd1 vccd1 _04083_ sky130_fd_sc_hd__or2_1
XFILLER_0_60_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10280_ net1312 net217 net386 vssd1 vssd1 vccd1 vccd1 _00458_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout693_X net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09385__A1 net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10334__S net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07396__B1 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08312__B net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout860_X net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout540 _01540_ vssd1 vssd1 vccd1 vccd1 net540 sky130_fd_sc_hd__clkbuf_4
Xfanout551 _01535_ vssd1 vssd1 vccd1 vccd1 net551 sky130_fd_sc_hd__buf_4
XANTENNA__09137__A1 top.pc\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout562 _01532_ vssd1 vssd1 vccd1 vccd1 net562 sky130_fd_sc_hd__buf_4
Xfanout573 _01519_ vssd1 vssd1 vccd1 vccd1 net573 sky130_fd_sc_hd__buf_6
XANTENNA__07148__B1 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_13_clk_A clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout584 _01513_ vssd1 vssd1 vccd1 vccd1 net584 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09688__A2 net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout595 _04966_ vssd1 vssd1 vccd1 vccd1 net595 sky130_fd_sc_hd__buf_4
XANTENNA__09424__A net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12921_ clknet_leaf_14_clk _00513_ net960 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[13\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12852_ clknet_leaf_57_clk _00444_ net1075 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[11\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_202_3474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_201_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_197_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_14_Left_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11803_ _05636_ _05683_ _05632_ vssd1 vssd1 vccd1 vccd1 _05686_ sky130_fd_sc_hd__a21o_1
XFILLER_0_185_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12783_ clknet_leaf_41_clk _00375_ net1045 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[8\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_139_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_185_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_28_clk_A clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_53_clk clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_53_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_68_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_302 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11734_ _05574_ _05611_ _05615_ _05616_ vssd1 vssd1 vccd1 vccd1 _05617_ sky130_fd_sc_hd__nor4_1
XANTENNA__09430__Y _04487_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07320__B1 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06674__A2 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11665_ _05546_ _05547_ vssd1 vssd1 vccd1 vccd1 _05548_ sky130_fd_sc_hd__nor2_1
XFILLER_0_193_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10509__S net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10616_ net200 net1929 net348 vssd1 vssd1 vccd1 vccd1 _00781_ sky130_fd_sc_hd__mux2_1
X_13404_ clknet_leaf_0_clk _00996_ net915 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[28\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11596_ _05443_ _05478_ vssd1 vssd1 vccd1 vccd1 _05479_ sky130_fd_sc_hd__nand2_1
XFILLER_0_153_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13335_ clknet_leaf_2_clk _00927_ net919 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[26\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_141_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10547_ net1341 net215 _04989_ vssd1 vssd1 vccd1 vccd1 _00714_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_23_Left_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13266_ clknet_leaf_31_clk _00858_ net1021 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[24\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_10478_ net1481 net188 net362 vssd1 vssd1 vccd1 vccd1 _00648_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_94_1852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_1863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12217_ top.lcd.cnt_20ms\[1\] top.lcd.cnt_20ms\[0\] top.lcd.cnt_20ms\[2\] vssd1 vssd1
+ vccd1 vccd1 _06061_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10244__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_714 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13197_ clknet_leaf_42_clk _00789_ net1064 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[21\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09318__B _04370_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07387__B1 net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12148_ _06011_ _06022_ _06024_ vssd1 vssd1 vccd1 vccd1 _06031_ sky130_fd_sc_hd__a21o_1
XANTENNA__09128__A1 top.pc\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12079_ _05957_ _05961_ vssd1 vssd1 vccd1 vccd1 _05962_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_10_Right_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_189_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_108_2059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_139_Right_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06640_ top.DUT.register\[13\]\[27\] net775 net764 top.DUT.register\[9\]\[27\] vssd1
+ vssd1 vccd1 vccd1 _01779_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_32_Left_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_188_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06571_ top.DUT.register\[3\]\[28\] net554 net457 top.DUT.register\[25\]\[28\] _01709_
+ vssd1 vssd1 vccd1 vccd1 _01710_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_121_2259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_44_clk clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_44_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_188_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08310_ _03413_ _03422_ _03412_ vssd1 vssd1 vccd1 vccd1 _03445_ sky130_fd_sc_hd__a21bo_1
X_09290_ _04353_ _04354_ vssd1 vssd1 vccd1 vccd1 _04355_ sky130_fd_sc_hd__nor2_1
XANTENNA__06693__A _01809_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07311__B1 net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10997__B2 top.a1.dataIn\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08241_ _03224_ _03228_ vssd1 vssd1 vccd1 vccd1 _03378_ sky130_fd_sc_hd__nand2_1
XFILLER_0_172_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06665__A2 net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10419__S net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_1992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08172_ _01940_ net299 vssd1 vssd1 vccd1 vccd1 _03310_ sky130_fd_sc_hd__nand2_1
XFILLER_0_70_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07123_ net807 net412 net437 vssd1 vssd1 vccd1 vccd1 _02262_ sky130_fd_sc_hd__o21ai_1
XANTENNA__06417__A2 net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_41_Left_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_2480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_2491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07054_ top.DUT.register\[26\]\[22\] net527 net507 top.DUT.register\[4\]\[22\] vssd1
+ vssd1 vccd1 vccd1 _02193_ sky130_fd_sc_hd__a22o_1
XANTENNA__09509__A _01854_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput110 net110 vssd1 vssd1 vccd1 vccd1 WE_O sky130_fd_sc_hd__buf_2
XANTENNA__07090__A2 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput121 net121 vssd1 vssd1 vccd1 vccd1 gpio_out[6] sky130_fd_sc_hd__buf_2
XFILLER_0_23_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_164 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09367__A1 net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10154__S net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07378__B1 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07917__A2 _02703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09005__A_N _03750_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07956_ _01790_ _03094_ vssd1 vssd1 vccd1 vccd1 _03095_ sky130_fd_sc_hd__nor2_1
X_06907_ net808 _02045_ net438 vssd1 vssd1 vccd1 vccd1 _02046_ sky130_fd_sc_hd__o21a_1
XPHY_EDGE_ROW_50_Left_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07887_ top.DUT.register\[2\]\[1\] net561 net520 top.DUT.register\[10\]\[1\] vssd1
+ vssd1 vccd1 vccd1 _03026_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout274_X net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout653_A _01610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_106_Right_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06838_ top.DUT.register\[2\]\[19\] net562 net461 top.DUT.register\[17\]\[19\] _01976_
+ vssd1 vssd1 vccd1 vccd1 _01977_ sky130_fd_sc_hd__a221o_1
X_09626_ _04670_ vssd1 vssd1 vccd1 vccd1 _04671_ sky130_fd_sc_hd__inv_2
XANTENNA__07550__B1 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_65_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09557_ _01722_ _04605_ vssd1 vssd1 vccd1 vccd1 _04606_ sky130_fd_sc_hd__nand2_1
X_06769_ top.DUT.register\[4\]\[24\] net670 net732 top.DUT.register\[14\]\[24\] vssd1
+ vssd1 vccd1 vccd1 _01908_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout441_X net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_35_clk clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_35_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout539_X net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08508_ _02386_ _03614_ vssd1 vssd1 vccd1 vccd1 _03636_ sky130_fd_sc_hd__nor2_1
X_09488_ _04537_ _04540_ vssd1 vssd1 vccd1 vccd1 _04541_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_65_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07302__B1 net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08439_ net886 top.pc\[8\] net697 _03569_ vssd1 vssd1 vccd1 vccd1 _03570_ sky130_fd_sc_hd__a22o_1
XANTENNA__06656__A2 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10329__S net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout706_X net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_519 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08307__B net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11450_ top.a1.dataIn\[17\] _05254_ _05293_ vssd1 vssd1 vccd1 vccd1 _05333_ sky130_fd_sc_hd__or3_1
XFILLER_0_18_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10401_ net1539 net257 net370 vssd1 vssd1 vccd1 vccd1 _00573_ sky130_fd_sc_hd__mux2_1
X_11381_ _05226_ _05257_ vssd1 vssd1 vccd1 vccd1 _05264_ sky130_fd_sc_hd__xor2_2
XFILLER_0_104_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_150_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13120_ clknet_leaf_115_clk _00712_ net964 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[19\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_10332_ net2177 net259 net379 vssd1 vssd1 vccd1 vccd1 _00508_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08323__A _03342_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_185_3219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13051_ clknet_leaf_126_clk _00643_ net929 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[17\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_10263_ net1751 net145 net385 vssd1 vssd1 vccd1 vccd1 _00441_ sky130_fd_sc_hd__mux2_1
XANTENNA__09138__B _02904_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10064__S net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07369__B1 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12002_ _05862_ net126 _05864_ vssd1 vssd1 vccd1 vccd1 _05885_ sky130_fd_sc_hd__a21o_1
X_10194_ net602 _04973_ net594 vssd1 vssd1 vccd1 vccd1 _04974_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_167_2952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08977__B net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08581__A2 top.pc\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_204_3503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout370 net372 vssd1 vssd1 vccd1 vccd1 net370 sky130_fd_sc_hd__buf_6
Xfanout381 net384 vssd1 vssd1 vccd1 vccd1 net381 sky130_fd_sc_hd__buf_6
Xfanout392 _04977_ vssd1 vssd1 vccd1 vccd1 net392 sky130_fd_sc_hd__clkbuf_8
X_12904_ clknet_leaf_7_clk _00496_ net946 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[12\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06895__A2 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12835_ clknet_leaf_53_clk _00427_ net1038 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[10\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_124_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_26_clk clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_26_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_69_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_185_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12766_ clknet_leaf_18_clk _00358_ net1031 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[8\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_655 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11717_ _05598_ _05599_ vssd1 vssd1 vccd1 vccd1 _05600_ sky130_fd_sc_hd__nand2_1
XANTENNA__10239__S net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12697_ clknet_leaf_14_clk _00289_ net955 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[6\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_182_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_140_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09046__B1 _03737_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11648_ _05514_ _05515_ _05507_ vssd1 vssd1 vccd1 vccd1 _05531_ sky130_fd_sc_hd__a21bo_1
Xinput12 DAT_I[19] vssd1 vssd1 vccd1 vccd1 net12 sky130_fd_sc_hd__buf_1
Xinput23 DAT_I[29] vssd1 vssd1 vccd1 vccd1 net23 sky130_fd_sc_hd__clkbuf_1
Xinput34 en vssd1 vssd1 vccd1 vccd1 net34 sky130_fd_sc_hd__clkbuf_2
X_11579_ _05447_ _05452_ _05460_ vssd1 vssd1 vccd1 vccd1 _05462_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_3_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold807 top.ramaddr\[26\] vssd1 vssd1 vccd1 vccd1 net1923 sky130_fd_sc_hd__dlygate4sd3_1
X_13318_ clknet_leaf_32_clk _00910_ net1044 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[25\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold818 top.DUT.register\[8\]\[0\] vssd1 vssd1 vccd1 vccd1 net1934 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07072__A2 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold829 top.DUT.register\[10\]\[12\] vssd1 vssd1 vccd1 vccd1 net1945 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_208_Right_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13249_ clknet_leaf_16_clk _00841_ net963 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[23\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11156__A1 top.a1.halfData\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_460 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07810_ top.a1.instruction\[21\] _01507_ net793 top.a1.instruction\[13\] _02948_
+ vssd1 vssd1 vccd1 vccd1 _02949_ sky130_fd_sc_hd__a221o_1
X_08790_ net281 _03204_ vssd1 vssd1 vccd1 vccd1 _03905_ sky130_fd_sc_hd__or2_1
XANTENNA__10702__S net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07780__B1 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07741_ _02857_ _02878_ net823 vssd1 vssd1 vccd1 vccd1 _02880_ sky130_fd_sc_hd__mux2_4
XFILLER_0_79_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07672_ top.DUT.register\[25\]\[4\] net780 net637 top.DUT.register\[6\]\[4\] vssd1
+ vssd1 vccd1 vccd1 _02811_ sky130_fd_sc_hd__a22o_1
XANTENNA__07532__B1 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09411_ _04456_ _04457_ _04454_ vssd1 vssd1 vccd1 vccd1 _04469_ sky130_fd_sc_hd__o21ai_1
X_06623_ top.DUT.register\[17\]\[27\] net461 net525 top.DUT.register\[11\]\[27\] _01761_
+ vssd1 vssd1 vccd1 vccd1 _01762_ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_17_clk clknet_4_12__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_17_clk
+ sky130_fd_sc_hd__clkbuf_8
X_09342_ _02580_ _02589_ _04403_ vssd1 vssd1 vccd1 vccd1 _04404_ sky130_fd_sc_hd__o21a_1
X_06554_ top.DUT.register\[1\]\[29\] net756 net712 top.DUT.register\[11\]\[29\] vssd1
+ vssd1 vccd1 vccd1 _01693_ sky130_fd_sc_hd__a22o_1
XFILLER_0_192_605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06638__A2 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09273_ _02286_ _04337_ vssd1 vssd1 vccd1 vccd1 _04339_ sky130_fd_sc_hd__nor2_1
XANTENNA__07835__A1 net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06485_ _01598_ _01607_ net792 vssd1 vssd1 vccd1 vccd1 _01624_ sky130_fd_sc_hd__and3b_4
XANTENNA__10149__S net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_2520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08224_ net292 _03226_ net304 vssd1 vssd1 vccd1 vccd1 _03361_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_60_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08155_ _02773_ net300 vssd1 vssd1 vccd1 vccd1 _03293_ sky130_fd_sc_hd__nand2_1
XFILLER_0_99_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_546 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07599__B1 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07106_ top.DUT.register\[15\]\[16\] net707 net699 top.DUT.register\[31\]\[16\] vssd1
+ vssd1 vccd1 vccd1 _02245_ sky130_fd_sc_hd__a22o_1
X_08086_ _02899_ net330 vssd1 vssd1 vccd1 vccd1 _03225_ sky130_fd_sc_hd__nand2_1
XANTENNA__07063__A2 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08143__A _02329_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07037_ net808 _02175_ net438 vssd1 vssd1 vccd1 vccd1 _02176_ sky130_fd_sc_hd__o21a_1
XANTENNA__06810__A2 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11147__A1 _02952_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09526__X _04577_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08430__X _03561_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout391_X net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout770_A _01614_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout489_X net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout868_A net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09760__A1 _04386_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10612__S net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_149_2682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_180_3149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08988_ _03256_ _03350_ vssd1 vssd1 vccd1 vccd1 _04063_ sky130_fd_sc_hd__nand2b_1
X_07939_ _02049_ _03077_ _03076_ vssd1 vssd1 vccd1 vccd1 _03078_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout656_X net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_162_2871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10950_ net2149 net149 net591 vssd1 vssd1 vccd1 vccd1 _01111_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_162_2882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07523__B1 net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09702__A net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09609_ net134 _04650_ _04651_ _04654_ vssd1 vssd1 vccd1 vccd1 _04655_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_211_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10881_ net170 net2105 net595 vssd1 vssd1 vccd1 vccd1 _01042_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout823_X net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_195_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12620_ clknet_leaf_62_clk _00212_ net1088 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[3\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_211_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09276__B1 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_195_3370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09815__A2 net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06629__A2 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12551_ clknet_leaf_6_clk _00143_ net937 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[1\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_182_126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10059__S net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_603 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11502_ _05274_ _05308_ vssd1 vssd1 vccd1 vccd1 _05385_ sky130_fd_sc_hd__xor2_1
XFILLER_0_19_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12482_ clknet_leaf_64_clk _00077_ net1092 vssd1 vssd1 vccd1 vccd1 top.ramstore\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_191_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_362 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11433_ _05274_ _05315_ vssd1 vssd1 vccd1 vccd1 _05316_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_78_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09579__B2 _04051_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11364_ top.a1.dataIn\[28\] _05239_ top.a1.dataIn\[29\] vssd1 vssd1 vccd1 vccd1 _05247_
+ sky130_fd_sc_hd__o21a_1
XANTENNA__07054__A2 net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10315_ net185 net1686 net382 vssd1 vssd1 vccd1 vccd1 _00492_ sky130_fd_sc_hd__mux2_1
X_13103_ clknet_leaf_21_clk _00695_ net1033 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[18\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13274__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11295_ top.a1.row1\[12\] _05123_ _05131_ vssd1 vssd1 vccd1 vccd1 _05184_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_210_3595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11138__A1 net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13034_ clknet_leaf_115_clk _00626_ net957 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[16\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_10246_ net226 net2209 net390 vssd1 vssd1 vccd1 vccd1 _00425_ sky130_fd_sc_hd__mux2_1
XANTENNA__08003__A1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08554__A2 net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08952__A1_N _02521_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10522__S net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10177_ net1912 net143 net604 vssd1 vssd1 vccd1 vccd1 _00376_ sky130_fd_sc_hd__mux2_1
XANTENNA__06565__A1 top.DUT.register\[6\]\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08306__A2 _03440_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_105_2018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07514__B1 net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08967__A1_N _02131_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_198_292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12818_ clknet_leaf_23_clk _00410_ net1021 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[10\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13798_ clknet_leaf_68_clk _01367_ vssd1 vssd1 vccd1 vccd1 top.pad.button_control.r_counter\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_33_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12749_ clknet_leaf_43_clk _00341_ net1063 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[7\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_155_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_1940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_1951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09758__S net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06270_ top.ramload\[31\] net853 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedData\[31\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_170_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_42_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold604 top.DUT.register\[13\]\[21\] vssd1 vssd1 vccd1 vccd1 net1720 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07045__A2 net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold615 top.DUT.register\[3\]\[10\] vssd1 vssd1 vccd1 vccd1 net1731 sky130_fd_sc_hd__dlygate4sd3_1
Xhold626 top.DUT.register\[18\]\[4\] vssd1 vssd1 vccd1 vccd1 net1742 sky130_fd_sc_hd__dlygate4sd3_1
Xhold637 top.DUT.register\[14\]\[9\] vssd1 vssd1 vccd1 vccd1 net1753 sky130_fd_sc_hd__dlygate4sd3_1
Xhold648 top.DUT.register\[12\]\[21\] vssd1 vssd1 vccd1 vccd1 net1764 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08793__A2 _03902_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11101__B net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12657__RESET_B net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09960_ net1465 net191 net628 vssd1 vssd1 vccd1 vccd1 _00168_ sky130_fd_sc_hd__mux2_1
Xhold659 top.DUT.register\[3\]\[3\] vssd1 vssd1 vccd1 vccd1 net1775 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_6_clk clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_6_clk
+ sky130_fd_sc_hd__clkbuf_8
X_08911_ net274 _03859_ _04016_ _04019_ vssd1 vssd1 vccd1 vccd1 _04020_ sky130_fd_sc_hd__a211o_1
X_09891_ _04898_ _04899_ vssd1 vssd1 vccd1 vccd1 _04900_ sky130_fd_sc_hd__and2b_1
X_08842_ _01833_ _03935_ _01831_ vssd1 vssd1 vccd1 vccd1 _03954_ sky130_fd_sc_hd__o21ba_1
XANTENNA__10432__S net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_191_Right_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07753__B1 net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08773_ _02136_ _03888_ vssd1 vssd1 vccd1 vccd1 _03889_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_26_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12791__CLK clknet_leaf_128_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07724_ top.DUT.register\[29\]\[3\] net724 _02860_ _02862_ vssd1 vssd1 vccd1 vccd1
+ _02863_ sky130_fd_sc_hd__a211o_1
XANTENNA__11301__A1 top.lcd.nextState\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07741__S net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09522__A top.pc\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06859__A2 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07655_ top.DUT.register\[17\]\[5\] net746 net742 top.DUT.register\[2\]\[5\] vssd1
+ vssd1 vccd1 vccd1 _02794_ sky130_fd_sc_hd__a22o_1
XFILLER_0_189_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout351_A net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1093_A net1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06606_ _01743_ _01744_ vssd1 vssd1 vccd1 vccd1 _01745_ sky130_fd_sc_hd__nand2b_2
XANTENNA_fanout449_A _01562_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07586_ top.a1.instruction\[26\] net789 vssd1 vssd1 vccd1 vccd1 _02725_ sky130_fd_sc_hd__and2_1
XFILLER_0_48_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09325_ _02623_ _02632_ _04386_ vssd1 vssd1 vccd1 vccd1 _04388_ sky130_fd_sc_hd__or3_1
X_06537_ top.DUT.register\[13\]\[29\] net464 net521 top.DUT.register\[10\]\[29\] _01675_
+ vssd1 vssd1 vccd1 vccd1 _01676_ sky130_fd_sc_hd__a221o_1
XFILLER_0_47_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_146_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout616_A _04954_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09256_ _04321_ _04322_ vssd1 vssd1 vccd1 vccd1 _04323_ sky130_fd_sc_hd__xnor2_1
XANTENNA_clkbuf_4_10__f_clk_A clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08481__A1 _03370_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06468_ top.a1.instruction\[22\] top.a1.instruction\[23\] vssd1 vssd1 vccd1 vccd1
+ _01607_ sky130_fd_sc_hd__and2_2
XFILLER_0_90_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07284__A2 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08425__X _03556_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08207_ net330 _03122_ vssd1 vssd1 vccd1 vccd1 _03345_ sky130_fd_sc_hd__or2_1
XFILLER_0_141_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06492__B1 net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09187_ _04254_ _04256_ _04257_ vssd1 vssd1 vccd1 vccd1 _04258_ sky130_fd_sc_hd__or3_1
XANTENNA__10607__S net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout404_X net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06399_ top.DUT.register\[2\]\[30\] net561 net556 top.DUT.register\[28\]\[30\] _01537_
+ vssd1 vssd1 vccd1 vccd1 _01538_ sky130_fd_sc_hd__a221o_1
X_08138_ _03272_ _03275_ net289 vssd1 vssd1 vccd1 vccd1 _03276_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_522 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout985_A net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08751__A2_N _03861_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11011__B net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08069_ _03206_ _03207_ vssd1 vssd1 vccd1 vccd1 _03208_ sky130_fd_sc_hd__nand2_1
XANTENNA__07983__Y _03122_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10100_ net1506 net201 net613 vssd1 vssd1 vccd1 vccd1 _00301_ sky130_fd_sc_hd__mux2_1
XANTENNA__07992__B1 net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11080_ net97 net871 net835 net1149 vssd1 vssd1 vccd1 vccd1 _01191_ sky130_fd_sc_hd__a22o_1
XFILLER_0_101_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout773_X net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_164_2900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09733__A1 _03594_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10031_ net1673 net217 net622 vssd1 vssd1 vccd1 vccd1 _00234_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_164_2911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10342__S net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12123__A top.a1.dataIn\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07744__B1 net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11982_ top.a1.dataIn\[4\] _05835_ _05852_ _05861_ vssd1 vssd1 vccd1 vccd1 _05865_
+ sky130_fd_sc_hd__or4b_2
X_13721_ clknet_leaf_98_clk _01292_ net986 vssd1 vssd1 vccd1 vccd1 top.a1.row2\[35\]
+ sky130_fd_sc_hd__dfrtp_1
X_10933_ net1475 net208 net591 vssd1 vssd1 vccd1 vccd1 _01094_ sky130_fd_sc_hd__mux2_1
XANTENNA__08319__Y _03454_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10864_ net235 net2173 net595 vssd1 vssd1 vccd1 vccd1 _01025_ sky130_fd_sc_hd__mux2_1
X_13652_ clknet_leaf_74_clk _01231_ net1078 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[61\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_155_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12603_ clknet_leaf_126_clk _00195_ net929 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[3\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11056__B1 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13583_ clknet_leaf_106_clk net1194 net968 vssd1 vssd1 vccd1 vccd1 net74 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10795_ net261 net2205 net601 vssd1 vssd1 vccd1 vccd1 _00956_ sky130_fd_sc_hd__mux2_1
X_12534_ clknet_leaf_4_clk _00126_ net940 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[1\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07275__A2 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_163_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10517__S net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12465_ clknet_leaf_106_clk _00060_ net968 vssd1 vssd1 vccd1 vccd1 top.ramstore\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_151_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07027__A2 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11416_ _05292_ _05297_ vssd1 vssd1 vccd1 vccd1 _05299_ sky130_fd_sc_hd__nor2_1
X_12396_ clknet_leaf_102_clk top.ru.next_FetchedInstr\[8\] net974 vssd1 vssd1 vccd1
+ vccd1 top.a1.instruction\[8\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_22_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_270 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11347_ _05228_ _05229_ vssd1 vssd1 vccd1 vccd1 _05230_ sky130_fd_sc_hd__nand2_1
XANTENNA__08775__A2 top.pc\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09607__A net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11278_ _05121_ _05164_ _05166_ _05168_ vssd1 vssd1 vccd1 vccd1 _05169_ sky130_fd_sc_hd__or4_1
XANTENNA__08527__A2 _03122_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09724__A1 _04172_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10229_ _04947_ _04958_ net399 vssd1 vssd1 vccd1 vccd1 _04977_ sky130_fd_sc_hd__nand3_1
X_13017_ clknet_leaf_15_clk _00609_ net959 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[16\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10252__S net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07735__B1 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1 top.ramload\[8\] vssd1 vssd1 vccd1 vccd1 net1117 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_6_Left_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_169_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_18_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07440_ top.DUT.register\[23\]\[15\] net573 net556 top.DUT.register\[28\]\[15\] _02578_
+ vssd1 vssd1 vccd1 vccd1 _02579_ sky130_fd_sc_hd__a221o_1
XFILLER_0_76_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_8_Right_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11047__B1 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07371_ top.DUT.register\[20\]\[8\] net664 net739 top.DUT.register\[12\]\[8\] _02507_
+ vssd1 vssd1 vccd1 vccd1 _02510_ sky130_fd_sc_hd__a221o_1
XFILLER_0_174_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06972__Y _02111_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09110_ _01406_ _03000_ vssd1 vssd1 vccd1 vccd1 _04185_ sky130_fd_sc_hd__nor2_1
X_06322_ top.pad.count\[0\] top.pad.count\[1\] vssd1 vssd1 vccd1 vccd1 net120 sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_118_2209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07266__A2 net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08463__B2 net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09041_ _01790_ _01834_ _02754_ _03519_ vssd1 vssd1 vccd1 vccd1 _04116_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_40_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06253_ top.ramload\[14\] net852 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedData\[14\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_182_490 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10427__S net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07018__A2 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_2409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold401 top.DUT.register\[21\]\[26\] vssd1 vssd1 vccd1 vccd1 net1517 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06184_ _01423_ vssd1 vssd1 vccd1 vccd1 top.a1.nextHex\[7\] sky130_fd_sc_hd__inv_2
XFILLER_0_111_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_170_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold412 top.DUT.register\[20\]\[7\] vssd1 vssd1 vccd1 vccd1 net1528 sky130_fd_sc_hd__dlygate4sd3_1
Xhold423 top.DUT.register\[15\]\[4\] vssd1 vssd1 vccd1 vccd1 net1539 sky130_fd_sc_hd__dlygate4sd3_1
Xhold434 top.DUT.register\[13\]\[31\] vssd1 vssd1 vccd1 vccd1 net1550 sky130_fd_sc_hd__dlygate4sd3_1
Xhold445 top.DUT.register\[8\]\[19\] vssd1 vssd1 vccd1 vccd1 net1561 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12491__RESET_B net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold456 top.ramaddr\[2\] vssd1 vssd1 vccd1 vccd1 net1572 sky130_fd_sc_hd__dlygate4sd3_1
Xhold467 top.DUT.register\[23\]\[9\] vssd1 vssd1 vccd1 vccd1 net1583 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09517__A top.pc\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold478 top.DUT.register\[2\]\[3\] vssd1 vssd1 vccd1 vccd1 net1594 sky130_fd_sc_hd__dlygate4sd3_1
X_09943_ top.a1.instruction\[7\] top.a1.instruction\[8\] _04708_ vssd1 vssd1 vccd1
+ vccd1 _04947_ sky130_fd_sc_hd__and3b_2
Xhold489 top.DUT.register\[13\]\[22\] vssd1 vssd1 vccd1 vccd1 net1605 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout903 top.i_ready vssd1 vssd1 vccd1 vccd1 net903 sky130_fd_sc_hd__clkbuf_4
Xfanout914 net915 vssd1 vssd1 vccd1 vccd1 net914 sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_39_Right_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout925 net935 vssd1 vssd1 vccd1 vccd1 net925 sky130_fd_sc_hd__buf_2
XFILLER_0_110_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout399_A net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout936 net939 vssd1 vssd1 vccd1 vccd1 net936 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09715__A1 _03514_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10162__S net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09874_ _03929_ net406 net491 _04884_ vssd1 vssd1 vccd1 vccd1 _04885_ sky130_fd_sc_hd__o211a_1
Xfanout947 net952 vssd1 vssd1 vccd1 vccd1 net947 sky130_fd_sc_hd__buf_2
Xfanout958 net966 vssd1 vssd1 vccd1 vccd1 net958 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07726__B1 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1101 top.DUT.register\[8\]\[30\] vssd1 vssd1 vccd1 vccd1 net2217 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09951__S net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout969 net970 vssd1 vssd1 vccd1 vccd1 net969 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_146_2630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1112 top.DUT.register\[22\]\[28\] vssd1 vssd1 vccd1 vccd1 net2228 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_146_2641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08825_ _03898_ _03937_ net290 vssd1 vssd1 vccd1 vccd1 _03938_ sky130_fd_sc_hd__mux2_1
Xhold1123 top.DUT.register\[4\]\[4\] vssd1 vssd1 vccd1 vccd1 net2239 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1134 top.DUT.register\[26\]\[15\] vssd1 vssd1 vccd1 vccd1 net2250 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1145 top.DUT.register\[25\]\[25\] vssd1 vssd1 vccd1 vccd1 net2261 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout566_A _01528_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11782__A top.a1.dataIn\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1156 top.DUT.register\[14\]\[2\] vssd1 vssd1 vccd1 vccd1 net2272 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_197_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1167 top.DUT.register\[14\]\[17\] vssd1 vssd1 vccd1 vccd1 net2283 sky130_fd_sc_hd__dlygate4sd3_1
X_08756_ _02136_ _03871_ vssd1 vssd1 vccd1 vccd1 _03872_ sky130_fd_sc_hd__xnor2_1
Xhold1178 top.DUT.register\[21\]\[3\] vssd1 vssd1 vccd1 vccd1 net2294 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1189 top.DUT.register\[29\]\[4\] vssd1 vssd1 vccd1 vccd1 net2305 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09252__A _02329_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11286__B1 _05149_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07707_ top.DUT.register\[2\]\[4\] net561 net548 top.DUT.register\[18\]\[4\] vssd1
+ vssd1 vccd1 vccd1 _02846_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout733_A _01627_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08687_ net497 _03790_ _03803_ _03806_ vssd1 vssd1 vccd1 vccd1 _03807_ sky130_fd_sc_hd__o211ai_4
XANTENNA_fanout354_X net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1096_X net1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07638_ top.a1.instruction\[26\] net805 _02775_ _02776_ vssd1 vssd1 vccd1 vccd1 _02777_
+ sky130_fd_sc_hd__a22oi_4
XFILLER_0_193_711 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_48_Right_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_165_424 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout521_X net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07569_ top.DUT.register\[23\]\[6\] net571 net543 top.DUT.register\[16\]\[6\] _02707_
+ vssd1 vssd1 vccd1 vccd1 _02708_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout900_A net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout619_X net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_192_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09308_ _02399_ _02408_ _04370_ vssd1 vssd1 vccd1 vccd1 _04372_ sky130_fd_sc_hd__o21ai_1
X_10580_ net1458 net216 net350 vssd1 vssd1 vccd1 vccd1 _00746_ sky130_fd_sc_hd__mux2_1
XANTENNA__07257__A2 net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12687__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12579__RESET_B net1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09239_ _04303_ _04306_ vssd1 vssd1 vccd1 vccd1 _04307_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10337__S net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12118__A top.a1.dataIn\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_9__f_clk_A clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_354 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12250_ _06080_ _06081_ vssd1 vssd1 vccd1 vccd1 _01325_ sky130_fd_sc_hd__nor2_1
XANTENNA__07009__A2 net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08206__A1 net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12508__RESET_B net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout890_X net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout988_X net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11201_ net845 _05012_ _05024_ vssd1 vssd1 vccd1 vccd1 _05107_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_170_2992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12181_ net1281 net846 net796 _05879_ vssd1 vssd1 vccd1 vccd1 _01289_ sky130_fd_sc_hd__a22o_1
XFILLER_0_31_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_57_Right_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07965__B1 net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11132_ net907 net1489 net862 _05071_ vssd1 vssd1 vccd1 vccd1 _01217_ sky130_fd_sc_hd__a31o_1
XANTENNA__06403__X _01542_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold990 top.DUT.register\[27\]\[21\] vssd1 vssd1 vccd1 vccd1 net2106 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11063_ net78 net870 net834 net1143 vssd1 vssd1 vccd1 vccd1 _01174_ sky130_fd_sc_hd__a22o_1
XANTENNA__10072__S net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10014_ net1691 net147 net619 vssd1 vssd1 vccd1 vccd1 _00217_ sky130_fd_sc_hd__mux2_1
XFILLER_0_204_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10800__S net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_203_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_86_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11965_ _05814_ _05821_ _05819_ vssd1 vssd1 vccd1 vccd1 _05848_ sky130_fd_sc_hd__o21a_1
XFILLER_0_58_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_66_Right_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13704_ clknet_leaf_96_clk _01275_ net984 vssd1 vssd1 vccd1 vccd1 top.a1.row2\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_10916_ net2234 net157 net481 vssd1 vssd1 vccd1 vccd1 _01077_ sky130_fd_sc_hd__mux2_1
XANTENNA__07496__A2 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11896_ _05770_ _05773_ _05774_ _05775_ _05767_ vssd1 vssd1 vccd1 vccd1 _05779_ sky130_fd_sc_hd__o41a_2
XFILLER_0_86_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_184_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13635_ clknet_leaf_72_clk _01222_ net1080 vssd1 vssd1 vccd1 vccd1 net63 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_132_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10847_ net1740 net177 net475 vssd1 vssd1 vccd1 vccd1 _01008_ sky130_fd_sc_hd__mux2_1
XFILLER_0_144_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08445__A1 _02498_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13566_ clknet_leaf_105_clk _01153_ net969 vssd1 vssd1 vccd1 vccd1 top.ramload\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_171_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_444 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10778_ net1348 net203 net484 vssd1 vssd1 vccd1 vccd1 _00939_ sky130_fd_sc_hd__mux2_1
XANTENNA__09101__S _04142_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12517_ clknet_leaf_87_clk _00109_ net1083 vssd1 vssd1 vccd1 vccd1 top.pc\[29\] sky130_fd_sc_hd__dfstp_2
XANTENNA__10247__S net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13497_ clknet_leaf_15_clk _01089_ net961 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[31\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12448_ clknet_leaf_72_clk _00044_ net1080 vssd1 vssd1 vccd1 vccd1 top.ramaddr\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_75_Right_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11289__D top.lcd.nextState\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10193__D net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_2139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_1894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12379_ clknet_leaf_108_clk top.ru.next_FetchedData\[23\] net975 vssd1 vssd1 vccd1
+ vccd1 top.a1.dataIn\[23\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_1_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07420__A2 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06940_ top.DUT.register\[10\]\[21\] net773 net740 top.DUT.register\[12\]\[21\] vssd1
+ vssd1 vccd1 vccd1 _02079_ sky130_fd_sc_hd__a22o_1
XFILLER_0_157_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07708__B1 net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09173__A2 _02849_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06871_ top.DUT.register\[20\]\[18\] net565 net525 top.DUT.register\[11\]\[18\] vssd1
+ vssd1 vccd1 vccd1 _02010_ sky130_fd_sc_hd__a22o_1
XFILLER_0_207_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_206_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_128_2360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08610_ net308 _03649_ vssd1 vssd1 vccd1 vccd1 _03733_ sky130_fd_sc_hd__or2_1
XFILLER_0_179_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_2371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10710__S net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09590_ top.pc\[30\] _04620_ vssd1 vssd1 vccd1 vccd1 _04637_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_50_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_84_Right_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_179_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08541_ _02474_ _03659_ vssd1 vssd1 vccd1 vccd1 _03667_ sky130_fd_sc_hd__or2_1
XFILLER_0_77_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_141_2560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08472_ _03551_ _03600_ net292 vssd1 vssd1 vccd1 vccd1 _03601_ sky130_fd_sc_hd__mux2_1
XANTENNA__08684__A1 _02049_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07487__A2 net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07423_ top.DUT.register\[20\]\[9\] net663 net770 top.DUT.register\[10\]\[9\] _02561_
+ vssd1 vssd1 vccd1 vccd1 _02562_ sky130_fd_sc_hd__a221o_1
XFILLER_0_147_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout147_A _04724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_175_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07354_ top.DUT.register\[7\]\[8\] net516 net444 top.DUT.register\[1\]\[8\] _02492_
+ vssd1 vssd1 vccd1 vccd1 _02493_ sky130_fd_sc_hd__a221o_1
XANTENNA__07239__A2 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_287 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06305_ _01459_ _01460_ vssd1 vssd1 vccd1 vccd1 _01461_ sky130_fd_sc_hd__nor2_1
XFILLER_0_33_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_21_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10157__S net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07285_ top.DUT.register\[10\]\[13\] net772 net736 top.DUT.register\[16\]\[13\] vssd1
+ vssd1 vccd1 vccd1 _02424_ sky130_fd_sc_hd__a22o_1
XFILLER_0_127_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout314_A _02924_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09024_ _01962_ _02048_ _02090_ _02265_ vssd1 vssd1 vccd1 vccd1 _04099_ sky130_fd_sc_hd__nand4_1
XPHY_EDGE_ROW_93_Right_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06236_ top.ramload\[30\] net859 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedInstr\[30\]
+ sky130_fd_sc_hd__and2_1
XANTENNA__09946__S net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_198_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_57_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold220 top.DUT.register\[31\]\[18\] vssd1 vssd1 vccd1 vccd1 net1336 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11777__A top.a1.dataIn\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06167_ top.a1.state\[1\] top.a1.state\[2\] top.a1.state\[0\] vssd1 vssd1 vccd1 vccd1
+ _01409_ sky130_fd_sc_hd__or3b_2
XFILLER_0_198_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold231 top.DUT.register\[4\]\[16\] vssd1 vssd1 vccd1 vccd1 net1347 sky130_fd_sc_hd__dlygate4sd3_1
Xhold242 top.DUT.register\[30\]\[3\] vssd1 vssd1 vccd1 vccd1 net1358 sky130_fd_sc_hd__dlygate4sd3_1
Xhold253 top.DUT.register\[28\]\[8\] vssd1 vssd1 vccd1 vccd1 net1369 sky130_fd_sc_hd__dlygate4sd3_1
Xhold264 top.DUT.register\[5\]\[25\] vssd1 vssd1 vccd1 vccd1 net1380 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13335__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07411__A2 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08151__A _02944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold275 top.DUT.register\[6\]\[25\] vssd1 vssd1 vccd1 vccd1 net1391 sky130_fd_sc_hd__dlygate4sd3_1
Xhold286 top.DUT.register\[15\]\[19\] vssd1 vssd1 vccd1 vccd1 net1402 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_582 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout700 _01643_ vssd1 vssd1 vccd1 vccd1 net700 sky130_fd_sc_hd__clkbuf_8
Xhold297 top.DUT.register\[26\]\[19\] vssd1 vssd1 vccd1 vccd1 net1413 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_70_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout711 _01638_ vssd1 vssd1 vccd1 vccd1 net711 sky130_fd_sc_hd__buf_4
XANTENNA__13807__RESET_B net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout722 _01630_ vssd1 vssd1 vccd1 vccd1 net722 sky130_fd_sc_hd__clkbuf_8
X_09926_ top.pc\[30\] _04628_ vssd1 vssd1 vccd1 vccd1 _04932_ sky130_fd_sc_hd__nor2_1
Xfanout733 _01627_ vssd1 vssd1 vccd1 vccd1 net733 sky130_fd_sc_hd__clkbuf_4
Xfanout744 _01623_ vssd1 vssd1 vccd1 vccd1 net744 sky130_fd_sc_hd__clkbuf_8
Xfanout755 _01620_ vssd1 vssd1 vccd1 vccd1 net755 sky130_fd_sc_hd__clkbuf_4
Xfanout766 net769 vssd1 vssd1 vccd1 vccd1 net766 sky130_fd_sc_hd__clkbuf_8
Xfanout777 _01608_ vssd1 vssd1 vccd1 vccd1 net777 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout850_A net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09857_ top.pc\[24\] _04543_ vssd1 vssd1 vccd1 vccd1 _04869_ sky130_fd_sc_hd__xor2_1
Xfanout788 _01591_ vssd1 vssd1 vccd1 vccd1 net788 sky130_fd_sc_hd__buf_2
Xfanout799 _04150_ vssd1 vssd1 vccd1 vccd1 net799 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout569_X net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13460__RESET_B net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08808_ net284 net429 vssd1 vssd1 vccd1 vccd1 _03922_ sky130_fd_sc_hd__nand2_1
XANTENNA__09613__D_N top.a1.halfData\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10620__S net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09788_ top.pc\[17\] _04438_ vssd1 vssd1 vccd1 vccd1 _04807_ sky130_fd_sc_hd__nor2_1
X_08739_ _03206_ _03210_ vssd1 vssd1 vccd1 vccd1 _03856_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_1_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout736_X net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_368 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11750_ _05603_ _05619_ vssd1 vssd1 vccd1 vccd1 _05633_ sky130_fd_sc_hd__nor2_1
XANTENNA__07478__A2 net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09872__B1 _04151_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_159_2832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06686__B1 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10701_ net1491 net253 net334 vssd1 vssd1 vccd1 vccd1 _00862_ sky130_fd_sc_hd__mux2_1
XFILLER_0_165_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11681_ _05530_ _05549_ _05533_ vssd1 vssd1 vccd1 vccd1 _05564_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout903_X net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13420_ clknet_leaf_49_clk _01012_ net1060 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[28\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_181_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10632_ net260 net1624 net344 vssd1 vssd1 vccd1 vccd1 _00796_ sky130_fd_sc_hd__mux2_1
XANTENNA__08427__B2 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10067__S net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10563_ net1777 net146 net353 vssd1 vssd1 vccd1 vccd1 _00729_ sky130_fd_sc_hd__mux2_1
X_13351_ clknet_leaf_8_clk _00943_ net947 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[26\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_118_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_180_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12302_ top.pad.button_control.r_counter\[0\] net790 vssd1 vssd1 vccd1 vccd1 _01352_
+ sky130_fd_sc_hd__and2b_1
XANTENNA__09856__S net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13282_ clknet_leaf_25_clk _00874_ net1012 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[24\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_10494_ net1623 net140 net363 vssd1 vssd1 vccd1 vccd1 _00664_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_184 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12233_ net2167 _06069_ net978 vssd1 vssd1 vccd1 vccd1 _06071_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_121_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12164_ _06036_ _06043_ vssd1 vssd1 vccd1 vccd1 _06046_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09157__A _02808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08061__A _01897_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07402__A2 net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11115_ net48 net865 vssd1 vssd1 vccd1 vccd1 _05063_ sky130_fd_sc_hd__and2_1
XANTENNA__06610__B1 net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12095_ _05960_ _05968_ _05973_ _05977_ vssd1 vssd1 vccd1 vccd1 _05978_ sky130_fd_sc_hd__a22o_2
XTAP_TAPCELL_ROW_207_3545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11046_ wb.curr_state\[1\] net905 wb.curr_state\[2\] vssd1 vssd1 vccd1 vccd1 _05045_
+ sky130_fd_sc_hd__and3b_2
XTAP_TAPCELL_ROW_207_3556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07166__A1 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_204_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_188_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_207_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12997_ clknet_leaf_33_clk _00589_ net1046 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[15\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_143_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_379 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11948_ _05812_ _05829_ vssd1 vssd1 vccd1 vccd1 _05831_ sky130_fd_sc_hd__xnor2_2
XANTENNA__09042__D net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_96_Left_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_123_2290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06677__B1 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10473__A1 net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_184_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13208__CLK clknet_leaf_128_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11879_ _05744_ _05761_ vssd1 vssd1 vccd1 vccd1 _05762_ sky130_fd_sc_hd__or2_1
XFILLER_0_172_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_157_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_591 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13618_ clknet_leaf_75_clk _01205_ net1079 vssd1 vssd1 vccd1 vccd1 net44 sky130_fd_sc_hd__dfrtp_1
XANTENNA__06429__B1 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_1934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13549_ clknet_leaf_104_clk _01136_ net973 vssd1 vssd1 vccd1 vccd1 top.ramload\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_201_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07070_ top.DUT.register\[14\]\[22\] net731 net726 top.DUT.register\[18\]\[22\] vssd1
+ vssd1 vccd1 vccd1 _02209_ sky130_fd_sc_hd__a22o_1
XANTENNA__07641__A2 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10705__S net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12192__S _06049_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09394__A2 _02679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_379 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_168_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07972_ _03104_ _03106_ _03108_ _03110_ vssd1 vssd1 vccd1 vccd1 _03111_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_52_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09711_ net1452 net251 net631 vssd1 vssd1 vccd1 vccd1 _00126_ sky130_fd_sc_hd__mux2_1
X_06923_ top.DUT.register\[25\]\[21\] net457 net525 top.DUT.register\[11\]\[21\] vssd1
+ vssd1 vccd1 vccd1 _02062_ sky130_fd_sc_hd__a22o_1
X_09642_ top.pad.keyCode\[4\] top.pad.keyCode\[5\] top.pad.keyCode\[6\] top.pad.keyCode\[7\]
+ vssd1 vssd1 vccd1 vccd1 _04684_ sky130_fd_sc_hd__or4b_2
XANTENNA__10440__S net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06854_ top.DUT.register\[15\]\[19\] net709 net701 top.DUT.register\[31\]\[19\] vssd1
+ vssd1 vccd1 vccd1 _01993_ sky130_fd_sc_hd__a22o_1
XFILLER_0_179_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06785_ top.DUT.register\[26\]\[17\] net527 net524 top.DUT.register\[11\]\[17\] vssd1
+ vssd1 vccd1 vccd1 _01924_ sky130_fd_sc_hd__a22o_1
X_09573_ _01678_ _04620_ vssd1 vssd1 vccd1 vccd1 _04621_ sky130_fd_sc_hd__xor2_1
XANTENNA_fanout264_A _04729_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08524_ net309 _03553_ _03650_ vssd1 vssd1 vccd1 vccd1 _03651_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_26_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06668__B1 net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08455_ _03347_ _03533_ _03584_ vssd1 vssd1 vccd1 vccd1 _03585_ sky130_fd_sc_hd__a21o_1
XFILLER_0_148_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout431_A net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout529_A net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_172_3029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07406_ top.a1.instruction\[30\] net789 net410 vssd1 vssd1 vccd1 vccd1 _02545_ sky130_fd_sc_hd__a21o_1
XFILLER_0_9_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08386_ _02678_ _02704_ vssd1 vssd1 vccd1 vccd1 _03518_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_63_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire408 net409 vssd1 vssd1 vccd1 vccd1 net408 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_190_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07337_ _02474_ _02475_ vssd1 vssd1 vccd1 vccd1 _02476_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_154_2751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_154_2762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07268_ top.DUT.register\[13\]\[13\] net465 net449 top.DUT.register\[21\]\[13\] _02406_
+ vssd1 vssd1 vccd1 vccd1 _02407_ sky130_fd_sc_hd__a221o_1
XFILLER_0_143_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07632__A2 net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout898_A net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09007_ _03443_ _03473_ _03508_ _03532_ vssd1 vssd1 vccd1 vccd1 _04082_ sky130_fd_sc_hd__or4b_1
X_06219_ net2312 net856 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedInstr\[13\] sky130_fd_sc_hd__and2_1
XFILLER_0_5_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06840__B1 net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10615__S net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07199_ _01480_ _02336_ vssd1 vssd1 vccd1 vccd1 _02338_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_187_3250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_491 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_699 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout530 _01550_ vssd1 vssd1 vccd1 vccd1 net530 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_6_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09137__A2 _02952_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout541 _01540_ vssd1 vssd1 vccd1 vccd1 net541 sky130_fd_sc_hd__clkbuf_8
X_09909_ net1598 net158 net634 vssd1 vssd1 vccd1 vccd1 _00149_ sky130_fd_sc_hd__mux2_1
Xfanout552 _01535_ vssd1 vssd1 vccd1 vccd1 net552 sky130_fd_sc_hd__clkbuf_4
Xfanout563 _01528_ vssd1 vssd1 vccd1 vccd1 net563 sky130_fd_sc_hd__buf_6
XANTENNA_fanout853_X net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout574 _01519_ vssd1 vssd1 vccd1 vccd1 net574 sky130_fd_sc_hd__buf_4
XANTENNA__08345__B1 net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout585 _01513_ vssd1 vssd1 vccd1 vccd1 net585 sky130_fd_sc_hd__clkbuf_8
XANTENNA__10350__S net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12920_ clknet_leaf_128_clk _00512_ net911 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[13\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout596 _04966_ vssd1 vssd1 vccd1 vccd1 net596 sky130_fd_sc_hd__buf_6
XANTENNA__07699__A2 net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12851_ clknet_leaf_123_clk _00443_ net926 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[11\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_202_3475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11802_ _05632_ _05684_ vssd1 vssd1 vccd1 vccd1 _05685_ sky130_fd_sc_hd__and2b_1
XFILLER_0_198_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12782_ clknet_leaf_41_clk _00374_ net1047 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[8\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_96_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_200_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06659__B1 net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11733_ _05579_ _05612_ vssd1 vssd1 vccd1 vccd1 _05616_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_83_314 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11664_ _05487_ _05518_ vssd1 vssd1 vccd1 vccd1 _05547_ sky130_fd_sc_hd__xor2_1
XANTENNA__07871__A2 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13500__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13403_ clknet_leaf_124_clk _00995_ net925 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[28\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_10615_ net184 net2256 net348 vssd1 vssd1 vccd1 vccd1 _00780_ sky130_fd_sc_hd__mux2_1
X_11595_ _05462_ net239 net234 _05476_ vssd1 vssd1 vccd1 vccd1 _05478_ sky130_fd_sc_hd__a22oi_2
X_13334_ clknet_leaf_4_clk _00926_ net938 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[26\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07623__A2 net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10546_ net1516 net223 net356 vssd1 vssd1 vccd1 vccd1 _00713_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_611 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06831__B1 net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10525__S net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13265_ clknet_leaf_115_clk _00857_ net966 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[24\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_10477_ net1922 net198 net362 vssd1 vssd1 vccd1 vccd1 _00647_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_94_1853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12216_ _06059_ _06060_ net980 vssd1 vssd1 vccd1 vccd1 _01312_ sky130_fd_sc_hd__o21a_1
X_13196_ clknet_leaf_47_clk _00788_ net1069 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[21\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_209_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11183__A2 net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12147_ _06022_ _06026_ vssd1 vssd1 vccd1 vccd1 _06030_ sky130_fd_sc_hd__xnor2_1
X_12078_ _05931_ _05952_ _05956_ vssd1 vssd1 vccd1 vccd1 _05961_ sky130_fd_sc_hd__or3_1
XANTENNA__09533__C1 net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10260__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11029_ net8 net838 net816 net1204 vssd1 vssd1 vccd1 vccd1 _01141_ sky130_fd_sc_hd__o22a_1
XANTENNA__09334__B _04386_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06898__B1 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09039__D_N _01659_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13030__CLK clknet_leaf_40_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06570_ top.DUT.register\[14\]\[28\] net585 net446 top.DUT.register\[1\]\[28\] vssd1
+ vssd1 vccd1 vccd1 _01709_ sky130_fd_sc_hd__a22o_1
XFILLER_0_177_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_686 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08240_ _03376_ vssd1 vssd1 vccd1 vccd1 _03377_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_157_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07862__A2 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_103_1993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08171_ _03307_ _03308_ vssd1 vssd1 vccd1 vccd1 _03309_ sky130_fd_sc_hd__nand2_1
XFILLER_0_103_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07122_ net807 net412 net437 vssd1 vssd1 vccd1 vccd1 _02261_ sky130_fd_sc_hd__o21a_1
XFILLER_0_12_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07075__B1 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08811__A1 _03260_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_2481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_136_2492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06822__B1 net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07053_ top.DUT.register\[2\]\[22\] net560 net460 top.DUT.register\[17\]\[22\] _02191_
+ vssd1 vssd1 vccd1 vccd1 _02192_ sky130_fd_sc_hd__a221o_1
XANTENNA__10435__S net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput100 net100 vssd1 vssd1 vccd1 vccd1 DAT_O[5] sky130_fd_sc_hd__buf_2
XANTENNA__09509__B _04560_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput111 net111 vssd1 vssd1 vccd1 vccd1 gpio_out[0] sky130_fd_sc_hd__buf_2
XFILLER_0_11_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput122 net122 vssd1 vssd1 vccd1 vccd1 gpio_out[7] sky130_fd_sc_hd__buf_2
XFILLER_0_2_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1019_A net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09525__A net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07955_ _01810_ _01830_ _03093_ vssd1 vssd1 vccd1 vccd1 _03094_ sky130_fd_sc_hd__a21oi_1
XANTENNA__06501__X _01640_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout381_A net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_182_3180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout479_A _04964_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06906_ _02035_ _02044_ vssd1 vssd1 vccd1 vccd1 _02045_ sky130_fd_sc_hd__nor2_1
XANTENNA__10170__S net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07886_ top.DUT.register\[13\]\[1\] net465 net458 top.DUT.register\[25\]\[1\] _03024_
+ vssd1 vssd1 vccd1 vccd1 _03025_ sky130_fd_sc_hd__a221o_1
XANTENNA__09812__X _04829_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06889__B1 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09625_ _04656_ _04669_ vssd1 vssd1 vccd1 vccd1 _04670_ sky130_fd_sc_hd__nor2_1
X_06837_ top.DUT.register\[6\]\[19\] net570 net517 top.DUT.register\[7\]\[19\] vssd1
+ vssd1 vccd1 vccd1 _01976_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout646_A _01613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09556_ top.a1.instruction\[28\] net822 net422 vssd1 vssd1 vccd1 vccd1 _04605_ sky130_fd_sc_hd__a21o_2
X_06768_ top.DUT.register\[16\]\[24\] net735 net700 top.DUT.register\[31\]\[24\] vssd1
+ vssd1 vccd1 vccd1 _01907_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_65_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08507_ _03263_ _03623_ _03633_ _03634_ vssd1 vssd1 vccd1 vccd1 _03635_ sky130_fd_sc_hd__a211o_1
XFILLER_0_78_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06699_ top.DUT.register\[13\]\[25\] net463 net531 top.DUT.register\[12\]\[25\] _01837_
+ vssd1 vssd1 vccd1 vccd1 _01838_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout813_A net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09487_ _04538_ _04539_ vssd1 vssd1 vccd1 vccd1 _04540_ sky130_fd_sc_hd__and2b_1
XANTENNA_fanout434_X net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08438_ net423 _03550_ _03568_ _03334_ _03564_ vssd1 vssd1 vccd1 vccd1 _03569_ sky130_fd_sc_hd__a221o_2
XFILLER_0_18_230 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07853__A2 net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08369_ _03230_ _03234_ vssd1 vssd1 vccd1 vccd1 _03502_ sky130_fd_sc_hd__nand2_1
XFILLER_0_92_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout601_X net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_594 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10400_ net1625 net259 net370 vssd1 vssd1 vccd1 vccd1 _00572_ sky130_fd_sc_hd__mux2_1
X_11380_ _05230_ _05261_ vssd1 vssd1 vccd1 vccd1 _05263_ sky130_fd_sc_hd__xnor2_2
XANTENNA__07605__A2 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10331_ net2091 net266 net377 vssd1 vssd1 vccd1 vccd1 _00507_ sky130_fd_sc_hd__mux2_1
XANTENNA__06813__B1 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10345__S net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_491 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10262_ _04155_ _04958_ net399 vssd1 vssd1 vccd1 vccd1 _04978_ sky130_fd_sc_hd__and3_4
X_13050_ clknet_leaf_4_clk _00642_ net936 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[17\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_76_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12001_ _05861_ _05883_ vssd1 vssd1 vccd1 vccd1 _05884_ sky130_fd_sc_hd__xor2_1
X_10193_ net482 net478 net474 net593 vssd1 vssd1 vccd1 vccd1 _04973_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_167_2953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_204_3504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout360 _04987_ vssd1 vssd1 vccd1 vccd1 net360 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_205_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout371 net372 vssd1 vssd1 vccd1 vccd1 net371 sky130_fd_sc_hd__buf_2
XANTENNA__06592__A2 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10080__S net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout382 net384 vssd1 vssd1 vccd1 vccd1 net382 sky130_fd_sc_hd__buf_6
Xfanout393 net396 vssd1 vssd1 vccd1 vccd1 net393 sky130_fd_sc_hd__buf_6
XANTENNA__09154__B _02857_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12903_ clknet_leaf_8_clk _00495_ net945 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[12\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12513__SET_B net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12834_ clknet_leaf_10_clk _00426_ net949 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[10\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_33_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12765_ clknet_leaf_119_clk _00357_ net930 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[8\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09294__A1 net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_173_319 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_204_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11716_ _05560_ _05593_ vssd1 vssd1 vccd1 vccd1 _05599_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_83_133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07844__A2 net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_667 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12696_ clknet_leaf_125_clk _00288_ net923 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[6\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_224 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09046__A1 net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11647_ _05522_ _05528_ vssd1 vssd1 vccd1 vccd1 _05530_ sky130_fd_sc_hd__nand2_1
Xinput13 DAT_I[1] vssd1 vssd1 vccd1 vccd1 net13 sky130_fd_sc_hd__buf_1
XFILLER_0_114_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput24 DAT_I[2] vssd1 vssd1 vccd1 vccd1 net24 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07057__B1 net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput35 gpio_in[15] vssd1 vssd1 vccd1 vccd1 net35 sky130_fd_sc_hd__clkbuf_1
X_11578_ _05460_ vssd1 vssd1 vccd1 vccd1 _05461_ sky130_fd_sc_hd__inv_2
XFILLER_0_52_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13317_ clknet_leaf_33_clk _00909_ net1043 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[25\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06804__B1 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold808 top.DUT.register\[12\]\[23\] vssd1 vssd1 vccd1 vccd1 net1924 sky130_fd_sc_hd__dlygate4sd3_1
X_10529_ _04712_ _04949_ net400 vssd1 vssd1 vccd1 vccd1 _04989_ sky130_fd_sc_hd__and3_4
XANTENNA__10255__S net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold819 top.DUT.register\[30\]\[23\] vssd1 vssd1 vccd1 vccd1 net1935 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_172_Right_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13248_ clknet_leaf_79_clk _00840_ net1073 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[23\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_149_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11156__A2 net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_199_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13179_ clknet_leaf_120_clk _00771_ net931 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[21\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08309__B1 _03437_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07740_ _02858_ _02877_ net823 vssd1 vssd1 vccd1 vccd1 _02879_ sky130_fd_sc_hd__mux2_1
XFILLER_0_165_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_74_clk_A clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07671_ top.DUT.register\[13\]\[4\] net775 net708 top.DUT.register\[15\]\[4\] vssd1
+ vssd1 vccd1 vccd1 _02810_ sky130_fd_sc_hd__a22o_1
X_09410_ _04466_ _04467_ vssd1 vssd1 vccd1 vccd1 _04468_ sky130_fd_sc_hd__xnor2_1
X_06622_ top.DUT.register\[7\]\[27\] net518 net514 top.DUT.register\[24\]\[27\] vssd1
+ vssd1 vccd1 vccd1 _01761_ sky130_fd_sc_hd__a22o_1
XFILLER_0_204_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_177_647 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09080__A top.a1.instruction\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06553_ top.DUT.register\[23\]\[29\] net673 net708 top.DUT.register\[15\]\[29\] _01691_
+ vssd1 vssd1 vccd1 vccd1 _01692_ sky130_fd_sc_hd__a221o_1
X_09341_ _01577_ _02805_ _04335_ _04402_ vssd1 vssd1 vccd1 vccd1 _04403_ sky130_fd_sc_hd__o22a_2
XPHY_EDGE_ROW_188_Left_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_36_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_89_clk_A clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07296__B1 net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11092__A1 net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06484_ net787 _01611_ _01618_ vssd1 vssd1 vccd1 vccd1 _01623_ sky130_fd_sc_hd__and3_4
X_09272_ _02286_ _04337_ vssd1 vssd1 vccd1 vccd1 _04338_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_138_2510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_2521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08223_ net292 _03235_ vssd1 vssd1 vccd1 vccd1 _03360_ sky130_fd_sc_hd__or2_1
XFILLER_0_7_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_60_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_60_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10954__A net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_380 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_659 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07048__B1 net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08154_ _02678_ _02498_ net331 vssd1 vssd1 vccd1 vccd1 _03292_ sky130_fd_sc_hd__mux2_1
XFILLER_0_160_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_12_clk_A clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_396 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_151_2710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_350 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_99_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_160_558 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07105_ top.DUT.register\[23\]\[16\] net672 net779 top.DUT.register\[25\]\[16\] _02243_
+ vssd1 vssd1 vccd1 vccd1 _02244_ sky130_fd_sc_hd__a221o_1
X_08085_ _02944_ net330 vssd1 vssd1 vccd1 vccd1 _03224_ sky130_fd_sc_hd__or2_1
XANTENNA__10165__S net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07036_ _02167_ _02174_ vssd1 vssd1 vccd1 vccd1 _02175_ sky130_fd_sc_hd__nor2_2
XANTENNA__09954__S net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13233__RESET_B net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08711__X _03830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout596_A _04966_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_27_clk_A clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_180_3139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08987_ _04014_ _04032_ _04061_ vssd1 vssd1 vccd1 vccd1 _04062_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout763_A net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06574__A2 net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout384_X net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_149_2683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_199_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07938_ _01940_ _01961_ vssd1 vssd1 vccd1 vccd1 _03077_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_162_2872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout551_X net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07869_ top.DUT.register\[9\]\[1\] net763 net736 top.DUT.register\[16\]\[1\] vssd1
+ vssd1 vccd1 vccd1 _03008_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_162_2883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout649_X net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09608_ net138 _04652_ net902 vssd1 vssd1 vccd1 vccd1 _04654_ sky130_fd_sc_hd__o21a_1
XFILLER_0_167_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10880_ net175 net2190 net596 vssd1 vssd1 vccd1 vccd1 _01041_ sky130_fd_sc_hd__mux2_1
XFILLER_0_210_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09539_ top.pc\[27\] _04567_ vssd1 vssd1 vccd1 vccd1 _04589_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_195_3371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12550_ clknet_leaf_38_clk _00142_ net1054 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[1\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07287__B1 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07826__A2 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_176_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_182_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11501_ _05315_ _05345_ vssd1 vssd1 vccd1 vccd1 _05384_ sky130_fd_sc_hd__nand2_1
XFILLER_0_65_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12481_ clknet_leaf_66_clk _00076_ net1094 vssd1 vssd1 vccd1 vccd1 top.ramstore\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_136_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_374 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11432_ _05273_ _05307_ vssd1 vssd1 vccd1 vccd1 _05315_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_78_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_190_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10075__S net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11363_ _05237_ _05245_ vssd1 vssd1 vccd1 vccd1 _05246_ sky130_fd_sc_hd__nand2_1
XANTENNA__08251__A2 net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13102_ clknet_leaf_40_clk _00694_ net1055 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[18\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_10314_ net203 net1981 net382 vssd1 vssd1 vccd1 vccd1 _00491_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_91_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11294_ net1179 net814 _05183_ net1003 vssd1 vssd1 vccd1 vccd1 _01267_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_210_3596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13033_ clknet_leaf_52_clk _00625_ net1038 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[16\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10803__S net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10245_ net190 net1814 net389 vssd1 vssd1 vccd1 vccd1 _00424_ sky130_fd_sc_hd__mux2_1
XANTENNA__08003__A2 _03141_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10176_ net2217 net151 net605 vssd1 vssd1 vccd1 vccd1 _00375_ sky130_fd_sc_hd__mux2_1
XANTENNA__06565__A2 net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_201_Left_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout190 net191 vssd1 vssd1 vccd1 vccd1 net190 sky130_fd_sc_hd__buf_2
XFILLER_0_135_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_89_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07514__A1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11310__A2 _05130_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkload5_A clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09612__B net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12817_ clknet_leaf_116_clk _00409_ net958 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[10\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13797_ clknet_leaf_68_clk _01366_ vssd1 vssd1 vccd1 vccd1 top.pad.button_control.r_counter\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_186_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07278__B1 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12748_ clknet_leaf_64_clk _00340_ net1093 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[7\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07817__A2 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_210_Left_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_139_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_68 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_100_1941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_100_1952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08490__A2 net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12679_ clknet_leaf_7_clk _00271_ net944 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[5\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_154_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_136 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_42_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08244__A net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13099__CLK clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_133_2440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold605 top.DUT.register\[12\]\[1\] vssd1 vssd1 vccd1 vccd1 net1721 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold616 top.ramaddr\[24\] vssd1 vssd1 vccd1 vccd1 net1732 sky130_fd_sc_hd__dlygate4sd3_1
Xhold627 top.DUT.register\[2\]\[23\] vssd1 vssd1 vccd1 vccd1 net1743 sky130_fd_sc_hd__dlygate4sd3_1
Xhold638 top.DUT.register\[10\]\[6\] vssd1 vssd1 vccd1 vccd1 net1754 sky130_fd_sc_hd__dlygate4sd3_1
Xhold649 top.DUT.register\[27\]\[28\] vssd1 vssd1 vccd1 vccd1 net1765 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_150_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08910_ net308 _03938_ _04018_ net285 vssd1 vssd1 vccd1 vccd1 _04019_ sky130_fd_sc_hd__o211a_1
X_09890_ top.pc\[27\] _04590_ vssd1 vssd1 vccd1 vccd1 _04899_ sky130_fd_sc_hd__or2_1
XANTENNA__10713__S net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08250__Y _03387_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08841_ net1923 net831 net801 _03953_ vssd1 vssd1 vccd1 vccd1 _00044_ sky130_fd_sc_hd__a22o_1
XANTENNA__06556__A2 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08950__B1 _02748_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08772_ _02222_ _03864_ _03082_ vssd1 vssd1 vccd1 vccd1 _03888_ sky130_fd_sc_hd__a21oi_1
XANTENNA__06211__B net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07723_ top.DUT.register\[7\]\[3\] net660 net637 top.DUT.register\[6\]\[3\] _02861_
+ vssd1 vssd1 vccd1 vccd1 _02862_ sky130_fd_sc_hd__a221o_1
XANTENNA__11301__A2 net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_260 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07654_ top.DUT.register\[16\]\[5\] net734 net636 top.DUT.register\[6\]\[5\] _02792_
+ vssd1 vssd1 vccd1 vccd1 _02793_ sky130_fd_sc_hd__a221o_1
XANTENNA__09522__B _04560_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_189_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06605_ _01721_ _01742_ vssd1 vssd1 vccd1 vccd1 _01744_ sky130_fd_sc_hd__nand2_1
XANTENNA__09258__A1 net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07585_ _02723_ vssd1 vssd1 vccd1 vccd1 _02724_ sky130_fd_sc_hd__inv_2
XFILLER_0_192_403 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout344_A _04992_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1086_A net1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09324_ _02623_ _02632_ _04386_ vssd1 vssd1 vccd1 vccd1 _04387_ sky130_fd_sc_hd__o21ai_1
XANTENNA__09949__S net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06536_ top.DUT.register\[20\]\[29\] net565 net509 top.DUT.register\[4\]\[29\] vssd1
+ vssd1 vccd1 vccd1 _01675_ sky130_fd_sc_hd__a22o_1
XANTENNA__10955__Y _04998_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07610__X _02749_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09255_ _04303_ _04305_ _04304_ vssd1 vssd1 vccd1 vccd1 _04322_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout511_A _01559_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06467_ _01592_ _01594_ _01596_ vssd1 vssd1 vccd1 vccd1 _01606_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout132_X net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08481__A2 _03534_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout609_A _04956_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08206_ net436 net284 _03332_ _03343_ vssd1 vssd1 vccd1 vccd1 _03344_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_190_3290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09186_ top.pc\[6\] _02778_ vssd1 vssd1 vccd1 vccd1 _04257_ sky130_fd_sc_hd__and2_1
X_06398_ top.DUT.register\[3\]\[30\] net553 net548 top.DUT.register\[18\]\[30\] vssd1
+ vssd1 vccd1 vccd1 _01537_ sky130_fd_sc_hd__a22o_1
X_08137_ _03273_ _03274_ vssd1 vssd1 vccd1 vccd1 _03275_ sky130_fd_sc_hd__nand2_1
XFILLER_0_31_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08068_ _02111_ net327 vssd1 vssd1 vccd1 vccd1 _03207_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout880_A net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout599_X net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06795__A2 net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07019_ top.DUT.register\[2\]\[20\] net745 net725 top.DUT.register\[29\]\[20\] vssd1
+ vssd1 vccd1 vccd1 _02158_ sky130_fd_sc_hd__a22o_1
XFILLER_0_12_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10623__S net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10030_ net1347 net225 net620 vssd1 vssd1 vccd1 vccd1 _00233_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_164_2901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09733__A2 net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_164_2912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06402__A top.a1.instruction\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06547__A2 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout766_X net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_197_3400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11981_ _05859_ _05863_ vssd1 vssd1 vccd1 vccd1 _05864_ sky130_fd_sc_hd__and2b_1
XANTENNA__09497__A1 _01505_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13720_ clknet_leaf_98_clk _01291_ net986 vssd1 vssd1 vccd1 vccd1 top.a1.row2\[34\]
+ sky130_fd_sc_hd__dfrtp_1
X_10932_ net1690 net212 net593 vssd1 vssd1 vccd1 vccd1 _01093_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_196_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13651_ clknet_leaf_90_clk _01230_ net1002 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[59\]
+ sky130_fd_sc_hd__dfrtp_1
X_10863_ net248 net2187 net594 vssd1 vssd1 vccd1 vccd1 _01024_ sky130_fd_sc_hd__mux2_1
X_12602_ clknet_leaf_1_clk _00194_ net916 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[3\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_13582_ clknet_leaf_123_clk _01169_ net970 vssd1 vssd1 vccd1 vccd1 net104 sky130_fd_sc_hd__dfrtp_1
X_10794_ net264 top.DUT.register\[27\]\[2\] net598 vssd1 vssd1 vccd1 vccd1 _00955_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_183_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08990__C _03861_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12533_ clknet_leaf_30_clk _00125_ net1019 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[1\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13155__RESET_B net1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09168__A_N _02808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07680__B1 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12464_ clknet_leaf_121_clk _00059_ net933 vssd1 vssd1 vccd1 vccd1 top.ramstore\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_478 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11415_ top.a1.dataIn\[17\] _05293_ _05294_ _05295_ vssd1 vssd1 vccd1 vccd1 _05298_
+ sky130_fd_sc_hd__a2bb2o_1
X_12395_ clknet_leaf_104_clk top.ru.next_FetchedInstr\[7\] net972 vssd1 vssd1 vccd1
+ vccd1 top.a1.instruction\[7\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__08999__A _03505_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_794 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_2170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11346_ _05210_ _05213_ vssd1 vssd1 vccd1 vccd1 _05229_ sky130_fd_sc_hd__nand2_1
XFILLER_0_104_282 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06786__A2 net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10533__S net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11277_ top.a1.row2\[10\] _05139_ _05145_ top.a1.row2\[18\] _05167_ vssd1 vssd1 vccd1
+ vccd1 _05168_ sky130_fd_sc_hd__a221o_1
XANTENNA__09607__B net139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_207_802 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13016_ clknet_leaf_128_clk _00608_ net911 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[16\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_10228_ net142 net1902 net394 vssd1 vssd1 vccd1 vccd1 _00408_ sky130_fd_sc_hd__mux2_1
XFILLER_0_206_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold2 top.ru.state\[2\] vssd1 vssd1 vccd1 vccd1 net1118 sky130_fd_sc_hd__dlygate4sd3_1
X_10159_ net1531 net210 net604 vssd1 vssd1 vccd1 vccd1 _00358_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09623__A _04658_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_68 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07499__B1 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_742 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09061__C _03854_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06710__A2 net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_44_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07370_ top.DUT.register\[21\]\[8\] net656 net648 top.DUT.register\[22\]\[8\] _02508_
+ vssd1 vssd1 vccd1 vccd1 _02509_ sky130_fd_sc_hd__a221o_1
XFILLER_0_84_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06321_ top.pad.count\[0\] top.pad.count\[1\] vssd1 vssd1 vccd1 vccd1 net119 sky130_fd_sc_hd__and2b_1
XFILLER_0_29_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10708__S net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09660__A1 top.a1.halfData\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09040_ _03044_ _03145_ _03180_ _04114_ vssd1 vssd1 vccd1 vccd1 _04115_ sky130_fd_sc_hd__or4_1
X_06252_ net1684 net852 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedData\[13\] sky130_fd_sc_hd__and2_1
XFILLER_0_5_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07671__B1 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_107_Left_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06183_ top.a1.hexop\[3\] _01419_ _01422_ _01385_ vssd1 vssd1 vccd1 vccd1 _01423_
+ sky130_fd_sc_hd__o2bb2a_1
Xhold402 top.DUT.register\[14\]\[29\] vssd1 vssd1 vccd1 vccd1 net1518 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_331 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold413 top.DUT.register\[28\]\[0\] vssd1 vssd1 vccd1 vccd1 net1529 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07423__B1 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold424 top.DUT.register\[22\]\[13\] vssd1 vssd1 vccd1 vccd1 net1540 sky130_fd_sc_hd__dlygate4sd3_1
Xhold435 top.DUT.register\[25\]\[10\] vssd1 vssd1 vccd1 vccd1 net1551 sky130_fd_sc_hd__dlygate4sd3_1
Xhold446 top.DUT.register\[1\]\[17\] vssd1 vssd1 vccd1 vccd1 net1562 sky130_fd_sc_hd__dlygate4sd3_1
Xhold457 top.DUT.register\[24\]\[3\] vssd1 vssd1 vccd1 vccd1 net1573 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_187_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold468 top.DUT.register\[15\]\[6\] vssd1 vssd1 vccd1 vccd1 net1584 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09076__Y _04151_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09942_ net2290 net142 net633 vssd1 vssd1 vccd1 vccd1 _00152_ sky130_fd_sc_hd__mux2_1
XANTENNA__10443__S net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold479 top.DUT.register\[19\]\[30\] vssd1 vssd1 vccd1 vccd1 net1595 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout904 _01408_ vssd1 vssd1 vccd1 vccd1 net904 sky130_fd_sc_hd__clkbuf_4
Xfanout915 net922 vssd1 vssd1 vccd1 vccd1 net915 sky130_fd_sc_hd__clkbuf_4
Xfanout926 net928 vssd1 vssd1 vccd1 vccd1 net926 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_55_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09715__A2 net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout937 net939 vssd1 vssd1 vccd1 vccd1 net937 sky130_fd_sc_hd__clkbuf_4
X_09873_ _04882_ _04883_ _04878_ vssd1 vssd1 vccd1 vccd1 _04884_ sky130_fd_sc_hd__o21ai_1
Xfanout948 net951 vssd1 vssd1 vccd1 vccd1 net948 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_209_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout294_A net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout959 net962 vssd1 vssd1 vccd1 vccd1 net959 sky130_fd_sc_hd__clkbuf_4
X_08824_ _03198_ _03201_ vssd1 vssd1 vccd1 vccd1 _03937_ sky130_fd_sc_hd__and2_1
Xhold1102 top.DUT.register\[2\]\[31\] vssd1 vssd1 vccd1 vccd1 net2218 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_146_2631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1113 top.DUT.register\[4\]\[12\] vssd1 vssd1 vccd1 vccd1 net2229 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12460__RESET_B net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_146_2642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1124 top.DUT.register\[29\]\[13\] vssd1 vssd1 vccd1 vccd1 net2240 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1135 top.DUT.register\[25\]\[6\] vssd1 vssd1 vccd1 vccd1 net2251 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1146 top.DUT.register\[6\]\[6\] vssd1 vssd1 vccd1 vccd1 net2262 sky130_fd_sc_hd__dlygate4sd3_1
X_08755_ _02221_ _03851_ _02220_ vssd1 vssd1 vccd1 vccd1 _03871_ sky130_fd_sc_hd__a21oi_1
Xhold1157 top.DUT.register\[23\]\[11\] vssd1 vssd1 vccd1 vccd1 net2273 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_116_Left_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout461_A net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09479__A1 net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1168 top.DUT.register\[1\]\[4\] vssd1 vssd1 vccd1 vccd1 net2284 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_206_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1179 top.pad.keyCode\[3\] vssd1 vssd1 vccd1 vccd1 net2295 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09479__B2 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout559_A _01532_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11286__A1 top.a1.row2\[35\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07706_ top.DUT.register\[11\]\[4\] net525 net513 top.DUT.register\[24\]\[4\] _02844_
+ vssd1 vssd1 vccd1 vccd1 _02845_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_179_3130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08686_ net424 _03805_ vssd1 vssd1 vccd1 vccd1 _03806_ sky130_fd_sc_hd__nand2_1
X_07637_ net410 _02774_ net794 vssd1 vssd1 vccd1 vccd1 _02776_ sky130_fd_sc_hd__a21oi_2
XANTENNA_fanout726_A _01628_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout347_X net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06701__A2 net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11038__B2 top.ramload\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_192_3330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_436 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07568_ top.DUT.register\[18\]\[6\] net547 net503 top.DUT.register\[27\]\[6\] vssd1
+ vssd1 vccd1 vccd1 _02707_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_153_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09307_ _02399_ _02408_ _04370_ vssd1 vssd1 vccd1 vccd1 _04371_ sky130_fd_sc_hd__or3_1
X_06519_ _01571_ _01656_ vssd1 vssd1 vccd1 vccd1 _01658_ sky130_fd_sc_hd__nand2_1
XANTENNA__10618__S net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_192_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout514_X net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07499_ top.DUT.register\[4\]\[14\] net669 net724 top.DUT.register\[29\]\[14\] _02637_
+ vssd1 vssd1 vccd1 vccd1 _02638_ sky130_fd_sc_hd__a221o_1
X_09238_ _04304_ _04305_ vssd1 vssd1 vccd1 vccd1 _04306_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_118_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_125_Left_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_161_631 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08206__A2 net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09169_ top.pc\[5\] _02808_ vssd1 vssd1 vccd1 vccd1 _04241_ sky130_fd_sc_hd__and2b_1
XFILLER_0_133_366 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11200_ _05106_ net1270 net471 vssd1 vssd1 vccd1 vccd1 _01250_ sky130_fd_sc_hd__mux2_1
XANTENNA__07414__B1 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_170_2993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12180_ _05904_ _05083_ net848 net1852 vssd1 vssd1 vccd1 vccd1 _01288_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__06768__A2 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11131_ net57 net869 vssd1 vssd1 vccd1 vccd1 _05071_ sky130_fd_sc_hd__and2_1
XANTENNA__10353__S net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09427__B _04471_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold980 top.DUT.register\[16\]\[30\] vssd1 vssd1 vccd1 vccd1 net2096 sky130_fd_sc_hd__dlygate4sd3_1
Xhold991 top.DUT.register\[22\]\[5\] vssd1 vssd1 vccd1 vccd1 net2107 sky130_fd_sc_hd__dlygate4sd3_1
X_11062_ net77 net871 net835 net1199 vssd1 vssd1 vccd1 vccd1 _01173_ sky130_fd_sc_hd__a22o_1
XANTENNA__08914__B1 _03184_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10013_ net689 _04718_ _04952_ vssd1 vssd1 vccd1 vccd1 _04953_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_134_Left_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input22_A DAT_I[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06940__A2 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11964_ _05841_ _05843_ _05845_ _05825_ vssd1 vssd1 vccd1 vccd1 _05847_ sky130_fd_sc_hd__a31o_2
XANTENNA__08059__A _01810_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13703_ clknet_leaf_96_clk _01274_ net984 vssd1 vssd1 vccd1 vccd1 top.a1.row2\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10915_ net2277 net161 net481 vssd1 vssd1 vccd1 vccd1 _01076_ sky130_fd_sc_hd__mux2_1
XFILLER_0_168_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_184_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11895_ _05770_ _05777_ vssd1 vssd1 vccd1 vccd1 _05778_ sky130_fd_sc_hd__or2_1
XFILLER_0_196_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_184_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13634_ clknet_leaf_72_clk _01221_ net1084 vssd1 vssd1 vccd1 vccd1 net61 sky130_fd_sc_hd__dfrtp_1
X_10846_ net1643 net180 net477 vssd1 vssd1 vccd1 vccd1 _01007_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10595__Y _04991_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_767 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13565_ clknet_leaf_105_clk _01152_ net968 vssd1 vssd1 vccd1 vccd1 top.ramload\[26\]
+ sky130_fd_sc_hd__dfrtp_2
XPHY_EDGE_ROW_143_Left_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10777_ net1655 net216 net483 vssd1 vssd1 vccd1 vccd1 _00938_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12516_ clknet_leaf_76_clk _00108_ net1083 vssd1 vssd1 vccd1 vccd1 top.pc\[28\] sky130_fd_sc_hd__dfstp_2
XFILLER_0_125_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_23_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07653__B1 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13496_ clknet_leaf_125_clk _01088_ net923 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[31\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_112_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12447_ clknet_leaf_75_clk _00043_ net1080 vssd1 vssd1 vccd1 vccd1 top.ramaddr\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_139 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_1895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12378_ clknet_leaf_108_clk top.ru.next_FetchedData\[22\] net975 vssd1 vssd1 vccd1
+ vccd1 top.a1.dataIn\[22\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__06759__A2 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11329_ top.a1.dataIn\[22\] _05211_ vssd1 vssd1 vccd1 vccd1 _05212_ sky130_fd_sc_hd__nand2_1
XANTENNA__10263__S net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_572 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09905__X _04913_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_152_Left_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_56 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06870_ top.DUT.register\[25\]\[18\] net457 net505 top.DUT.register\[27\]\[18\] _02008_
+ vssd1 vssd1 vccd1 vccd1 _02009_ sky130_fd_sc_hd__a221o_1
XANTENNA__07184__A2 net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_2361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_2372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08540_ _02434_ _03665_ vssd1 vssd1 vccd1 vccd1 _03666_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_141_2561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08471_ _03248_ _03252_ vssd1 vssd1 vccd1 vccd1 _03600_ sky130_fd_sc_hd__and2_1
XANTENNA__11107__B net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_187_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_314 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07422_ top.DUT.register\[30\]\[9\] net758 net734 top.DUT.register\[16\]\[9\] vssd1
+ vssd1 vccd1 vccd1 _02561_ sky130_fd_sc_hd__a22o_1
XFILLER_0_147_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09800__B _04453_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07892__B1 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_161_Left_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkload79_A clknet_leaf_40_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_174_3060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07353_ top.DUT.register\[12\]\[8\] net532 net522 top.DUT.register\[10\]\[8\] vssd1
+ vssd1 vccd1 vccd1 _02492_ sky130_fd_sc_hd__a22o_1
XANTENNA__10438__S net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06304_ _01330_ _01329_ vssd1 vssd1 vccd1 vccd1 _01460_ sky130_fd_sc_hd__nor2_1
XFILLER_0_155_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07644__B1 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07284_ top.DUT.register\[29\]\[13\] net724 _02412_ _02422_ vssd1 vssd1 vccd1 vccd1
+ _02423_ sky130_fd_sc_hd__a211o_1
XFILLER_0_122_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06998__A2 net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09023_ _04094_ _04095_ _04096_ _04097_ vssd1 vssd1 vccd1 vccd1 _04098_ sky130_fd_sc_hd__or4_1
XFILLER_0_32_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06235_ top.ramload\[29\] net859 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedInstr\[29\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_86_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_170_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout307_A _02925_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_4_1__f_clk_X clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold210 top.DUT.register\[18\]\[17\] vssd1 vssd1 vccd1 vccd1 net1326 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09528__A _01810_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06504__X _01643_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold221 top.DUT.register\[31\]\[15\] vssd1 vssd1 vccd1 vccd1 net1337 sky130_fd_sc_hd__dlygate4sd3_1
X_06166_ net904 vssd1 vssd1 vccd1 vccd1 _00016_ sky130_fd_sc_hd__inv_2
XFILLER_0_41_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold232 top.DUT.register\[26\]\[18\] vssd1 vssd1 vccd1 vccd1 net1348 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold243 top.DUT.register\[19\]\[5\] vssd1 vssd1 vccd1 vccd1 net1359 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10173__S net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold254 top.a1.dataInTemp\[4\] vssd1 vssd1 vccd1 vccd1 net1370 sky130_fd_sc_hd__dlygate4sd3_1
Xhold265 top.DUT.register\[26\]\[20\] vssd1 vssd1 vccd1 vccd1 net1381 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_170_Left_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold276 top.DUT.register\[31\]\[26\] vssd1 vssd1 vccd1 vccd1 net1392 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_770 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold287 top.DUT.register\[17\]\[3\] vssd1 vssd1 vccd1 vccd1 net1403 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout701 _01643_ vssd1 vssd1 vccd1 vccd1 net701 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_70_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09962__S net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout712 net713 vssd1 vssd1 vccd1 vccd1 net712 sky130_fd_sc_hd__clkbuf_8
Xhold298 top.DUT.register\[11\]\[14\] vssd1 vssd1 vccd1 vccd1 net1414 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_594 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09925_ top.pc\[30\] _04628_ vssd1 vssd1 vccd1 vccd1 _04931_ sky130_fd_sc_hd__and2_1
XANTENNA__09815__X _04832_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout723 _01630_ vssd1 vssd1 vccd1 vccd1 net723 sky130_fd_sc_hd__clkbuf_4
Xfanout734 net737 vssd1 vssd1 vccd1 vccd1 net734 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout297_X net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout745 _01623_ vssd1 vssd1 vccd1 vccd1 net745 sky130_fd_sc_hd__buf_4
XANTENNA_fanout676_A _01548_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout756 net757 vssd1 vssd1 vccd1 vccd1 net756 sky130_fd_sc_hd__clkbuf_8
X_09856_ net1603 net176 net632 vssd1 vssd1 vccd1 vccd1 _00144_ sky130_fd_sc_hd__mux2_1
Xfanout767 net769 vssd1 vssd1 vccd1 vccd1 net767 sky130_fd_sc_hd__buf_4
XANTENNA__10901__S net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout778 net779 vssd1 vssd1 vccd1 vccd1 net778 sky130_fd_sc_hd__clkbuf_8
XANTENNA__06887__A _02016_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout789 _01508_ vssd1 vssd1 vccd1 vccd1 net789 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07175__A2 net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08807_ net281 _03328_ vssd1 vssd1 vccd1 vccd1 _03921_ sky130_fd_sc_hd__or2_1
X_09787_ top.pc\[16\] _04420_ _04799_ vssd1 vssd1 vccd1 vccd1 _04806_ sky130_fd_sc_hd__a21oi_1
X_06999_ top.DUT.register\[24\]\[20\] net514 net454 top.DUT.register\[29\]\[20\] _02137_
+ vssd1 vssd1 vccd1 vccd1 _02138_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout464_X net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06922__A2 net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08738_ net318 _03507_ vssd1 vssd1 vccd1 vccd1 _03855_ sky130_fd_sc_hd__nor2_1
XANTENNA_hold254_A top.a1.dataInTemp\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12397__Q top.a1.instruction\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08669_ _02047_ _03770_ vssd1 vssd1 vccd1 vccd1 _03789_ sky130_fd_sc_hd__and2b_1
XANTENNA_fanout631_X net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout729_X net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10700_ net1541 net258 net336 vssd1 vssd1 vccd1 vccd1 _00861_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_159_2833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11680_ _05530_ _05533_ _05549_ vssd1 vssd1 vccd1 vccd1 _05563_ sky130_fd_sc_hd__and3_1
XANTENNA__07883__B1 net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10631_ net264 net1662 net342 vssd1 vssd1 vccd1 vccd1 _00795_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_81_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10348__S net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09624__A1 _04658_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13350_ clknet_leaf_40_clk _00942_ net1047 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[26\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_119_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10562_ _04718_ _04952_ net399 vssd1 vssd1 vccd1 vccd1 _04990_ sky130_fd_sc_hd__and3_1
X_12301_ _01494_ _01495_ _06110_ _06111_ vssd1 vssd1 vccd1 vccd1 _06112_ sky130_fd_sc_hd__o211a_1
XFILLER_0_17_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_595 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06989__A2 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13281_ clknet_leaf_115_clk _00873_ net963 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[24\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10493_ net1707 net150 net363 vssd1 vssd1 vccd1 vccd1 _00663_ sky130_fd_sc_hd__mux2_1
XANTENNA__08613__Y _03736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_388 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12232_ top.lcd.cnt_20ms\[8\] _06069_ vssd1 vssd1 vccd1 vccd1 _06070_ sky130_fd_sc_hd__and2_1
XFILLER_0_133_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06414__X _01553_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12382__RESET_B net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12163_ net1289 net846 net796 _06045_ vssd1 vssd1 vccd1 vccd1 _01274_ sky130_fd_sc_hd__a22o_1
XANTENNA__09157__B _02849_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10083__S net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11114_ net905 net1611 net860 _05062_ vssd1 vssd1 vccd1 vccd1 _01208_ sky130_fd_sc_hd__a31o_1
XFILLER_0_102_594 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12094_ _05951_ _05974_ _05968_ _05962_ vssd1 vssd1 vccd1 vccd1 _05977_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_207_3546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11045_ net26 net838 net816 net2104 vssd1 vssd1 vccd1 vccd1 _01157_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_207_3557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10811__S net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07166__A2 _02304_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06913__A2 net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12996_ clknet_leaf_37_clk _00588_ net1051 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[15\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_99_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_204_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_12__f_clk_X clknet_4_12__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11947_ net128 _05818_ _05798_ _05812_ vssd1 vssd1 vccd1 vccd1 _05830_ sky130_fd_sc_hd__a211o_1
XFILLER_0_143_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_28_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09863__A1 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_2291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11878_ _05677_ _05708_ _05743_ vssd1 vssd1 vccd1 vccd1 _05761_ sky130_fd_sc_hd__and3_1
XFILLER_0_129_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08517__A net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_184_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13617_ clknet_leaf_71_clk _01204_ net1084 vssd1 vssd1 vccd1 vccd1 net43 sky130_fd_sc_hd__dfrtp_1
XANTENNA__10258__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10829_ net1593 net251 net477 vssd1 vssd1 vccd1 vccd1 _00990_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08418__A2 net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_1924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13548_ clknet_leaf_104_clk _01135_ net973 vssd1 vssd1 vccd1 vccd1 top.ramload\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07626__B1 net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_1935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_478 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13479_ clknet_leaf_8_clk _01071_ net945 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[30\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_124_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11230__X _05123_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09379__B1 _04438_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_678 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07971_ top.DUT.register\[10\]\[31\] net520 net453 top.DUT.register\[29\]\[31\] _03109_
+ vssd1 vssd1 vccd1 vccd1 _03110_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_52_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09710_ _03488_ net404 net490 _04740_ vssd1 vssd1 vccd1 vccd1 _04741_ sky130_fd_sc_hd__o211a_4
X_06922_ top.DUT.register\[8\]\[21\] net542 _02060_ vssd1 vssd1 vccd1 vccd1 _02061_
+ sky130_fd_sc_hd__a21o_1
XANTENNA__10721__S net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07157__A2 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08354__A1 _03342_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09083__A top.a1.instruction\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08354__B2 net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09641_ _04676_ _04679_ _04682_ vssd1 vssd1 vccd1 vccd1 _04683_ sky130_fd_sc_hd__or3_1
X_06853_ _01985_ _01988_ _01991_ vssd1 vssd1 vccd1 vccd1 _01992_ sky130_fd_sc_hd__or3_1
XANTENNA__06904__A2 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09572_ top.a1.instruction\[29\] net821 net422 vssd1 vssd1 vccd1 vccd1 _04620_ sky130_fd_sc_hd__a21o_2
XFILLER_0_89_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06784_ top.DUT.register\[17\]\[17\] net460 net512 top.DUT.register\[24\]\[17\] _01922_
+ vssd1 vssd1 vccd1 vccd1 _01923_ sky130_fd_sc_hd__a221o_1
X_08523_ net309 _03649_ vssd1 vssd1 vccd1 vccd1 _03650_ sky130_fd_sc_hd__nand2_1
XFILLER_0_148_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10957__A _04657_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08454_ net282 _03284_ _03314_ net280 vssd1 vssd1 vccd1 vccd1 _03584_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_9_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07865__B1 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_187_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_172_3019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07405_ _02534_ _02543_ vssd1 vssd1 vccd1 vccd1 _02544_ sky130_fd_sc_hd__nor2_8
XPHY_EDGE_ROW_186_Right_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10168__S net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08385_ _03516_ vssd1 vssd1 vccd1 vccd1 _03517_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout424_A net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10395__C net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09957__S net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire409 _02972_ vssd1 vssd1 vccd1 vccd1 net409 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_135_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07617__B1 net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07336_ _02443_ _02452_ _02473_ vssd1 vssd1 vccd1 vccd1 _02475_ sky130_fd_sc_hd__or3_1
XFILLER_0_116_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_154_2752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_154_2763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07267_ top.DUT.register\[20\]\[13\] net566 net526 top.DUT.register\[11\]\[13\] vssd1
+ vssd1 vccd1 vccd1 _02406_ sky130_fd_sc_hd__a22o_1
XFILLER_0_5_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09006_ _03785_ _03816_ vssd1 vssd1 vccd1 vccd1 _04081_ sky130_fd_sc_hd__nand2_1
X_06218_ top.ramload\[12\] net857 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedInstr\[12\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_20_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08162__A _01897_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07198_ _02336_ vssd1 vssd1 vccd1 vccd1 _02337_ sky130_fd_sc_hd__inv_2
XANTENNA__11177__B1 net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_187_3251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06149_ top.a1.instruction\[13\] vssd1 vssd1 vccd1 vccd1 _01392_ sky130_fd_sc_hd__inv_2
XANTENNA__07396__A2 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09692__S net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout581_X net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout520 net522 vssd1 vssd1 vccd1 vccd1 net520 sky130_fd_sc_hd__buf_4
Xfanout531 _01542_ vssd1 vssd1 vccd1 vccd1 net531 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_6_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout679_X net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout542 _01540_ vssd1 vssd1 vccd1 vccd1 net542 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10631__S net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09908_ _03987_ net404 net489 _04915_ vssd1 vssd1 vccd1 vccd1 _04916_ sky130_fd_sc_hd__o211a_4
Xfanout553 _01535_ vssd1 vssd1 vccd1 vccd1 net553 sky130_fd_sc_hd__clkbuf_8
Xfanout564 _01528_ vssd1 vssd1 vccd1 vccd1 net564 sky130_fd_sc_hd__clkbuf_4
Xfanout575 net578 vssd1 vssd1 vccd1 vccd1 net575 sky130_fd_sc_hd__clkbuf_8
XANTENNA__07148__A2 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout586 _01513_ vssd1 vssd1 vccd1 vccd1 net586 sky130_fd_sc_hd__buf_4
Xfanout597 _04966_ vssd1 vssd1 vccd1 vccd1 net597 sky130_fd_sc_hd__buf_4
X_09839_ _04843_ _04852_ _04851_ vssd1 vssd1 vccd1 vccd1 _04853_ sky130_fd_sc_hd__a21oi_1
X_12850_ clknet_leaf_22_clk _00442_ net1024 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[11\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_197_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11801_ _05636_ _05683_ vssd1 vssd1 vccd1 vccd1 _05684_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_202_3476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12781_ clknet_leaf_42_clk _00373_ net1057 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[8\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_96_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_200_148 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11732_ _05495_ _05614_ vssd1 vssd1 vccd1 vccd1 _05615_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_194_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06409__X _01548_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07320__A2 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_575 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11663_ _05498_ _05538_ _05544_ _05545_ vssd1 vssd1 vccd1 vccd1 _05546_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__10078__S net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_153_Right_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_166_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13402_ clknet_leaf_0_clk _00994_ net916 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[28\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_10614_ net205 net1828 net349 vssd1 vssd1 vccd1 vccd1 _00779_ sky130_fd_sc_hd__mux2_1
X_11594_ net234 _05476_ vssd1 vssd1 vccd1 vccd1 _05477_ sky130_fd_sc_hd__nand2_1
X_13333_ clknet_leaf_32_clk _00925_ net1044 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[26\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_106_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10545_ net2043 net188 net354 vssd1 vssd1 vccd1 vccd1 _00712_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_130_clk clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_130_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__10806__S net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_623 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13264_ clknet_leaf_29_clk _00856_ net1018 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[23\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_10476_ net1859 net207 net362 vssd1 vssd1 vccd1 vccd1 _00646_ sky130_fd_sc_hd__mux2_1
X_12215_ top.lcd.cnt_20ms\[1\] top.lcd.cnt_20ms\[0\] vssd1 vssd1 vccd1 vccd1 _06060_
+ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_94_1854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13195_ clknet_leaf_45_clk _00787_ net1069 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[21\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07387__A2 net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12146_ _06007_ _06026_ _06027_ vssd1 vssd1 vccd1 vccd1 _06029_ sky130_fd_sc_hd__or3_1
XFILLER_0_102_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_391 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06595__B1 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08800__A net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10541__S net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12077_ _05958_ _05959_ vssd1 vssd1 vccd1 vccd1 _05960_ sky130_fd_sc_hd__nor2_1
XANTENNA__09615__B _04657_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07139__A2 net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09107__S _04045_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11028_ net7 net841 net818 top.ramload\[14\] vssd1 vssd1 vccd1 vccd1 _01140_ sky130_fd_sc_hd__a22o_1
XFILLER_0_204_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_154_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_125_2320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_177_807 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09053__D _03626_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12979_ clknet_leaf_121_clk _00571_ net933 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[15\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08518__Y _03645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11225__X _05118_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07311__A2 net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_170_58 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_120_Right_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_103_1994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08170_ _02155_ net329 vssd1 vssd1 vccd1 vccd1 _03308_ sky130_fd_sc_hd__nand2_1
XFILLER_0_15_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_510 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_212 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07121_ _02244_ _02250_ _02259_ vssd1 vssd1 vccd1 vccd1 _02260_ sky130_fd_sc_hd__nor3_1
XFILLER_0_132_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_172_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10716__S net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_121_clk clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_121_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_125_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_179_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_2482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_136_2493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06822__A1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09078__A top.a1.instruction\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07052_ top.DUT.register\[18\]\[22\] net550 net516 top.DUT.register\[7\]\[22\] vssd1
+ vssd1 vccd1 vccd1 _02191_ sky130_fd_sc_hd__a22o_1
XFILLER_0_70_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput101 net101 vssd1 vssd1 vccd1 vccd1 DAT_O[6] sky130_fd_sc_hd__buf_2
XFILLER_0_42_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput112 net112 vssd1 vssd1 vccd1 vccd1 gpio_out[10] sky130_fd_sc_hd__buf_2
Xoutput123 net123 vssd1 vssd1 vccd1 vccd1 gpio_out[8] sky130_fd_sc_hd__buf_2
XFILLER_0_140_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07378__A2 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06586__B1 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_195_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10451__S net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07954_ _01834_ _03092_ vssd1 vssd1 vccd1 vccd1 _03093_ sky130_fd_sc_hd__nor2_1
XFILLER_0_49_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_182_3170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_182_3181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06905_ top.DUT.register\[1\]\[18\] net756 _02036_ _02037_ _02043_ vssd1 vssd1 vccd1
+ vccd1 _02044_ sky130_fd_sc_hd__a2111o_1
XANTENNA__06230__A top.ramload\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07885_ top.DUT.register\[7\]\[1\] net517 net441 top.DUT.register\[5\]\[1\] vssd1
+ vssd1 vccd1 vccd1 _03024_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout374_A _04981_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_207_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09624_ _04658_ _04667_ _04660_ _04659_ vssd1 vssd1 vccd1 vccd1 _04669_ sky130_fd_sc_hd__o211a_1
XFILLER_0_97_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06836_ top.DUT.register\[22\]\[19\] net577 _01974_ vssd1 vssd1 vccd1 vccd1 _01975_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_168_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07550__A2 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09555_ _04600_ _04603_ vssd1 vssd1 vccd1 vccd1 _04604_ sky130_fd_sc_hd__xor2_1
X_06767_ _01901_ _01903_ _01904_ _01905_ vssd1 vssd1 vccd1 vccd1 _01906_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout541_A _01540_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout639_A _01619_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08506_ _02310_ net494 _03626_ net428 _03624_ vssd1 vssd1 vccd1 vccd1 _03634_ sky130_fd_sc_hd__a221o_1
XANTENNA__07838__B1 net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09486_ top.pc\[24\] _01584_ vssd1 vssd1 vccd1 vccd1 _04539_ sky130_fd_sc_hd__or2_1
X_06698_ top.DUT.register\[19\]\[25\] net535 net519 top.DUT.register\[10\]\[25\] vssd1
+ vssd1 vccd1 vccd1 _01837_ sky130_fd_sc_hd__a22o_1
XANTENNA__07302__A2 net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08437_ _03566_ _03567_ vssd1 vssd1 vccd1 vccd1 _03568_ sky130_fd_sc_hd__nor2_1
XFILLER_0_92_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1071_X net1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout427_X net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_190_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_163_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08368_ net321 _03500_ _03495_ vssd1 vssd1 vccd1 vccd1 _03501_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_33_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07319_ top.DUT.register\[25\]\[12\] net778 net714 top.DUT.register\[27\]\[12\] vssd1
+ vssd1 vccd1 vccd1 _02458_ sky130_fd_sc_hd__a22o_1
XFILLER_0_151_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10626__S net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08299_ net311 _03236_ vssd1 vssd1 vccd1 vccd1 _03434_ sky130_fd_sc_hd__nand2_1
XFILLER_0_34_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_112_clk clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_112_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_6_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10330_ net1597 net269 net379 vssd1 vssd1 vccd1 vccd1 _00506_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10261_ net141 net2116 net390 vssd1 vssd1 vccd1 vccd1 _00440_ sky130_fd_sc_hd__mux2_1
XANTENNA__09212__C1 net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12000_ _05862_ _05864_ net126 vssd1 vssd1 vccd1 vccd1 _05883_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_76_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07369__A2 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10192_ _04154_ _04156_ net689 net786 vssd1 vssd1 vccd1 vccd1 _04972_ sky130_fd_sc_hd__or4b_2
XANTENNA__06577__B1 net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_167_2954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout350 net353 vssd1 vssd1 vccd1 vccd1 net350 sky130_fd_sc_hd__buf_8
XTAP_TAPCELL_ROW_204_3505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout361 net364 vssd1 vssd1 vccd1 vccd1 net361 sky130_fd_sc_hd__buf_4
XANTENNA__09515__B1 _04051_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout372 _04983_ vssd1 vssd1 vccd1 vccd1 net372 sky130_fd_sc_hd__buf_4
Xfanout383 net384 vssd1 vssd1 vccd1 vccd1 net383 sky130_fd_sc_hd__buf_4
Xfanout394 net396 vssd1 vssd1 vccd1 vccd1 net394 sky130_fd_sc_hd__clkbuf_8
X_12902_ clknet_leaf_40_clk _00494_ net1046 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[12\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_107_2050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12833_ clknet_leaf_55_clk _00425_ net1030 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[10\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_158_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09279__C1 net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12764_ clknet_leaf_130_clk _00356_ net909 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[8\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07829__B1 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08067__A _02198_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_120_2250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11715_ _05562_ _05590_ vssd1 vssd1 vccd1 vccd1 _05598_ sky130_fd_sc_hd__xnor2_1
X_12695_ clknet_leaf_3_clk _00287_ net919 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[6\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_72_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11646_ _05526_ _05527_ _05522_ vssd1 vssd1 vccd1 vccd1 _05529_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_126_236 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput14 DAT_I[20] vssd1 vssd1 vccd1 vccd1 net14 sky130_fd_sc_hd__clkbuf_1
Xinput25 DAT_I[30] vssd1 vssd1 vccd1 vccd1 net25 sky130_fd_sc_hd__clkbuf_1
Xinput36 gpio_in[16] vssd1 vssd1 vccd1 vccd1 net36 sky130_fd_sc_hd__clkbuf_1
XANTENNA__10536__S net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_103_clk clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_103_clk
+ sky130_fd_sc_hd__clkbuf_8
X_11577_ _05457_ _05458_ _05454_ _05455_ vssd1 vssd1 vccd1 vccd1 _05460_ sky130_fd_sc_hd__a211o_1
XFILLER_0_107_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13316_ clknet_leaf_36_clk _00908_ net1050 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[25\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_10528_ _04712_ _04949_ net400 vssd1 vssd1 vccd1 vccd1 _04988_ sky130_fd_sc_hd__and3_1
XFILLER_0_122_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold809 top.DUT.register\[24\]\[17\] vssd1 vssd1 vccd1 vccd1 net1925 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_149_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13247_ clknet_leaf_24_clk _00839_ net1013 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[23\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_10459_ net152 net1948 net366 vssd1 vssd1 vccd1 vccd1 _00630_ sky130_fd_sc_hd__mux2_1
X_13178_ clknet_leaf_1_clk _00770_ net916 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[21\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06568__B1 net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12129_ _05995_ _06001_ _06004_ vssd1 vssd1 vccd1 vccd1 _06012_ sky130_fd_sc_hd__or3_1
XANTENNA__10271__S net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09798__B1_N _04815_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07780__A2 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07670_ top.DUT.register\[19\]\[4\] net720 net700 top.DUT.register\[31\]\[4\] vssd1
+ vssd1 vccd1 vccd1 _02809_ sky130_fd_sc_hd__a22o_1
XFILLER_0_79_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07532__A2 net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06621_ top.DUT.register\[12\]\[27\] net534 net450 top.DUT.register\[21\]\[27\] _01759_
+ vssd1 vssd1 vccd1 vccd1 _01760_ sky130_fd_sc_hd__a221o_1
XANTENNA__09361__A _02232_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06740__B1 net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09340_ net821 _02854_ vssd1 vssd1 vccd1 vccd1 _04402_ sky130_fd_sc_hd__and2_1
XFILLER_0_75_602 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_659 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06552_ top.DUT.register\[22\]\[29\] net650 net735 top.DUT.register\[16\]\[29\] vssd1
+ vssd1 vccd1 vccd1 _01691_ sky130_fd_sc_hd__a22o_1
XANTENNA__09080__B top.a1.instruction\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12495__Q top.pc\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09271_ _01580_ _02950_ _01583_ vssd1 vssd1 vccd1 vccd1 _04337_ sky130_fd_sc_hd__o21ai_1
XANTENNA__11115__B net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06483_ net788 _01602_ _01618_ vssd1 vssd1 vccd1 vccd1 _01622_ sky130_fd_sc_hd__and3_4
XFILLER_0_173_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09690__C1 net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_2511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06209__B net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_2522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08222_ _03232_ _03253_ net276 vssd1 vssd1 vccd1 vccd1 _03359_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_16_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12414__RESET_B net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12865__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_690 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_578 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08153_ net293 _03287_ net312 vssd1 vssd1 vccd1 vccd1 _03291_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_43_532 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10446__S net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_151_2711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07599__A2 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07104_ top.DUT.register\[30\]\[16\] net759 net727 top.DUT.register\[18\]\[16\] vssd1
+ vssd1 vccd1 vccd1 _02243_ sky130_fd_sc_hd__a22o_1
XFILLER_0_70_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08084_ _03205_ _03222_ net296 vssd1 vssd1 vccd1 vccd1 _03223_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07035_ _02169_ _02171_ _02173_ vssd1 vssd1 vccd1 vccd1 _02174_ sky130_fd_sc_hd__or3_1
XFILLER_0_140_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10970__A top.a1.halfData\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_184_3210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12344__A2 net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11147__A3 _02993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout491_A _04721_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08986_ _03975_ _03993_ _04060_ _03955_ vssd1 vssd1 vccd1 vccd1 _04061_ sky130_fd_sc_hd__and4b_1
XANTENNA__09970__S net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_149_2684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07771__A2 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09823__X _04839_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07937_ _02026_ _02046_ vssd1 vssd1 vccd1 vccd1 _03076_ sky130_fd_sc_hd__and2b_1
XFILLER_0_199_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout756_A net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout377_X net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07868_ top.DUT.register\[30\]\[1\] net760 net757 top.DUT.register\[1\]\[1\] vssd1
+ vssd1 vccd1 vccd1 _03007_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_162_2873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07523__A2 net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09607_ net899 net139 vssd1 vssd1 vccd1 vccd1 _04653_ sky130_fd_sc_hd__nand2_1
XFILLER_0_97_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06819_ top.DUT.register\[25\]\[17\] net779 _01955_ _01957_ vssd1 vssd1 vccd1 vccd1
+ _01958_ sky130_fd_sc_hd__a211o_1
X_07799_ top.DUT.register\[29\]\[2\] net451 net503 top.DUT.register\[27\]\[2\] _02937_
+ vssd1 vssd1 vccd1 vccd1 _02938_ sky130_fd_sc_hd__a221o_1
XANTENNA__06731__B1 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout544_X net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_195_434 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09538_ _04586_ _04587_ vssd1 vssd1 vccd1 vccd1 _04588_ sky130_fd_sc_hd__or2_1
XFILLER_0_210_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_195_3372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout711_X net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09469_ _04521_ _04522_ vssd1 vssd1 vccd1 vccd1 _04523_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout809_X net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11500_ _05349_ _05354_ _05382_ _05351_ vssd1 vssd1 vccd1 vccd1 _05383_ sky130_fd_sc_hd__a22o_1
X_12480_ clknet_leaf_63_clk _00075_ net1090 vssd1 vssd1 vccd1 vccd1 top.ramstore\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_163_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11431_ _05313_ vssd1 vssd1 vccd1 vccd1 _05314_ sky130_fd_sc_hd__inv_2
XFILLER_0_136_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10356__S net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08236__B1 _03367_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_190_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_78_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08787__A1 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11362_ top.a1.dataIn\[27\] _05240_ _05241_ _05243_ vssd1 vssd1 vccd1 vccd1 _05245_
+ sky130_fd_sc_hd__and4b_1
XANTENNA__08251__A3 _03387_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06798__B1 net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13101_ clknet_leaf_42_clk _00693_ net1058 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[18\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10313_ net216 net1696 net384 vssd1 vssd1 vccd1 vccd1 _00490_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11293_ _05173_ _05177_ _05182_ vssd1 vssd1 vccd1 vccd1 _05183_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_91_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08621__Y _03744_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_210_3597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13032_ clknet_leaf_7_clk _00624_ net946 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[16\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11138__A3 net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10244_ net196 net1557 net390 vssd1 vssd1 vccd1 vccd1 _00423_ sky130_fd_sc_hd__mux2_1
XANTENNA__06422__X _01561_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10091__S net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10175_ net2153 net152 net605 vssd1 vssd1 vccd1 vccd1 _00374_ sky130_fd_sc_hd__mux2_1
XANTENNA__09733__X _04760_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout180 _04858_ vssd1 vssd1 vccd1 vccd1 net180 sky130_fd_sc_hd__clkbuf_2
XANTENNA__06970__B1 net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout191 _04796_ vssd1 vssd1 vccd1 vccd1 net191 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_44_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_89_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_604 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07514__A2 _02652_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08711__B2 _03829_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_186_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12816_ clknet_leaf_29_clk _00408_ net1017 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[9\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_202_788 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13796_ clknet_leaf_68_clk _01365_ vssd1 vssd1 vccd1 vccd1 top.pad.button_control.r_counter\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12747_ clknet_leaf_44_clk _00339_ net1065 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[7\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_1942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12678_ clknet_leaf_38_clk _00270_ net1054 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[5\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_13_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_1953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11629_ _05489_ _05511_ vssd1 vssd1 vccd1 vccd1 _05512_ sky130_fd_sc_hd__nor2_1
XFILLER_0_71_148 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10266__S net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09908__X _04916_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold606 top.DUT.register\[20\]\[18\] vssd1 vssd1 vccd1 vccd1 net1722 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06789__B1 net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_2441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold617 top.ru.state\[6\] vssd1 vssd1 vccd1 vccd1 net1733 sky130_fd_sc_hd__dlygate4sd3_1
Xhold628 top.DUT.register\[13\]\[25\] vssd1 vssd1 vccd1 vccd1 net1744 sky130_fd_sc_hd__dlygate4sd3_1
Xhold639 top.DUT.register\[31\]\[28\] vssd1 vssd1 vccd1 vccd1 net1755 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09727__B1 _04752_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07428__X _02567_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07147__Y _02286_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08840_ net694 _03951_ _03952_ top.pc\[26\] net884 vssd1 vssd1 vccd1 vccd1 _03953_
+ sky130_fd_sc_hd__a32o_1
XPHY_EDGE_ROW_29_Left_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07753__A2 net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08771_ net323 net429 _03530_ _03885_ vssd1 vssd1 vccd1 vccd1 _03887_ sky130_fd_sc_hd__a31o_1
XANTENNA__08950__B2 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06961__B1 net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07722_ top.DUT.register\[12\]\[3\] net741 net717 top.DUT.register\[27\]\[3\] vssd1
+ vssd1 vccd1 vccd1 _02861_ sky130_fd_sc_hd__a22o_1
XFILLER_0_79_204 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08702__A1 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11301__A3 _05128_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07653_ top.DUT.register\[9\]\[5\] net765 net739 top.DUT.register\[12\]\[5\] vssd1
+ vssd1 vccd1 vccd1 _02792_ sky130_fd_sc_hd__a22o_1
XFILLER_0_189_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06604_ _01721_ _01742_ vssd1 vssd1 vccd1 vccd1 _01743_ sky130_fd_sc_hd__nor2_1
X_07584_ _02713_ _02722_ vssd1 vssd1 vccd1 vccd1 _02723_ sky130_fd_sc_hd__nor2_8
X_09323_ net804 _02854_ _04335_ _04385_ vssd1 vssd1 vccd1 vccd1 _04386_ sky130_fd_sc_hd__o22a_2
XFILLER_0_87_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06535_ top.DUT.register\[28\]\[29\] net557 net461 top.DUT.register\[17\]\[29\] _01673_
+ vssd1 vssd1 vccd1 vccd1 _01674_ sky130_fd_sc_hd__a221o_1
XFILLER_0_165_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_123 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_38_Left_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout337_A _04995_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_459 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09254_ _04319_ _04320_ vssd1 vssd1 vccd1 vccd1 _04321_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout1079_A net1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06466_ _01595_ _01604_ vssd1 vssd1 vccd1 vccd1 _01605_ sky130_fd_sc_hd__nor2_4
XFILLER_0_173_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08205_ _03334_ _03336_ net494 _03044_ _03337_ vssd1 vssd1 vccd1 vccd1 _03343_ sky130_fd_sc_hd__a221o_1
XFILLER_0_16_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10176__S net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13043__CLK clknet_leaf_120_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09185_ _04255_ vssd1 vssd1 vccd1 vccd1 _04256_ sky130_fd_sc_hd__inv_2
XANTENNA__06492__A2 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06397_ net685 _01512_ _01531_ vssd1 vssd1 vccd1 vccd1 _01536_ sky130_fd_sc_hd__and3_1
XFILLER_0_90_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout504_A _01567_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_190_3291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08769__A1 net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08136_ _02633_ net327 vssd1 vssd1 vccd1 vccd1 _03274_ sky130_fd_sc_hd__nand2_1
XANTENNA__09965__S net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_160_367 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08067_ _02198_ net300 vssd1 vssd1 vccd1 vccd1 _03206_ sky130_fd_sc_hd__nand2_1
XFILLER_0_31_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10904__S net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07018_ top.DUT.register\[21\]\[20\] net658 net721 top.DUT.register\[19\]\[20\] vssd1
+ vssd1 vccd1 vccd1 _02157_ sky130_fd_sc_hd__a22o_1
XANTENNA__09718__B1 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07992__A2 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08170__A _02155_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout873_A net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout494_X net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_164_2902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_164_2913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07744__A2 net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout661_X net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08969_ net415 net691 net1162 net875 vssd1 vssd1 vccd1 vccd1 _00075_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA_fanout759_X net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11980_ _05755_ _05851_ _05835_ vssd1 vssd1 vccd1 vccd1 _05863_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_197_3401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10931_ net1507 net221 net593 vssd1 vssd1 vccd1 vccd1 _01092_ sky130_fd_sc_hd__mux2_1
X_10862_ net243 net1770 net594 vssd1 vssd1 vccd1 vccd1 _01023_ sky130_fd_sc_hd__mux2_1
X_13650_ clknet_leaf_89_clk _01229_ net1004 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[58\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_195_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06180__B2 net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12601_ clknet_leaf_14_clk _00193_ net955 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[3\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11056__A2 net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13581_ clknet_leaf_75_clk net1293 net1081 vssd1 vssd1 vccd1 vccd1 net103 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10793_ net270 net1682 net601 vssd1 vssd1 vccd1 vccd1 _00954_ sky130_fd_sc_hd__mux2_1
XFILLER_0_149_692 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12532_ clknet_leaf_54_clk _00124_ net1037 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[1\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_170_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_191_470 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10086__S net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12463_ clknet_leaf_75_clk _00058_ net1083 vssd1 vssd1 vccd1 vccd1 top.ramstore\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11414_ top.a1.dataIn\[17\] _05293_ _05296_ vssd1 vssd1 vccd1 vccd1 _05297_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_50_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09875__S net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12394_ clknet_leaf_95_clk top.ru.next_FetchedInstr\[6\] net981 vssd1 vssd1 vccd1
+ vccd1 top.a1.instruction\[6\] sky130_fd_sc_hd__dfrtp_2
XANTENNA_clkbuf_leaf_73_clk_A clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11345_ _05212_ _05219_ top.a1.dataIn\[23\] vssd1 vssd1 vccd1 vccd1 _05228_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_132_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10814__S net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_2171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08080__A _01940_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11276_ top.a1.row2\[26\] _05142_ _05150_ top.a1.row1\[106\] vssd1 vssd1 vccd1 vccd1
+ _05167_ sky130_fd_sc_hd__a22o_1
X_13015_ clknet_leaf_129_clk _00607_ net912 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[16\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_10227_ net149 net2069 net394 vssd1 vssd1 vccd1 vccd1 _00407_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_88_clk_A clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_207_814 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07735__A2 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10158_ net2087 net211 net602 vssd1 vssd1 vccd1 vccd1 _00357_ sky130_fd_sc_hd__mux2_1
XFILLER_0_146_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06943__B1 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold3 top.pad.button_control.debounce vssd1 vssd1 vccd1 vccd1 net1119 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09623__B net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10089_ net2155 net231 net612 vssd1 vssd1 vccd1 vccd1 _00290_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_11_clk_A clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_202_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_18_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_754 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_202_563 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_174_404 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13066__CLK clknet_leaf_120_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_26_clk_A clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13779_ clknet_leaf_69_clk _01350_ net1097 vssd1 vssd1 vccd1 vccd1 top.pad.count\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08526__Y _03653_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06320_ top.pad.count\[1\] top.pad.count\[0\] vssd1 vssd1 vccd1 vccd1 net118 sky130_fd_sc_hd__and2b_1
XFILLER_0_29_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_155_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06251_ top.ramload\[12\] net852 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedData\[12\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_154_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_619 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_362 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06182_ net888 _01422_ _01419_ net1464 vssd1 vssd1 vccd1 vccd1 _00008_ sky130_fd_sc_hd__a2bb2o_1
Xhold403 top.DUT.register\[20\]\[5\] vssd1 vssd1 vccd1 vccd1 net1519 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold414 top.DUT.register\[28\]\[27\] vssd1 vssd1 vccd1 vccd1 net1530 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10724__S net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold425 top.DUT.register\[24\]\[4\] vssd1 vssd1 vccd1 vccd1 net1541 sky130_fd_sc_hd__dlygate4sd3_1
Xhold436 top.DUT.register\[13\]\[17\] vssd1 vssd1 vccd1 vccd1 net1552 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold447 top.DUT.register\[25\]\[8\] vssd1 vssd1 vccd1 vccd1 net1563 sky130_fd_sc_hd__dlygate4sd3_1
Xhold458 top.DUT.register\[1\]\[11\] vssd1 vssd1 vccd1 vccd1 net1574 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07974__A2 net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold469 top.DUT.register\[5\]\[12\] vssd1 vssd1 vccd1 vccd1 net1585 sky130_fd_sc_hd__dlygate4sd3_1
X_09941_ net491 _04939_ _04945_ vssd1 vssd1 vccd1 vccd1 _04946_ sky130_fd_sc_hd__and3_2
XFILLER_0_40_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout905 _01405_ vssd1 vssd1 vccd1 vccd1 net905 sky130_fd_sc_hd__clkbuf_4
Xfanout916 net922 vssd1 vssd1 vccd1 vccd1 net916 sky130_fd_sc_hd__clkbuf_4
Xfanout927 net928 vssd1 vssd1 vccd1 vccd1 net927 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_55_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09872_ _04879_ _04880_ _04881_ _04151_ vssd1 vssd1 vccd1 vccd1 _04883_ sky130_fd_sc_hd__a31o_1
XANTENNA__07187__B1 net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06222__B net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout938 net939 vssd1 vssd1 vccd1 vccd1 net938 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08923__A1 _01659_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12180__B1 net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout949 net951 vssd1 vssd1 vccd1 vccd1 net949 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07726__A2 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08823_ _01833_ _03935_ vssd1 vssd1 vccd1 vccd1 _03936_ sky130_fd_sc_hd__xnor2_2
Xhold1103 top.DUT.register\[27\]\[16\] vssd1 vssd1 vccd1 vccd1 net2219 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_146_2632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1114 top.DUT.register\[10\]\[10\] vssd1 vssd1 vccd1 vccd1 net2230 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06934__B1 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_146_2643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout287_A net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1125 top.DUT.register\[13\]\[11\] vssd1 vssd1 vccd1 vccd1 net2241 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1136 top.DUT.register\[12\]\[24\] vssd1 vssd1 vccd1 vccd1 net2252 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1147 top.a1.row2\[33\] vssd1 vssd1 vccd1 vccd1 net2263 sky130_fd_sc_hd__dlygate4sd3_1
X_08754_ net1296 net830 net800 _03870_ vssd1 vssd1 vccd1 vccd1 _00040_ sky130_fd_sc_hd__a22o_1
Xhold1158 top.DUT.register\[30\]\[26\] vssd1 vssd1 vccd1 vccd1 net2274 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1169 top.DUT.register\[26\]\[2\] vssd1 vssd1 vccd1 vccd1 net2285 sky130_fd_sc_hd__dlygate4sd3_1
X_07705_ top.DUT.register\[14\]\[4\] net585 net573 top.DUT.register\[23\]\[4\] vssd1
+ vssd1 vccd1 vccd1 _02844_ sky130_fd_sc_hd__a22o_1
X_08685_ _02007_ _03804_ vssd1 vssd1 vccd1 vccd1 _03805_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_179_3131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout454_A _01561_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_92_clk clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_92_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_95_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07636_ net410 _02725_ vssd1 vssd1 vccd1 vccd1 _02775_ sky130_fd_sc_hd__or2_1
XFILLER_0_48_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_178_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_192_3320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07567_ top.DUT.register\[14\]\[6\] net583 net467 top.DUT.register\[9\]\[6\] _02705_
+ vssd1 vssd1 vccd1 vccd1 _02706_ sky130_fd_sc_hd__a221o_1
XANTENNA__08439__B1 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_192_3331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout621_A net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09306_ net804 _02901_ _04335_ _04369_ vssd1 vssd1 vccd1 vccd1 _04370_ sky130_fd_sc_hd__o22a_2
XANTENNA_fanout719_A _01635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06518_ _01571_ _01656_ vssd1 vssd1 vccd1 vccd1 _01657_ sky130_fd_sc_hd__nor2_1
XFILLER_0_76_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08165__A _02069_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07498_ top.DUT.register\[23\]\[14\] net674 net772 top.DUT.register\[10\]\[14\] vssd1
+ vssd1 vccd1 vccd1 _02637_ sky130_fd_sc_hd__a22o_1
XFILLER_0_17_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09237_ _02544_ _02547_ vssd1 vssd1 vccd1 vccd1 _04305_ sky130_fd_sc_hd__or2_1
XFILLER_0_161_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06449_ net896 _01389_ _01390_ _01472_ vssd1 vssd1 vccd1 vccd1 _01588_ sky130_fd_sc_hd__or4_2
XFILLER_0_133_301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_157_2794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout507_X net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_643 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09168_ _02808_ top.pc\[5\] vssd1 vssd1 vccd1 vccd1 _04240_ sky130_fd_sc_hd__and2b_1
XANTENNA_fanout990_A net1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_378 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08119_ _03163_ _03167_ vssd1 vssd1 vccd1 vccd1 _03258_ sky130_fd_sc_hd__or2_2
XFILLER_0_114_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10634__S net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09099_ _02356_ _04173_ vssd1 vssd1 vccd1 vccd1 _04174_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_170_2994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07965__A2 net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11130_ net906 net1732 net861 _05070_ vssd1 vssd1 vccd1 vccd1 _01216_ sky130_fd_sc_hd__a31o_1
Xhold970 top.DUT.register\[14\]\[1\] vssd1 vssd1 vccd1 vccd1 net2086 sky130_fd_sc_hd__dlygate4sd3_1
Xhold981 top.DUT.register\[7\]\[23\] vssd1 vssd1 vccd1 vccd1 net2097 sky130_fd_sc_hd__dlygate4sd3_1
X_11061_ net76 net870 net834 net1202 vssd1 vssd1 vccd1 vccd1 _01172_ sky130_fd_sc_hd__a22o_1
Xhold992 top.DUT.register\[3\]\[14\] vssd1 vssd1 vccd1 vccd1 net2108 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07178__B1 net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10012_ top.a1.instruction\[10\] net786 top.a1.instruction\[9\] vssd1 vssd1 vccd1
+ vccd1 _04952_ sky130_fd_sc_hd__and3b_4
XTAP_TAPCELL_ROW_110_2090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06925__B1 net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input15_A DAT_I[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11963_ _05841_ _05843_ _05845_ vssd1 vssd1 vccd1 vccd1 _05846_ sky130_fd_sc_hd__and3_1
XANTENNA__13089__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13702_ clknet_leaf_92_clk _01273_ net998 vssd1 vssd1 vccd1 vccd1 top.a1.row2\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_10914_ net2274 net166 net481 vssd1 vssd1 vccd1 vccd1 _01075_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11894_ _05773_ _05774_ _05775_ vssd1 vssd1 vccd1 vccd1 _05777_ sky130_fd_sc_hd__or3_1
XANTENNA__07350__B1 net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10845_ net1401 net194 net476 vssd1 vssd1 vccd1 vccd1 _01006_ sky130_fd_sc_hd__mux2_1
X_13633_ clknet_leaf_75_clk _01220_ net1081 vssd1 vssd1 vccd1 vccd1 net60 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_168_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10809__S net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_183_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_560 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08075__A _02026_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13564_ clknet_leaf_105_clk _01151_ net968 vssd1 vssd1 vccd1 vccd1 top.ramload\[25\]
+ sky130_fd_sc_hd__dfrtp_2
X_10776_ net1840 net224 net483 vssd1 vssd1 vccd1 vccd1 _00937_ sky130_fd_sc_hd__mux2_1
XANTENNA__10788__A1 net156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_2200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13376__RESET_B net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12515_ clknet_leaf_76_clk _00107_ net1083 vssd1 vssd1 vccd1 vccd1 top.pc\[27\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_124_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08850__B1 _03427_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13495_ clknet_leaf_3_clk _01087_ net919 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[31\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_23_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13305__RESET_B net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12446_ clknet_leaf_72_clk _00042_ net1080 vssd1 vssd1 vccd1 vccd1 top.ramaddr\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08362__X _03495_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_130_2400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12377_ clknet_leaf_109_clk top.ru.next_FetchedData\[21\] net976 vssd1 vssd1 vccd1
+ vccd1 top.a1.dataIn\[21\] sky130_fd_sc_hd__dfrtp_2
XANTENNA__10544__S net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_1896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11328_ top.a1.dataIn\[21\] top.a1.dataIn\[20\] vssd1 vssd1 vccd1 vccd1 _05211_ sky130_fd_sc_hd__or2_1
XFILLER_0_157_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11259_ _05121_ _05138_ _05144_ _05151_ vssd1 vssd1 vccd1 vccd1 _05152_ sky130_fd_sc_hd__or4_1
XFILLER_0_66_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07708__A2 net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_207_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06916__B1 net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11228__X _05121_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09353__B _04403_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_2362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_2373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06392__A1 top.a1.instruction\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_167_Right_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_50_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_74_clk clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_74_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__09330__A1 net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08470_ _03372_ _03534_ _03587_ net298 _03598_ vssd1 vssd1 vccd1 vccd1 _03599_ sky130_fd_sc_hd__o221ai_4
XANTENNA__09330__B2 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_141_2562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07341__B1 net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_175_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07421_ top.DUT.register\[14\]\[9\] net730 _02548_ _02559_ vssd1 vssd1 vccd1 vccd1
+ _02560_ sky130_fd_sc_hd__a211o_1
XANTENNA__07441__X _02580_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10719__S net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_174_3050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07352_ top.DUT.register\[24\]\[8\] net512 _02488_ _02490_ vssd1 vssd1 vccd1 vccd1
+ _02491_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_174_3061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06303_ net1085 _01453_ vssd1 vssd1 vccd1 vccd1 _01329_ sky130_fd_sc_hd__and2_1
XFILLER_0_162_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_148 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11123__B net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07283_ top.DUT.register\[22\]\[13\] net649 net717 top.DUT.register\[27\]\[13\] _02411_
+ vssd1 vssd1 vccd1 vccd1 _02422_ sky130_fd_sc_hd__a221o_1
XANTENNA__06217__B net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09022_ _02387_ _02431_ _02475_ _02524_ vssd1 vssd1 vccd1 vccd1 _04097_ sky130_fd_sc_hd__or4_1
XFILLER_0_170_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06234_ top.ramload\[28\] net859 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedInstr\[28\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_143_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold200 top.DUT.register\[18\]\[30\] vssd1 vssd1 vccd1 vccd1 net1316 sky130_fd_sc_hd__dlygate4sd3_1
X_06165_ net36 net35 net38 net37 vssd1 vssd1 vccd1 vccd1 _01408_ sky130_fd_sc_hd__nor4_1
XANTENNA__10454__S net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold211 top.DUT.register\[8\]\[24\] vssd1 vssd1 vccd1 vccd1 net1327 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout202_A _04841_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09528__B _04577_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold222 top.DUT.register\[23\]\[12\] vssd1 vssd1 vccd1 vccd1 net1338 sky130_fd_sc_hd__dlygate4sd3_1
Xhold233 top.DUT.register\[20\]\[25\] vssd1 vssd1 vccd1 vccd1 net1349 sky130_fd_sc_hd__dlygate4sd3_1
Xhold244 top.DUT.register\[23\]\[23\] vssd1 vssd1 vccd1 vccd1 net1360 sky130_fd_sc_hd__dlygate4sd3_1
Xhold255 top.DUT.register\[25\]\[14\] vssd1 vssd1 vccd1 vccd1 net1371 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06233__A top.ramload\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold266 top.DUT.register\[14\]\[14\] vssd1 vssd1 vccd1 vccd1 net1382 sky130_fd_sc_hd__dlygate4sd3_1
Xhold277 top.DUT.register\[17\]\[18\] vssd1 vssd1 vccd1 vccd1 net1393 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09149__A1 top.pc\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold288 top.DUT.register\[5\]\[22\] vssd1 vssd1 vccd1 vccd1 net1404 sky130_fd_sc_hd__dlygate4sd3_1
Xhold299 top.DUT.register\[24\]\[7\] vssd1 vssd1 vccd1 vccd1 net1415 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout702 _01642_ vssd1 vssd1 vccd1 vccd1 net702 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_70_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09924_ _04918_ _04922_ _04924_ vssd1 vssd1 vccd1 vccd1 _04930_ sky130_fd_sc_hd__or3b_1
Xfanout713 _01638_ vssd1 vssd1 vccd1 vccd1 net713 sky130_fd_sc_hd__buf_4
XFILLER_0_0_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout724 _01630_ vssd1 vssd1 vccd1 vccd1 net724 sky130_fd_sc_hd__clkbuf_8
Xfanout735 net736 vssd1 vssd1 vccd1 vccd1 net735 sky130_fd_sc_hd__clkbuf_8
Xfanout746 _01622_ vssd1 vssd1 vccd1 vccd1 net746 sky130_fd_sc_hd__clkbuf_8
XANTENNA_input7_A DAT_I[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09855_ _03890_ net404 net490 _04867_ vssd1 vssd1 vccd1 vccd1 _04868_ sky130_fd_sc_hd__o211a_2
Xfanout757 _01620_ vssd1 vssd1 vccd1 vccd1 net757 sky130_fd_sc_hd__buf_4
XANTENNA__12681__RESET_B net1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout768 net769 vssd1 vssd1 vccd1 vccd1 net768 sky130_fd_sc_hd__buf_4
XANTENNA_fanout571_A _01519_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout779 _01603_ vssd1 vssd1 vccd1 vccd1 net779 sky130_fd_sc_hd__buf_4
XANTENNA__06887__B _02025_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout669_A _01599_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08806_ net324 _03579_ _03919_ vssd1 vssd1 vccd1 vccd1 _03920_ sky130_fd_sc_hd__o21ba_1
XANTENNA__13231__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06998_ top.DUT.register\[6\]\[20\] net570 net542 top.DUT.register\[8\]\[20\] vssd1
+ vssd1 vccd1 vccd1 _02137_ sky130_fd_sc_hd__a22o_1
X_09786_ net1602 net223 net632 vssd1 vssd1 vccd1 vccd1 _00137_ sky130_fd_sc_hd__mux2_1
XANTENNA__07580__B1 net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08737_ net322 _03500_ _03535_ vssd1 vssd1 vccd1 vccd1 _03854_ sky130_fd_sc_hd__a21oi_2
XPHY_EDGE_ROW_134_Right_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout836_A net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_65_clk clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_65_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout457_X net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_3_4_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08668_ net2146 net830 net800 _03788_ vssd1 vssd1 vccd1 vccd1 _00036_ sky130_fd_sc_hd__a22o_1
XANTENNA__06686__A2 net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07619_ top.DUT.register\[29\]\[5\] net451 net508 top.DUT.register\[4\]\[5\] _02757_
+ vssd1 vssd1 vccd1 vccd1 _02758_ sky130_fd_sc_hd__a221o_1
XFILLER_0_193_521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_159_2834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10629__S net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout624_X net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08599_ _03342_ _03708_ _03722_ net496 vssd1 vssd1 vccd1 vccd1 _03723_ sky130_fd_sc_hd__o22a_1
XFILLER_0_95_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_166_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10630_ net267 net1645 net344 vssd1 vssd1 vccd1 vccd1 _00794_ sky130_fd_sc_hd__mux2_1
XFILLER_0_165_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_81_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08872__A2_N net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07635__A1 top.a1.instruction\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10561_ net1428 net140 net356 vssd1 vssd1 vccd1 vccd1 _00728_ sky130_fd_sc_hd__mux2_1
XANTENNA__07635__B2 top.a1.instruction\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12300_ top.pad.button_control.debounce top.pad.button_control.noisy vssd1 vssd1
+ vccd1 vccd1 _06111_ sky130_fd_sc_hd__nand2_1
XFILLER_0_118_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09719__A net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13280_ clknet_leaf_114_clk _00872_ net992 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[24\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_10492_ top.DUT.register\[17\]\[29\] net154 net363 vssd1 vssd1 vccd1 vccd1 _00662_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout993_X net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12231_ _06069_ net978 _06068_ vssd1 vssd1 vccd1 vccd1 _01318_ sky130_fd_sc_hd__and3b_1
XANTENNA__10364__S net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09438__B _04487_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_2130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12162_ _06043_ _06044_ vssd1 vssd1 vccd1 vccd1 _06045_ sky130_fd_sc_hd__or2_1
XANTENNA__12769__RESET_B net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11113_ net47 net864 vssd1 vssd1 vccd1 vccd1 _05062_ sky130_fd_sc_hd__and2_1
XANTENNA__06610__A2 net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12093_ _05962_ _05968_ vssd1 vssd1 vccd1 vccd1 _05976_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_9_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_208_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11044_ net25 net841 net818 net2297 vssd1 vssd1 vccd1 vccd1 _01156_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_207_3547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_207_3558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07571__B1 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09741__X _04766_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_207_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_203_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_101_Right_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_56_clk clknet_4_12__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_56_clk
+ sky130_fd_sc_hd__clkbuf_8
X_12995_ clknet_leaf_57_clk _00587_ net1076 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[15\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09312__A1 net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11946_ net128 _05818_ _05798_ vssd1 vssd1 vccd1 vccd1 _05829_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_52_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07323__B1 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_404 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06677__A2 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_2292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10539__S net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11877_ _05747_ _05756_ vssd1 vssd1 vccd1 vccd1 _05760_ sky130_fd_sc_hd__xor2_1
XANTENNA__08517__B _03440_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13616_ clknet_leaf_90_clk _01203_ net1002 vssd1 vssd1 vccd1 vccd1 net42 sky130_fd_sc_hd__dfrtp_1
X_10828_ net1816 net256 net476 vssd1 vssd1 vccd1 vccd1 _00989_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06429__A2 net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_1925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13547_ clknet_4_5__leaf_clk _01134_ net980 vssd1 vssd1 vccd1 vccd1 top.ramload\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_99_1936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10759_ net1407 net142 net419 vssd1 vssd1 vccd1 vccd1 _00920_ sky130_fd_sc_hd__mux2_1
XFILLER_0_171_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13825__1109 vssd1 vssd1 vccd1 vccd1 _13825__1109/HI net1109 sky130_fd_sc_hd__conb_1
X_13478_ clknet_leaf_38_clk _01070_ net1053 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[30\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09379__A1 _01930_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10274__S net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12429_ clknet_leaf_87_clk _00025_ net1004 vssd1 vssd1 vccd1 vccd1 top.ramaddr\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_152_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_39_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07970_ top.DUT.register\[17\]\[31\] net462 net441 top.DUT.register\[5\]\[31\] vssd1
+ vssd1 vccd1 vccd1 _03109_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_52_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06921_ top.DUT.register\[15\]\[21\] net682 net678 top.DUT.register\[31\]\[21\] vssd1
+ vssd1 vccd1 vccd1 _02060_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_52_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09000__B1 _03176_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_0__f_clk clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_0__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_06852_ top.DUT.register\[4\]\[19\] net669 net776 top.DUT.register\[13\]\[19\] _01986_
+ vssd1 vssd1 vccd1 vccd1 _01991_ sky130_fd_sc_hd__a221o_1
X_09640_ _04680_ _04681_ vssd1 vssd1 vccd1 vccd1 _04682_ sky130_fd_sc_hd__nor2_1
XANTENNA__09083__B top.a1.instruction\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_77 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09571_ _04616_ _04618_ vssd1 vssd1 vccd1 vccd1 _04619_ sky130_fd_sc_hd__xnor2_1
X_06783_ top.DUT.register\[14\]\[17\] net583 net545 top.DUT.register\[16\]\[17\] vssd1
+ vssd1 vccd1 vccd1 _01922_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_47_clk clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_47_clk
+ sky130_fd_sc_hd__clkbuf_8
X_08522_ _03600_ _03648_ net289 vssd1 vssd1 vccd1 vccd1 _03649_ sky130_fd_sc_hd__mux2_1
XFILLER_0_179_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_210_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10957__B _04998_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08965__A1_N net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_187_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08453_ _03581_ _03582_ vssd1 vssd1 vccd1 vccd1 _03583_ sky130_fd_sc_hd__nand2_1
XANTENNA__06668__A2 net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10449__S net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_175_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout152_A _04929_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07404_ _02538_ _02540_ _02542_ vssd1 vssd1 vccd1 vccd1 _02543_ sky130_fd_sc_hd__or3_2
X_08384_ _02678_ _02704_ vssd1 vssd1 vccd1 vccd1 _03516_ sky130_fd_sc_hd__nand2_1
XANTENNA__06228__A top.ramload\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_610 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07335_ _02443_ _02452_ _02473_ vssd1 vssd1 vccd1 vccd1 _02474_ sky130_fd_sc_hd__o21a_1
XFILLER_0_163_749 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1061_A net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_154_2753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07266_ top.DUT.register\[9\]\[13\] net468 net462 top.DUT.register\[17\]\[13\] _02404_
+ vssd1 vssd1 vccd1 vccd1 _02405_ sky130_fd_sc_hd__a221o_1
XFILLER_0_33_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09005_ _03750_ _03778_ _03792_ _03818_ vssd1 vssd1 vccd1 vccd1 _04080_ sky130_fd_sc_hd__and4b_1
XFILLER_0_5_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06217_ net1256 net856 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedInstr\[11\] sky130_fd_sc_hd__and2_1
XFILLER_0_103_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06840__A2 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07197_ _01473_ _01573_ vssd1 vssd1 vccd1 vccd1 _02336_ sky130_fd_sc_hd__nand2_1
XANTENNA__09973__S net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06148_ net894 vssd1 vssd1 vccd1 vccd1 _01391_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_187_3252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08730__X _03848_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11300__C top.lcd.nextState\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_203_Right_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout786_A _04708_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12059__A_N top.a1.dataIn\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10912__S net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout510 _01565_ vssd1 vssd1 vccd1 vccd1 net510 sky130_fd_sc_hd__buf_4
Xfanout521 net522 vssd1 vssd1 vccd1 vccd1 net521 sky130_fd_sc_hd__buf_4
XFILLER_0_158_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_6_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09274__A _02286_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout532 _01542_ vssd1 vssd1 vccd1 vccd1 net532 sky130_fd_sc_hd__buf_2
X_09907_ _04913_ _04914_ vssd1 vssd1 vccd1 vccd1 _04915_ sky130_fd_sc_hd__or2_1
Xfanout543 net546 vssd1 vssd1 vccd1 vccd1 net543 sky130_fd_sc_hd__clkbuf_8
Xfanout554 _01535_ vssd1 vssd1 vccd1 vccd1 net554 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout953_A net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout565 net566 vssd1 vssd1 vccd1 vccd1 net565 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout574_X net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout576 net578 vssd1 vssd1 vccd1 vccd1 net576 sky130_fd_sc_hd__buf_4
Xfanout587 net588 vssd1 vssd1 vccd1 vccd1 net587 sky130_fd_sc_hd__buf_2
X_09838_ _04842_ _04844_ vssd1 vssd1 vccd1 vccd1 _04852_ sky130_fd_sc_hd__nand2_1
XFILLER_0_198_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout598 _04965_ vssd1 vssd1 vccd1 vccd1 net598 sky130_fd_sc_hd__buf_6
XANTENNA__07553__B1 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09769_ top.pc\[15\] _04403_ vssd1 vssd1 vccd1 vccd1 _04790_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout741_X net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_38_clk clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_38_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_201_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_201_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11800_ _05637_ _05656_ _05654_ vssd1 vssd1 vccd1 vccd1 _05683_ sky130_fd_sc_hd__a21boi_1
XTAP_TAPCELL_ROW_202_3477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12780_ clknet_leaf_65_clk _00372_ net1093 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[8\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07305__B1 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09943__A_N top.a1.instruction\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06659__A2 net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11731_ _05540_ _05571_ _05539_ vssd1 vssd1 vccd1 vccd1 _05614_ sky130_fd_sc_hd__o21ai_1
XANTENNA__10359__S net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_746 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11662_ _05483_ _05484_ vssd1 vssd1 vccd1 vccd1 _05545_ sky130_fd_sc_hd__xor2_1
XFILLER_0_83_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13401_ clknet_leaf_14_clk _00993_ net956 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[28\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_154_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11979__A top.a1.dataIn\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10613_ net216 net1863 net347 vssd1 vssd1 vccd1 vccd1 _00778_ sky130_fd_sc_hd__mux2_1
X_11593_ _05432_ _05437_ _05472_ _05435_ vssd1 vssd1 vccd1 vccd1 _05476_ sky130_fd_sc_hd__a22o_2
XFILLER_0_36_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10544_ net1588 net196 net356 vssd1 vssd1 vccd1 vccd1 _00711_ sky130_fd_sc_hd__mux2_1
X_13332_ clknet_leaf_55_clk _00924_ net1073 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[26\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06425__X _01564_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06292__B1 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10094__S net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06831__A2 net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10475_ net1860 net211 net361 vssd1 vssd1 vccd1 vccd1 _00645_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13263_ clknet_leaf_22_clk _00855_ net1035 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[23\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12214_ _01384_ _06059_ net980 vssd1 vssd1 vccd1 vccd1 _01311_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_94_1855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13194_ clknet_leaf_118_clk _00786_ net954 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[21\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_121_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12145_ _06026_ _06027_ vssd1 vssd1 vccd1 vccd1 _06028_ sky130_fd_sc_hd__nor2_1
XANTENNA__10822__S net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07792__B1 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12076_ _05920_ _05957_ _05923_ vssd1 vssd1 vccd1 vccd1 _05959_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_47_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11027_ net6 net839 net817 net1684 vssd1 vssd1 vccd1 vccd1 _01139_ sky130_fd_sc_hd__o22a_1
XANTENNA__09533__A1 net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07544__B1 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10194__C_N net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06898__A2 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_29_clk clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_29_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_204_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_819 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09297__B1 top.pc\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12978_ clknet_leaf_23_clk _00570_ net1014 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[15\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10269__S net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11929_ _05810_ _05811_ vssd1 vssd1 vccd1 vccd1 _05812_ sky130_fd_sc_hd__or2_1
XFILLER_0_185_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08815__X _03929_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_103_1984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_1995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_64 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07120_ _02255_ _02256_ _02257_ _02258_ vssd1 vssd1 vccd1 vccd1 _02259_ sky130_fd_sc_hd__or4_1
XFILLER_0_70_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07075__A2 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07051_ top.DUT.register\[12\]\[22\] net532 _02189_ vssd1 vssd1 vccd1 vccd1 _02190_
+ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_136_2483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06822__A2 _01960_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09078__B top.a1.instruction\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_179_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput102 net102 vssd1 vssd1 vccd1 vccd1 DAT_O[7] sky130_fd_sc_hd__buf_2
XANTENNA__11159__B2 net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput113 net113 vssd1 vssd1 vccd1 vccd1 gpio_out[11] sky130_fd_sc_hd__buf_2
Xoutput124 net124 vssd1 vssd1 vccd1 vccd1 gpio_out[9] sky130_fd_sc_hd__buf_2
XFILLER_0_2_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_10_Left_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10732__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_195_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07953_ _01854_ _01873_ _03091_ vssd1 vssd1 vccd1 vccd1 _03092_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_182_3171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06904_ top.DUT.register\[3\]\[18\] net705 _02038_ _02039_ _02042_ vssd1 vssd1 vccd1
+ vccd1 _02043_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_182_3182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07884_ top.DUT.register\[11\]\[1\] net526 net510 top.DUT.register\[4\]\[1\] _03022_
+ vssd1 vssd1 vccd1 vccd1 _03023_ sky130_fd_sc_hd__a221o_1
XANTENNA__06230__B net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07535__B1 net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09623_ _04658_ net848 vssd1 vssd1 vccd1 vccd1 _04668_ sky130_fd_sc_hd__nor2_2
XANTENNA__09822__A net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06835_ top.DUT.register\[15\]\[19\] net682 net678 top.DUT.register\[31\]\[19\] vssd1
+ vssd1 vccd1 vccd1 _01974_ sky130_fd_sc_hd__a22o_1
XANTENNA__06889__A2 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout367_A net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06766_ top.DUT.register\[20\]\[24\] net666 net740 top.DUT.register\[12\]\[24\] _01900_
+ vssd1 vssd1 vccd1 vccd1 _01905_ sky130_fd_sc_hd__a221o_1
X_09554_ _04601_ _04602_ vssd1 vssd1 vccd1 vccd1 _04603_ sky130_fd_sc_hd__nand2_1
XFILLER_0_179_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08505_ net434 _03632_ vssd1 vssd1 vccd1 vccd1 _03633_ sky130_fd_sc_hd__nor2_1
XFILLER_0_144_71 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_176_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06697_ top.DUT.register\[22\]\[25\] net578 net555 top.DUT.register\[28\]\[25\] _01835_
+ vssd1 vssd1 vccd1 vccd1 _01836_ sky130_fd_sc_hd__a221o_1
X_09485_ top.pc\[24\] _01584_ vssd1 vssd1 vccd1 vccd1 _04538_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout534_A _01542_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09968__S net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08436_ _02525_ _03565_ vssd1 vssd1 vccd1 vccd1 _03567_ sky130_fd_sc_hd__and2_1
XFILLER_0_148_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08367_ net316 _03499_ _03497_ vssd1 vssd1 vccd1 vccd1 _03500_ sky130_fd_sc_hd__a21oi_2
XANTENNA__10907__S net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout701_A _01643_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_708 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07318_ top.DUT.register\[21\]\[12\] net655 net730 top.DUT.register\[14\]\[12\] _02456_
+ vssd1 vssd1 vccd1 vccd1 _02457_ sky130_fd_sc_hd__a221o_1
XFILLER_0_73_371 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07066__A2 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08298_ net311 _03221_ _03432_ vssd1 vssd1 vccd1 vccd1 _03433_ sky130_fd_sc_hd__o21ai_1
XANTENNA__08173__A _02026_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07249_ _02386_ _02387_ vssd1 vssd1 vccd1 vccd1 _02388_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_61_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06813__A2 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09556__X _04605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10260_ net151 net1710 net390 vssd1 vssd1 vccd1 vccd1 _00439_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout789_X net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10191_ top.a1.instruction\[11\] _04153_ _04949_ vssd1 vssd1 vccd1 vccd1 _04971_
+ sky130_fd_sc_hd__and3_4
XANTENNA__10642__S net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07774__B1 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_167_2944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07938__A_N _01940_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_167_2955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout956_X net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout340 _04993_ vssd1 vssd1 vccd1 vccd1 net340 sky130_fd_sc_hd__clkbuf_8
Xfanout351 net353 vssd1 vssd1 vccd1 vccd1 net351 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_204_3506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout362 net364 vssd1 vssd1 vccd1 vccd1 net362 sky130_fd_sc_hd__buf_4
XANTENNA__09515__B2 top.pc\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout373 _04981_ vssd1 vssd1 vccd1 vccd1 net373 sky130_fd_sc_hd__buf_6
Xfanout384 _04979_ vssd1 vssd1 vccd1 vccd1 net384 sky130_fd_sc_hd__clkbuf_8
XANTENNA__07526__B1 net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout395 net396 vssd1 vssd1 vccd1 vccd1 net395 sky130_fd_sc_hd__clkbuf_8
X_12901_ clknet_leaf_35_clk _00493_ net1040 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[12\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07804__X _02943_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13824__1108 vssd1 vssd1 vccd1 vccd1 _13824__1108/HI net1108 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_107_2051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12832_ clknet_leaf_17_clk _00424_ net964 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[10\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_96_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_201_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10089__S net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12763_ clknet_leaf_120_clk _00355_ net931 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[8\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_201_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_167_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_120_2240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_532 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06139__Y _01382_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_2251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11714_ _05589_ _05595_ vssd1 vssd1 vccd1 vccd1 _05597_ sky130_fd_sc_hd__nand2_1
X_12694_ clknet_leaf_11_clk _00286_ net948 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[6\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_83_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_204_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11645_ _05526_ _05527_ vssd1 vssd1 vccd1 vccd1 _05528_ sky130_fd_sc_hd__nand2_1
XANTENNA__10817__S net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08354__Y _03488_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08254__A1 _03263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput15 DAT_I[21] vssd1 vssd1 vccd1 vccd1 net15 sky130_fd_sc_hd__clkbuf_1
XANTENNA__07057__A2 net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08254__B2 net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11576_ _05457_ _05458_ vssd1 vssd1 vccd1 vccd1 _05459_ sky130_fd_sc_hd__nand2_1
Xinput26 DAT_I[31] vssd1 vssd1 vccd1 vccd1 net26 sky130_fd_sc_hd__clkbuf_1
Xinput37 gpio_in[17] vssd1 vssd1 vccd1 vccd1 net37 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11996__X _05879_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13315_ clknet_leaf_49_clk _00907_ net1061 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[25\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06804__A2 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10527_ net1921 net142 net358 vssd1 vssd1 vccd1 vccd1 _00696_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10458_ net158 net1861 net367 vssd1 vssd1 vccd1 vccd1 _00629_ sky130_fd_sc_hd__mux2_1
XANTENNA__09907__A _04913_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13246_ clknet_leaf_20_clk _00838_ net1029 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[23\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08557__A2 top.pc\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09754__B2 net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10552__S net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10389_ net2299 net161 net376 vssd1 vssd1 vccd1 vccd1 _00564_ sky130_fd_sc_hd__mux2_1
X_13177_ clknet_leaf_14_clk _00769_ net959 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[21\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06602__Y _01741_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12128_ _06010_ vssd1 vssd1 vccd1 vccd1 _06011_ sky130_fd_sc_hd__inv_2
XFILLER_0_165_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08309__A2 _03441_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12059_ top.a1.dataIn\[3\] _05941_ vssd1 vssd1 vccd1 vccd1 _05942_ sky130_fd_sc_hd__nand2b_2
X_06620_ top.DUT.register\[23\]\[27\] net573 net565 top.DUT.register\[20\]\[27\] vssd1
+ vssd1 vccd1 vccd1 _01759_ sky130_fd_sc_hd__a22o_1
XFILLER_0_205_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_487 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06551_ top.DUT.register\[30\]\[29\] net761 net721 top.DUT.register\[19\]\[29\] _01689_
+ vssd1 vssd1 vccd1 vccd1 _01690_ sky130_fd_sc_hd__a221o_1
XFILLER_0_47_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_47_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09270_ _01580_ _02950_ _01583_ vssd1 vssd1 vccd1 vccd1 _04336_ sky130_fd_sc_hd__o21a_1
X_06482_ net788 _01600_ _01611_ vssd1 vssd1 vccd1 vccd1 _01621_ sky130_fd_sc_hd__and3_4
XANTENNA__07296__A2 net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_185_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11092__A3 net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_2512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08221_ _03355_ _03357_ net311 vssd1 vssd1 vccd1 vccd1 _03358_ sky130_fd_sc_hd__mux2_1
XFILLER_0_173_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_16_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_2523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10727__S net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_546 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08152_ _03288_ _03289_ net287 vssd1 vssd1 vccd1 vccd1 _03290_ sky130_fd_sc_hd__and3b_1
XANTENNA__11412__A top.a1.dataIn\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07048__A2 net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_544 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07103_ _02232_ _02241_ vssd1 vssd1 vccd1 vccd1 _02242_ sky130_fd_sc_hd__nor2_4
XTAP_TAPCELL_ROW_151_2712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11131__B net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08083_ _03213_ _03221_ net311 vssd1 vssd1 vccd1 vccd1 _03222_ sky130_fd_sc_hd__mux2_1
XANTENNA__08796__A2 top.pc\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_9_clk clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_9_clk
+ sky130_fd_sc_hd__clkbuf_8
X_07034_ top.DUT.register\[14\]\[20\] net733 net716 top.DUT.register\[27\]\[20\] _02172_
+ vssd1 vssd1 vccd1 vccd1 _02173_ sky130_fd_sc_hd__a221o_1
XFILLER_0_30_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08721__A net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_184_3200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_184_3211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09745__B2 net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07756__B1 net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1024_A net1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06241__A top.ramload\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08985_ _03568_ _03896_ _03913_ _04059_ vssd1 vssd1 vccd1 vccd1 _04060_ sky130_fd_sc_hd__and4b_1
XANTENNA_fanout484_A _04962_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_149_2674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_149_2685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07936_ _01983_ _02003_ vssd1 vssd1 vccd1 vccd1 _03075_ sky130_fd_sc_hd__and2_1
XANTENNA__07508__B1 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout651_A _01610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07867_ top.DUT.register\[23\]\[1\] net674 net720 top.DUT.register\[19\]\[1\] _03005_
+ vssd1 vssd1 vccd1 vccd1 _03006_ sky130_fd_sc_hd__a221o_1
XFILLER_0_211_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_162_2874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout749_A _01622_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09606_ top.pc\[31\] _04633_ vssd1 vssd1 vccd1 vccd1 _04652_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_3_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06818_ top.DUT.register\[24\]\[17\] net644 net762 top.DUT.register\[9\]\[17\] _01956_
+ vssd1 vssd1 vccd1 vccd1 _01957_ sky130_fd_sc_hd__a221o_1
X_07798_ top.DUT.register\[13\]\[2\] net463 net459 top.DUT.register\[17\]\[2\] vssd1
+ vssd1 vccd1 vccd1 _02937_ sky130_fd_sc_hd__a22o_1
XFILLER_0_210_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09537_ _04584_ _04585_ vssd1 vssd1 vccd1 vccd1 _04587_ sky130_fd_sc_hd__nor2_1
XFILLER_0_195_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06749_ top.DUT.register\[15\]\[24\] net682 net678 top.DUT.register\[31\]\[24\] vssd1
+ vssd1 vccd1 vccd1 _01888_ sky130_fd_sc_hd__a22o_1
XFILLER_0_149_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout916_A net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout537_X net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_195_3373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_705 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09468_ top.pc\[23\] _04506_ vssd1 vssd1 vccd1 vccd1 _04522_ sky130_fd_sc_hd__nor2_1
XANTENNA__07287__A2 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10291__A1 net156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06495__B1 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08419_ _02525_ _03057_ vssd1 vssd1 vccd1 vccd1 _03550_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10637__S net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout704_X net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09399_ _04456_ _04457_ vssd1 vssd1 vccd1 vccd1 _04458_ sky130_fd_sc_hd__xnor2_1
XANTENNA__08236__A1 net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11430_ _05310_ _05312_ _05309_ vssd1 vssd1 vccd1 vccd1 _05313_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_151_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_78_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11361_ _05243_ vssd1 vssd1 vccd1 vccd1 _05244_ sky130_fd_sc_hd__inv_2
XFILLER_0_61_352 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13100_ clknet_leaf_62_clk _00692_ net1093 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[18\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_10312_ net226 net1318 net382 vssd1 vssd1 vccd1 vccd1 _00489_ sky130_fd_sc_hd__mux2_1
XANTENNA__07995__B1 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11292_ _05117_ _05181_ _05121_ vssd1 vssd1 vccd1 vccd1 _05182_ sky130_fd_sc_hd__o21bai_2
XANTENNA__09197__C1 net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_210_3598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13031_ clknet_leaf_6_clk _00623_ net944 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[16\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_10243_ net207 net1637 net390 vssd1 vssd1 vccd1 vccd1 _00422_ sky130_fd_sc_hd__mux2_1
XANTENNA__10372__S net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07747__B1 net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07247__A _02329_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10174_ net1567 net156 net605 vssd1 vssd1 vccd1 vccd1 _00373_ sky130_fd_sc_hd__mux2_1
Xfanout170 net171 vssd1 vssd1 vccd1 vccd1 net170 sky130_fd_sc_hd__buf_2
Xfanout181 _04858_ vssd1 vssd1 vccd1 vccd1 net181 sky130_fd_sc_hd__buf_1
Xfanout192 _04850_ vssd1 vssd1 vccd1 vccd1 net192 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_44_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_89_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13465__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09612__D top.a1.halfData\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11059__B1 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_201_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12815_ clknet_leaf_22_clk _00407_ net1035 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[9\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_13795_ clknet_leaf_68_clk net1232 vssd1 vssd1 vccd1 vccd1 top.pad.button_control.r_counter\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_400 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_167_660 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12746_ clknet_leaf_118_clk _00338_ net955 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[7\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07278__A2 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_154_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10547__S _04989_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12677_ clknet_leaf_33_clk _00269_ net1042 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[5\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_100_1943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11628_ _05507_ _05510_ _05497_ vssd1 vssd1 vccd1 vccd1 _05511_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_170_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_503 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11559_ _05411_ _05415_ _05430_ net249 _05407_ vssd1 vssd1 vccd1 vccd1 _05442_ sky130_fd_sc_hd__a41o_1
XTAP_TAPCELL_ROW_133_2442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold607 top.DUT.register\[18\]\[2\] vssd1 vssd1 vccd1 vccd1 net1723 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07986__B1 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold618 top.DUT.register\[13\]\[4\] vssd1 vssd1 vccd1 vccd1 net1734 sky130_fd_sc_hd__dlygate4sd3_1
Xhold629 top.DUT.register\[13\]\[14\] vssd1 vssd1 vccd1 vccd1 net1745 sky130_fd_sc_hd__dlygate4sd3_1
X_13229_ clknet_leaf_44_clk _00821_ net1063 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[22\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10282__S net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09727__B2 top.a1.dataIn\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06410__B1 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08950__A2 net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08770_ _03121_ net281 vssd1 vssd1 vccd1 vccd1 _03886_ sky130_fd_sc_hd__nand2_1
X_07721_ top.DUT.register\[24\]\[3\] net645 net760 top.DUT.register\[30\]\[3\] vssd1
+ vssd1 vccd1 vccd1 _02860_ sky130_fd_sc_hd__a22o_1
XFILLER_0_109_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07652_ top.DUT.register\[5\]\[5\] net651 _02779_ _02790_ vssd1 vssd1 vccd1 vccd1
+ _02791_ sky130_fd_sc_hd__a211o_1
XFILLER_0_149_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06603_ net808 _01741_ net438 vssd1 vssd1 vccd1 vccd1 _01742_ sky130_fd_sc_hd__o21a_1
X_07583_ _02715_ _02717_ _02719_ _02721_ vssd1 vssd1 vccd1 vccd1 _02722_ sky130_fd_sc_hd__or4_2
X_06534_ top.DUT.register\[23\]\[29\] net574 net542 top.DUT.register\[8\]\[29\] vssd1
+ vssd1 vccd1 vccd1 _01673_ sky130_fd_sc_hd__a22o_1
X_09322_ net822 _02901_ vssd1 vssd1 vccd1 vccd1 _04385_ sky130_fd_sc_hd__and2_1
XFILLER_0_75_422 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_660 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_192_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10965__B net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06465_ top.a1.instruction\[20\] top.a1.instruction\[21\] top.a1.instruction\[24\]
+ _01590_ vssd1 vssd1 vccd1 vccd1 _01604_ sky130_fd_sc_hd__or4bb_4
X_09253_ _02329_ _02365_ vssd1 vssd1 vccd1 vccd1 _04320_ sky130_fd_sc_hd__nand2_1
XANTENNA__10457__S net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout232_A _04760_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08204_ _03167_ _03182_ vssd1 vssd1 vccd1 vccd1 _03342_ sky130_fd_sc_hd__or2_4
X_09184_ top.pc\[6\] _02778_ vssd1 vssd1 vccd1 vccd1 _04255_ sky130_fd_sc_hd__or2_1
XFILLER_0_173_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06396_ top.a1.instruction\[16\] net683 _01522_ _01531_ vssd1 vssd1 vccd1 vccd1 _01535_
+ sky130_fd_sc_hd__and4_4
XFILLER_0_90_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06236__A top.ramload\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_190_3292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08135_ _02409_ net299 vssd1 vssd1 vccd1 vccd1 _03273_ sky130_fd_sc_hd__nand2_1
XANTENNA__08769__A2 _03881_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11222__B1 net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13823__1107 vssd1 vssd1 vccd1 vccd1 _13823__1107/HI net1107 sky130_fd_sc_hd__conb_1
XANTENNA__07977__B1 net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08066_ _03204_ vssd1 vssd1 vccd1 vccd1 _03205_ sky130_fd_sc_hd__inv_2
XFILLER_0_160_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09718__A1 top.a1.dataIn\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09179__C1 net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout699_A _01643_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07017_ _02155_ vssd1 vssd1 vccd1 vccd1 _02156_ sky130_fd_sc_hd__inv_2
XANTENNA__09718__B2 top.pc\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_295 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09981__S net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_164_2903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout866_A _01427_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08968_ _01916_ net692 net1130 net875 vssd1 vssd1 vccd1 vccd1 _00074_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__09282__A top.pc\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07919_ _03057_ vssd1 vssd1 vccd1 vccd1 _03058_ sky130_fd_sc_hd__inv_2
XANTENNA__08154__A0 _02678_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout654_X net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08899_ _03988_ _04008_ vssd1 vssd1 vccd1 vccd1 _04009_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_197_3402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10930_ net227 top.DUT.register\[31\]\[10\] _04972_ vssd1 vssd1 vccd1 vccd1 _01091_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_104_2010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10861_ net253 net1718 net594 vssd1 vssd1 vccd1 vccd1 _01022_ sky130_fd_sc_hd__mux2_1
X_12600_ clknet_leaf_128_clk _00192_ net918 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[3\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_13580_ clknet_leaf_123_clk net1208 net927 vssd1 vssd1 vccd1 vccd1 net102 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_66_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10792_ net146 net1455 net598 vssd1 vssd1 vccd1 vccd1 _00953_ sky130_fd_sc_hd__mux2_1
X_12531_ clknet_leaf_123_clk _00123_ net927 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[1\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_66_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10367__S net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12376__RESET_B net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12462_ clknet_leaf_123_clk _00057_ net926 vssd1 vssd1 vccd1 vccd1 top.ramstore\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_10_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07680__A2 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_482 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11413_ _05294_ _05295_ vssd1 vssd1 vccd1 vccd1 _05296_ sky130_fd_sc_hd__and2_1
XANTENNA__11213__B1 _04668_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12393_ clknet_leaf_94_clk top.ru.next_FetchedInstr\[5\] net982 vssd1 vssd1 vccd1
+ vccd1 top.a1.instruction\[5\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_34_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07968__B1 net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11344_ _05224_ _05226_ vssd1 vssd1 vccd1 vccd1 _05227_ sky130_fd_sc_hd__and2_1
XFILLER_0_104_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_2172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11198__S net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06640__B1 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11275_ top.a1.row2\[34\] _05140_ _05149_ top.a1.row1\[122\] _05165_ vssd1 vssd1
+ vccd1 vccd1 _05166_ sky130_fd_sc_hd__a221o_1
XANTENNA__12705__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13014_ clknet_leaf_13_clk _00606_ net942 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[16\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_148_Right_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10226_ net155 net2292 net395 vssd1 vssd1 vccd1 vccd1 _00406_ sky130_fd_sc_hd__mux2_1
XFILLER_0_207_826 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08932__A2 net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10157_ net2264 net220 net602 vssd1 vssd1 vccd1 vccd1 _00356_ sky130_fd_sc_hd__mux2_1
XANTENNA__10830__S net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold4 top.a1.dataInTemp\[0\] vssd1 vssd1 vccd1 vccd1 net1120 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12855__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10088_ net1604 net236 net611 vssd1 vssd1 vccd1 vccd1 _00289_ sky130_fd_sc_hd__mux2_1
XANTENNA__07499__A2 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_202_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_187_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_187_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_591 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_44_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13778_ clknet_leaf_99_clk _01349_ vssd1 vssd1 vccd1 vccd1 top.lcd.cnt_500hz\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_44_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12729_ clknet_leaf_14_clk _00321_ net959 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[7\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10277__S net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06250_ net1256 net852 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedData\[11\] sky130_fd_sc_hd__and2_1
XFILLER_0_72_447 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07671__A2 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09948__A1 net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06181_ _01412_ _01419_ vssd1 vssd1 vccd1 vccd1 _01422_ sky130_fd_sc_hd__or2_1
XFILLER_0_25_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold404 top.DUT.register\[23\]\[4\] vssd1 vssd1 vccd1 vccd1 net1520 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07423__A2 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold415 top.DUT.register\[8\]\[13\] vssd1 vssd1 vccd1 vccd1 net1531 sky130_fd_sc_hd__dlygate4sd3_1
Xhold426 top.DUT.register\[5\]\[8\] vssd1 vssd1 vccd1 vccd1 net1542 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold437 top.DUT.register\[9\]\[13\] vssd1 vssd1 vccd1 vccd1 net1553 sky130_fd_sc_hd__dlygate4sd3_1
Xhold448 top.DUT.register\[25\]\[5\] vssd1 vssd1 vccd1 vccd1 net1564 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06631__B1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold459 top.DUT.register\[17\]\[23\] vssd1 vssd1 vccd1 vccd1 net1575 sky130_fd_sc_hd__dlygate4sd3_1
X_09940_ net798 _04942_ _04943_ _04944_ vssd1 vssd1 vccd1 vccd1 _04945_ sky130_fd_sc_hd__a211o_1
XFILLER_0_0_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_232 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_115_Right_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout906 net908 vssd1 vssd1 vccd1 vccd1 net906 sky130_fd_sc_hd__buf_2
Xfanout917 net922 vssd1 vssd1 vccd1 vccd1 net917 sky130_fd_sc_hd__clkbuf_2
X_09871_ _04880_ _04881_ _04879_ vssd1 vssd1 vccd1 vccd1 _04882_ sky130_fd_sc_hd__a21oi_1
Xfanout928 net935 vssd1 vssd1 vccd1 vccd1 net928 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_55_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout939 net967 vssd1 vssd1 vccd1 vccd1 net939 sky130_fd_sc_hd__clkbuf_2
X_08822_ _03894_ _03934_ _01874_ vssd1 vssd1 vccd1 vccd1 _03935_ sky130_fd_sc_hd__a21o_1
XANTENNA__08923__A2 _04013_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10740__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1104 top.DUT.register\[22\]\[0\] vssd1 vssd1 vccd1 vccd1 net2220 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_146_2633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1115 top.DUT.register\[17\]\[6\] vssd1 vssd1 vccd1 vccd1 net2231 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1126 top.DUT.register\[1\]\[3\] vssd1 vssd1 vccd1 vccd1 net2242 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1137 top.DUT.register\[11\]\[10\] vssd1 vssd1 vccd1 vccd1 net2253 sky130_fd_sc_hd__dlygate4sd3_1
X_08753_ net883 top.pc\[22\] net694 _03869_ vssd1 vssd1 vccd1 vccd1 _03870_ sky130_fd_sc_hd__a22o_1
Xhold1148 top.DUT.register\[8\]\[11\] vssd1 vssd1 vccd1 vccd1 net2264 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1159 top.DUT.register\[16\]\[11\] vssd1 vssd1 vccd1 vccd1 net2275 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout182_A _04858_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07704_ top.DUT.register\[7\]\[4\] net518 net441 top.DUT.register\[5\]\[4\] _02842_
+ vssd1 vssd1 vccd1 vccd1 _02843_ sky130_fd_sc_hd__a221o_1
XANTENNA__08687__A1 net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08684_ _02049_ _03784_ _03076_ vssd1 vssd1 vccd1 vccd1 _03804_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_179_3132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06698__B1 net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07635_ top.a1.instruction\[25\] net789 net793 top.a1.instruction\[17\] vssd1 vssd1
+ vccd1 vccd1 _02774_ sky130_fd_sc_hd__a22oi_4
XFILLER_0_95_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1091_A net1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout447_A _01562_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08439__A1 net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07566_ top.DUT.register\[12\]\[6\] net531 net511 top.DUT.register\[24\]\[6\] vssd1
+ vssd1 vccd1 vccd1 _02705_ sky130_fd_sc_hd__a22o_1
XANTENNA__08439__B2 _03569_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_192_3321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_192_3332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09305_ net822 _02949_ vssd1 vssd1 vccd1 vccd1 _04369_ sky130_fd_sc_hd__and2_1
XFILLER_0_76_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06517_ net807 _01655_ net437 vssd1 vssd1 vccd1 vccd1 _01656_ sky130_fd_sc_hd__o21a_1
XANTENNA__11443__B1 top.a1.dataIn\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout614_A _04955_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07497_ top.DUT.register\[21\]\[14\] net657 net749 top.DUT.register\[17\]\[14\] vssd1
+ vssd1 vccd1 vccd1 _02636_ sky130_fd_sc_hd__a22o_1
XFILLER_0_180_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09976__S net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09236_ _02544_ _02547_ vssd1 vssd1 vccd1 vccd1 _04304_ sky130_fd_sc_hd__and2_1
X_06448_ net809 _01584_ vssd1 vssd1 vccd1 vccd1 _01587_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_17_Right_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_157_2795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_184 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06870__B1 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10915__S net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06379_ top.a1.instruction\[15\] top.a1.instruction\[16\] vssd1 vssd1 vccd1 vccd1
+ _01518_ sky130_fd_sc_hd__and2_1
X_09167_ _04225_ _04228_ _04226_ vssd1 vssd1 vccd1 vccd1 _04239_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_44_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_2_Left_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08118_ _03163_ _03167_ vssd1 vssd1 vccd1 vccd1 _03257_ sky130_fd_sc_hd__nor2_1
XANTENNA__08611__A1 net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07414__A2 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_0_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09098_ _04149_ _04172_ vssd1 vssd1 vccd1 vccd1 _04173_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_170_2995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout983_A net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06622__B1 net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08049_ _03177_ net433 net501 _03179_ vssd1 vssd1 vccd1 vccd1 _03188_ sky130_fd_sc_hd__a22o_1
XFILLER_0_102_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold960 top.DUT.register\[1\]\[2\] vssd1 vssd1 vccd1 vccd1 net2076 sky130_fd_sc_hd__dlygate4sd3_1
Xhold971 top.DUT.register\[8\]\[12\] vssd1 vssd1 vccd1 vccd1 net2087 sky130_fd_sc_hd__dlygate4sd3_1
Xhold982 top.DUT.register\[16\]\[24\] vssd1 vssd1 vccd1 vccd1 net2098 sky130_fd_sc_hd__dlygate4sd3_1
X_11060_ net1180 net866 net837 top.ramstore\[11\] vssd1 vssd1 vccd1 vccd1 _01171_
+ sky130_fd_sc_hd__a22o_1
Xhold993 top.DUT.register\[6\]\[10\] vssd1 vssd1 vccd1 vccd1 net2109 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout771_X net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08375__B1 _03495_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout869_X net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10011_ net140 net1913 net624 vssd1 vssd1 vccd1 vccd1 _00216_ sky130_fd_sc_hd__mux2_1
XFILLER_0_177_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10650__S net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_2091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_26_Right_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11962_ _05782_ _05806_ _05844_ vssd1 vssd1 vccd1 vccd1 _05845_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_86_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_733 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13701_ clknet_leaf_71_clk _01272_ vssd1 vssd1 vccd1 vccd1 top.lcd.lcd_rs sky130_fd_sc_hd__dfxtp_1
XFILLER_0_168_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10913_ net1711 net168 net478 vssd1 vssd1 vccd1 vccd1 _01074_ sky130_fd_sc_hd__mux2_1
X_11893_ _05774_ _05775_ vssd1 vssd1 vccd1 vccd1 _05776_ sky130_fd_sc_hd__or2_1
XFILLER_0_67_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_731 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13632_ clknet_leaf_72_clk _01219_ net1085 vssd1 vssd1 vccd1 vccd1 net59 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_211_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10844_ net1680 net200 net476 vssd1 vssd1 vccd1 vccd1 _01005_ sky130_fd_sc_hd__mux2_1
XFILLER_0_169_799 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06428__X _01567_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13563_ clknet_leaf_105_clk _01150_ net968 vssd1 vssd1 vccd1 vccd1 top.ramload\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10097__S net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_572 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10775_ net2250 net190 net484 vssd1 vssd1 vccd1 vccd1 _00936_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_35_Right_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_734 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09886__S net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12514_ clknet_leaf_86_clk _00106_ net1006 vssd1 vssd1 vccd1 vccd1 top.pc\[26\] sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_117_2201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08643__X _03765_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13494_ clknet_leaf_3_clk _01086_ net920 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[31\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07653__A2 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06861__B1 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12445_ clknet_leaf_75_clk _00041_ net1081 vssd1 vssd1 vccd1 vccd1 top.ramaddr\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10825__S net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_57_Left_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_322 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_491 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12376_ clknet_leaf_109_clk top.ru.next_FetchedData\[20\] net976 vssd1 vssd1 vccd1
+ vccd1 top.a1.dataIn\[20\] sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_130_2401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06604__A _01721_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_1897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06613__B1 net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11327_ _05206_ _05208_ _05209_ _05205_ _05204_ vssd1 vssd1 vccd1 vccd1 _05210_ sky130_fd_sc_hd__a32o_1
XFILLER_0_22_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13345__RESET_B net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11258_ top.a1.row1\[120\] _05149_ _05150_ top.a1.row1\[104\] _05147_ vssd1 vssd1
+ vccd1 vccd1 _05151_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_44_Right_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10209_ net211 net2066 net393 vssd1 vssd1 vccd1 vccd1 _00389_ sky130_fd_sc_hd__mux2_1
XANTENNA__10560__S net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11189_ net1250 net587 net473 _05101_ vssd1 vssd1 vccd1 vccd1 _01244_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_128_2363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_66_Left_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_173_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06392__A2 top.a1.instruction\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_50_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12980__RESET_B net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13822__1106 vssd1 vssd1 vccd1 vccd1 _13822__1106/HI net1106 sky130_fd_sc_hd__conb_1
XFILLER_0_82_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_wire415_A net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_141_2563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07420_ top.DUT.register\[7\]\[9\] net659 net754 top.DUT.register\[1\]\[9\] _02555_
+ vssd1 vssd1 vccd1 vccd1 _02559_ sky130_fd_sc_hd__a221o_1
XFILLER_0_187_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_175_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07892__A2 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_53_Right_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07170__A _02286_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07351_ top.DUT.register\[2\]\[8\] net560 net543 top.DUT.register\[16\]\[8\] _02489_
+ vssd1 vssd1 vccd1 vccd1 _02490_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_174_3051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_174_3062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09796__S net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06302_ _01331_ _01453_ vssd1 vssd1 vccd1 vccd1 _01459_ sky130_fd_sc_hd__and2_1
XFILLER_0_45_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07282_ _02414_ _02416_ _02419_ _02420_ vssd1 vssd1 vccd1 vccd1 _02421_ sky130_fd_sc_hd__or4_1
XFILLER_0_143_600 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07644__A2 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_75_Left_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06233_ top.ramload\[27\] net858 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedInstr\[27\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_115_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09021_ _02568_ _02800_ _02851_ _02946_ vssd1 vssd1 vccd1 vccd1 _04096_ sky130_fd_sc_hd__or4b_1
XANTENNA__06852__B1 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10735__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09809__B _04471_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06164_ net2031 vssd1 vssd1 vccd1 vccd1 _01407_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_57_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold201 top.ramaddr\[27\] vssd1 vssd1 vccd1 vccd1 net1317 sky130_fd_sc_hd__dlygate4sd3_1
Xhold212 top.DUT.register\[31\]\[2\] vssd1 vssd1 vccd1 vccd1 net1328 sky130_fd_sc_hd__dlygate4sd3_1
Xhold223 top.DUT.register\[18\]\[27\] vssd1 vssd1 vccd1 vccd1 net1339 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold234 top.a1.row1\[109\] vssd1 vssd1 vccd1 vccd1 net1350 sky130_fd_sc_hd__dlygate4sd3_1
Xhold245 top.DUT.register\[4\]\[19\] vssd1 vssd1 vccd1 vccd1 net1361 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold256 top.DUT.register\[2\]\[5\] vssd1 vssd1 vccd1 vccd1 net1372 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06233__B net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_62_Right_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold267 top.DUT.register\[15\]\[22\] vssd1 vssd1 vccd1 vccd1 net1383 sky130_fd_sc_hd__dlygate4sd3_1
Xhold278 top.DUT.register\[25\]\[30\] vssd1 vssd1 vccd1 vccd1 net1394 sky130_fd_sc_hd__dlygate4sd3_1
X_09923_ top.DUT.register\[1\]\[29\] net154 net634 vssd1 vssd1 vccd1 vccd1 _00150_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_70_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout703 _01642_ vssd1 vssd1 vccd1 vccd1 net703 sky130_fd_sc_hd__clkbuf_4
Xhold289 top.DUT.register\[11\]\[31\] vssd1 vssd1 vccd1 vccd1 net1405 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout714 _01637_ vssd1 vssd1 vccd1 vccd1 net714 sky130_fd_sc_hd__clkbuf_8
Xfanout725 _01630_ vssd1 vssd1 vccd1 vccd1 net725 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_0_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout736 net737 vssd1 vssd1 vccd1 vccd1 net736 sky130_fd_sc_hd__buf_6
XANTENNA__10470__S net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout747 _01622_ vssd1 vssd1 vccd1 vccd1 net747 sky130_fd_sc_hd__buf_4
X_09854_ _04865_ _04866_ _04860_ vssd1 vssd1 vccd1 vccd1 _04867_ sky130_fd_sc_hd__o21ai_1
XANTENNA__06520__Y _01659_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout758 _01617_ vssd1 vssd1 vccd1 vccd1 net758 sky130_fd_sc_hd__clkbuf_8
Xfanout769 _01615_ vssd1 vssd1 vccd1 vccd1 net769 sky130_fd_sc_hd__buf_4
XPHY_EDGE_ROW_84_Left_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08805_ net274 _03757_ _03918_ net285 vssd1 vssd1 vccd1 vccd1 _03919_ sky130_fd_sc_hd__a22o_1
X_09785_ _03745_ net403 net491 _04804_ vssd1 vssd1 vccd1 vccd1 _04805_ sky130_fd_sc_hd__o211a_2
XFILLER_0_147_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06997_ _02133_ _02135_ vssd1 vssd1 vccd1 vccd1 _02136_ sky130_fd_sc_hd__or2_2
XANTENNA_fanout564_A _01528_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08736_ net496 _03852_ vssd1 vssd1 vccd1 vccd1 _03853_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_1_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_72_clk_A clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout731_A _01627_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08667_ net883 top.pc\[18\] net694 _03787_ vssd1 vssd1 vccd1 vccd1 _03788_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout352_X net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_71_Right_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07618_ top.DUT.register\[26\]\[5\] net530 net447 top.DUT.register\[21\]\[5\] vssd1
+ vssd1 vccd1 vccd1 _02757_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_159_2824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_159_2835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07883__A2 net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08598_ _02614_ _03721_ vssd1 vssd1 vccd1 vccd1 _03722_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_193_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_166_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07549_ top.DUT.register\[25\]\[7\] net778 net722 top.DUT.register\[29\]\[7\] vssd1
+ vssd1 vccd1 vccd1 _02688_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_81_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_81_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_87_clk_A clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout617_X net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07096__B1 net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07635__A2 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10560_ net1595 net150 net355 vssd1 vssd1 vccd1 vccd1 _00727_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_244 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_130_clk_A clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_575 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09219_ top.pc\[8\] _02682_ vssd1 vssd1 vccd1 vccd1 _04288_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_20_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10645__S net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10491_ net1423 net158 net364 vssd1 vssd1 vccd1 vccd1 _00661_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_20_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07079__X _02218_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12230_ top.lcd.cnt_20ms\[7\] top.lcd.cnt_20ms\[6\] _06053_ vssd1 vssd1 vccd1 vccd1
+ _06069_ sky130_fd_sc_hd__and3_1
XFILLER_0_44_491 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_10_clk_A clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout986_X net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_80_Right_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_112_2120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12161_ top.a1.dataIn\[1\] _06035_ _06041_ vssd1 vssd1 vccd1 vccd1 _06044_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_112_2131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11112_ net905 net1629 net860 _05061_ vssd1 vssd1 vccd1 vccd1 _01207_ sky130_fd_sc_hd__a31o_1
X_12092_ _05970_ _05974_ vssd1 vssd1 vccd1 vccd1 _05975_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_9_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold790 top.DUT.register\[29\]\[15\] vssd1 vssd1 vccd1 vccd1 net1906 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_25_clk_A clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11043_ net23 net838 net816 net2112 vssd1 vssd1 vccd1 vccd1 _01155_ sky130_fd_sc_hd__o22a_1
XANTENNA__10380__S net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12161__A top.a1.dataIn\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_207_3548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07020__B1 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_204_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08638__X _03760_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12994_ clknet_leaf_11_clk _00586_ net951 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[15\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_98_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09470__A top.pc\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_530 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11945_ _05801_ _05826_ vssd1 vssd1 vccd1 vccd1 _05828_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_28_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08520__B1 _03645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_123_2293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08086__A _02899_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11876_ _05758_ vssd1 vssd1 vccd1 vccd1 _05759_ sky130_fd_sc_hd__inv_2
XANTENNA__07874__A2 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13615_ clknet_leaf_91_clk _01202_ net999 vssd1 vssd1 vccd1 vccd1 net41 sky130_fd_sc_hd__dfrtp_1
X_10827_ net1351 net259 net475 vssd1 vssd1 vccd1 vccd1 _00988_ sky130_fd_sc_hd__mux2_1
XANTENNA__07087__B1 net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13546_ clknet_leaf_104_clk _01133_ net972 vssd1 vssd1 vccd1 vccd1 top.ramload\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_10758_ net1394 net150 net420 vssd1 vssd1 vccd1 vccd1 _00919_ sky130_fd_sc_hd__mux2_1
XANTENNA__07626__A2 net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_1926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_1937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_290 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13477_ clknet_leaf_35_clk _01069_ net1042 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[30\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_152_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10689_ net1560 net159 net341 vssd1 vssd1 vccd1 vccd1 _00852_ sky130_fd_sc_hd__mux2_1
XANTENNA__11240__A top.lcd.nextState\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12428_ clknet_leaf_88_clk _00024_ net1001 vssd1 vssd1 vccd1 vccd1 top.ramaddr\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09379__A2 _01939_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_168_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12359_ clknet_leaf_94_clk top.ru.next_FetchedData\[3\] net982 vssd1 vssd1 vccd1
+ vccd1 top.a1.dataIn\[3\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_77_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10290__S net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06920_ _02052_ _02054_ _02056_ _02058_ vssd1 vssd1 vccd1 vccd1 _02059_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_52_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09000__A1 net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06340__Y top.lcd.lcd_en vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07011__B1 net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09932__X _04938_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06851_ top.DUT.register\[5\]\[19\] net653 net704 top.DUT.register\[3\]\[19\] _01989_
+ vssd1 vssd1 vccd1 vccd1 _01990_ sky130_fd_sc_hd__a221o_1
XANTENNA__09551__A2 _04577_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_207_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09570_ _04602_ _04617_ vssd1 vssd1 vccd1 vccd1 _04618_ sky130_fd_sc_hd__nand2_1
X_06782_ _01918_ _01919_ vssd1 vssd1 vccd1 vccd1 _01921_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_93_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08521_ _03245_ _03249_ vssd1 vssd1 vccd1 vccd1 _03648_ sky130_fd_sc_hd__and2_1
XFILLER_0_26_72 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_303 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08511__B1 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08452_ _02571_ net492 _03580_ net434 vssd1 vssd1 vccd1 vccd1 _03582_ sky130_fd_sc_hd__o22a_1
XANTENNA__07612__B _02749_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07865__A2 net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_175_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkload84_A clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07403_ top.DUT.register\[10\]\[9\] net519 net447 top.DUT.register\[21\]\[9\] _02541_
+ vssd1 vssd1 vccd1 vccd1 _02542_ sky130_fd_sc_hd__a221o_1
XFILLER_0_18_403 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08383_ net1537 net833 net803 _03515_ vssd1 vssd1 vccd1 vccd1 _00024_ sky130_fd_sc_hd__a22o_1
XFILLER_0_18_425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_60 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06228__B net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout145_A net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_268 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07334_ net823 _02472_ _01586_ vssd1 vssd1 vccd1 vccd1 _02473_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_63_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07617__A2 net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_622 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_154_2754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10465__S net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07265_ top.DUT.register\[2\]\[13\] net561 net545 top.DUT.register\[16\]\[13\] vssd1
+ vssd1 vccd1 vccd1 _02404_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout312_A net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_154 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09004_ _04069_ _04070_ _04071_ _04078_ vssd1 vssd1 vccd1 vccd1 _04079_ sky130_fd_sc_hd__or4_1
XFILLER_0_131_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_171_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06216_ net2313 net856 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedInstr\[10\] sky130_fd_sc_hd__and2_1
X_07196_ _02333_ _02334_ vssd1 vssd1 vccd1 vccd1 _02335_ sky130_fd_sc_hd__nor2_1
XFILLER_0_5_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06147_ top.a1.instruction\[6\] vssd1 vssd1 vccd1 vccd1 _01390_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_187_3253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_92_Left_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12126__A1 top.a1.dataIn\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout681_A _01547_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout500 net502 vssd1 vssd1 vccd1 vccd1 net500 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout779_A _01603_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout511 _01559_ vssd1 vssd1 vccd1 vccd1 net511 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_111_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout522 _01555_ vssd1 vssd1 vccd1 vccd1 net522 sky130_fd_sc_hd__clkbuf_8
X_09906_ net828 _04599_ _04911_ _04912_ vssd1 vssd1 vccd1 vccd1 _04914_ sky130_fd_sc_hd__o22ai_1
XTAP_TAPCELL_ROW_6_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout533 _01542_ vssd1 vssd1 vccd1 vccd1 net533 sky130_fd_sc_hd__clkbuf_8
Xfanout544 net545 vssd1 vssd1 vccd1 vccd1 net544 sky130_fd_sc_hd__clkbuf_8
Xfanout555 net558 vssd1 vssd1 vccd1 vccd1 net555 sky130_fd_sc_hd__clkbuf_8
XANTENNA__07002__B1 net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout566 _01528_ vssd1 vssd1 vccd1 vccd1 net566 sky130_fd_sc_hd__buf_4
Xfanout577 net578 vssd1 vssd1 vccd1 vccd1 net577 sky130_fd_sc_hd__buf_4
X_09837_ top.pc\[22\] _04514_ vssd1 vssd1 vccd1 vccd1 _04851_ sky130_fd_sc_hd__xnor2_1
Xfanout588 _05097_ vssd1 vssd1 vccd1 vccd1 net588 sky130_fd_sc_hd__buf_2
XANTENNA_fanout567_X net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08130__B1_N net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout599 _04965_ vssd1 vssd1 vccd1 vccd1 net599 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout946_A net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08750__B1 net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09768_ top.pc\[14\] _04386_ _04785_ vssd1 vssd1 vccd1 vccd1 _04789_ sky130_fd_sc_hd__a21o_1
X_08719_ _03795_ _03836_ net287 vssd1 vssd1 vccd1 vccd1 _03837_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_202_3478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout734_X net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09699_ _04716_ _04731_ vssd1 vssd1 vccd1 vccd1 _04732_ sky130_fd_sc_hd__or2_1
XFILLER_0_96_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11730_ _05579_ _05612_ _05575_ vssd1 vssd1 vccd1 vccd1 _05613_ sky130_fd_sc_hd__o21a_1
XFILLER_0_95_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_656 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_758 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11661_ _05493_ _05543_ vssd1 vssd1 vccd1 vccd1 _05544_ sky130_fd_sc_hd__nor2_1
XFILLER_0_126_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13400_ clknet_leaf_127_clk _00992_ net929 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[28\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_64_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10612_ net223 net2033 net347 vssd1 vssd1 vccd1 vccd1 _00777_ sky130_fd_sc_hd__mux2_1
XANTENNA__08805__A1 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11592_ _05462_ net240 _05474_ _05444_ vssd1 vssd1 vccd1 vccd1 _05475_ sky130_fd_sc_hd__a211o_1
XANTENNA__08805__B2 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13331_ clknet_leaf_120_clk _00923_ net933 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[26\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06816__B1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10543_ net1421 net209 net356 vssd1 vssd1 vccd1 vccd1 _00710_ sky130_fd_sc_hd__mux2_1
XANTENNA__10375__S net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06292__A1 net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13262_ clknet_leaf_43_clk _00854_ net1062 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[23\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_121_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10474_ net1527 net221 net361 vssd1 vssd1 vccd1 vccd1 _00644_ sky130_fd_sc_hd__mux2_1
XANTENNA__06154__A top.a1.dataIn\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12213_ _06054_ _06058_ vssd1 vssd1 vccd1 vccd1 _06059_ sky130_fd_sc_hd__nor2_2
X_13821__1105 vssd1 vssd1 vccd1 vccd1 _13821__1105/HI net1105 sky130_fd_sc_hd__conb_1
XFILLER_0_20_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_1856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13193_ clknet_leaf_54_clk _00785_ net1037 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[21\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07241__B1 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12144_ _06010_ _06023_ _06024_ vssd1 vssd1 vccd1 vccd1 _06027_ sky130_fd_sc_hd__and3_1
XFILLER_0_209_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06595__A2 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09184__B _02778_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12075_ _05920_ _05923_ _05957_ vssd1 vssd1 vccd1 vccd1 _05958_ sky130_fd_sc_hd__and3_1
X_11026_ net5 net839 net817 net2131 vssd1 vssd1 vccd1 vccd1 _01138_ sky130_fd_sc_hd__o22a_1
XANTENNA__09533__A2 top.pc\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_2__f_clk_A clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09912__B _04620_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12501__RESET_B net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12977_ clknet_leaf_116_clk _00569_ net958 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[15\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09297__A1 top.pc\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11235__A top.lcd.nextState\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_371 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11928_ _05759_ _05770_ _05786_ _05775_ vssd1 vssd1 vccd1 vccd1 _05811_ sky130_fd_sc_hd__o31a_1
XANTENNA__07847__A2 net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11859_ _05715_ _05741_ vssd1 vssd1 vccd1 vccd1 _05742_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_129_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_171_3010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_103_1985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_1996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_350 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06807__B1 net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_160_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13529_ clknet_leaf_93_clk _01116_ net998 vssd1 vssd1 vccd1 vccd1 top.a1.data\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_103_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10285__S net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07050_ top.DUT.register\[15\]\[22\] net680 net676 top.DUT.register\[31\]\[22\] vssd1
+ vssd1 vccd1 vccd1 _02189_ sky130_fd_sc_hd__a22o_1
XANTENNA__07480__B1 net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_136_2484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_149_Left_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_472 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09757__C1 _04779_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput103 net103 vssd1 vssd1 vccd1 vccd1 DAT_O[8] sky130_fd_sc_hd__buf_2
Xoutput114 net114 vssd1 vssd1 vccd1 vccd1 gpio_out[12] sky130_fd_sc_hd__buf_2
XFILLER_0_2_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07232__B1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06586__A2 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12939__CLK clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07952_ _01878_ _03090_ vssd1 vssd1 vccd1 vccd1 _03091_ sky130_fd_sc_hd__nor2_1
X_06903_ top.DUT.register\[28\]\[18\] net768 _02027_ _02041_ vssd1 vssd1 vccd1 vccd1
+ _02042_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_182_3172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11129__B net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_182_3183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07883_ top.DUT.register\[23\]\[1\] net573 net506 top.DUT.register\[27\]\[1\] vssd1
+ vssd1 vccd1 vccd1 _03022_ sky130_fd_sc_hd__a22o_1
X_09622_ net850 net843 vssd1 vssd1 vccd1 vccd1 _04667_ sky130_fd_sc_hd__nor2_2
X_06834_ _01966_ _01968_ _01970_ _01972_ vssd1 vssd1 vccd1 vccd1 _01973_ sky130_fd_sc_hd__or4_1
XPHY_EDGE_ROW_158_Left_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_179_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11619__B1 top.a1.dataIn\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09553_ top.pc\[28\] _04590_ vssd1 vssd1 vccd1 vccd1 _04602_ sky130_fd_sc_hd__or2_1
X_06765_ top.DUT.register\[10\]\[24\] net773 net709 top.DUT.register\[15\]\[24\] _01899_
+ vssd1 vssd1 vccd1 vccd1 _01904_ sky130_fd_sc_hd__a221o_1
XANTENNA__09288__A1 _02443_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_195_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout262_A _04733_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_50 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08504_ net324 _03631_ vssd1 vssd1 vccd1 vccd1 _03632_ sky130_fd_sc_hd__nand2_1
XANTENNA__07299__B1 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07838__A2 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09484_ top.pc\[23\] _04514_ _04526_ vssd1 vssd1 vccd1 vccd1 _04537_ sky130_fd_sc_hd__a21o_1
X_06696_ top.DUT.register\[6\]\[25\] net567 net515 top.DUT.register\[7\]\[25\] vssd1
+ vssd1 vccd1 vccd1 _01835_ sky130_fd_sc_hd__a22o_1
XFILLER_0_144_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08435_ _02525_ _03565_ vssd1 vssd1 vccd1 vccd1 _03566_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout527_A net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06510__A2 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08366_ net303 net333 _03326_ _03498_ vssd1 vssd1 vccd1 vccd1 _03499_ sky130_fd_sc_hd__a211o_1
X_07317_ top.DUT.register\[13\]\[12\] net774 net734 top.DUT.register\[16\]\[12\] vssd1
+ vssd1 vccd1 vccd1 _02456_ sky130_fd_sc_hd__a22o_1
XFILLER_0_73_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08297_ net305 _03247_ vssd1 vssd1 vccd1 vccd1 _03432_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout315_X net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_4_13__f_clk_A clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09984__S net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07248_ _02329_ _02385_ vssd1 vssd1 vccd1 vccd1 _02387_ sky130_fd_sc_hd__nand2_1
XFILLER_0_143_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_30_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09212__A1 net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07179_ top.DUT.register\[14\]\[10\] net583 net439 top.DUT.register\[5\]\[10\] _02317_
+ vssd1 vssd1 vccd1 vccd1 _02318_ sky130_fd_sc_hd__a221o_1
XANTENNA__10923__S net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10190_ _04712_ _04952_ net689 vssd1 vssd1 vccd1 vccd1 _04970_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_76_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06577__A2 net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_167_2945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_167_2956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout330 net332 vssd1 vssd1 vccd1 vccd1 net330 sky130_fd_sc_hd__buf_2
Xfanout341 _04993_ vssd1 vssd1 vccd1 vccd1 net341 sky130_fd_sc_hd__buf_4
Xfanout352 net353 vssd1 vssd1 vccd1 vccd1 net352 sky130_fd_sc_hd__clkbuf_8
XANTENNA__09572__X _04620_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_204_3507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout851_X net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout363 net364 vssd1 vssd1 vccd1 vccd1 net363 sky130_fd_sc_hd__buf_8
Xfanout374 _04981_ vssd1 vssd1 vccd1 vccd1 net374 sky130_fd_sc_hd__clkbuf_4
Xfanout385 _04978_ vssd1 vssd1 vccd1 vccd1 net385 sky130_fd_sc_hd__buf_6
X_12900_ clknet_leaf_38_clk _00492_ net1050 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[12\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08723__B1 _03185_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout396 _04976_ vssd1 vssd1 vccd1 vccd1 net396 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_107_2052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12831_ clknet_leaf_24_clk _00423_ net1013 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[10\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09279__A1 net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11086__A1 net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12762_ clknet_leaf_2_clk _00354_ net914 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[8\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07829__A2 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_2241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_544 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11713_ _05586_ _05587_ _05595_ vssd1 vssd1 vccd1 vccd1 _05596_ sky130_fd_sc_hd__a21boi_1
XTAP_TAPCELL_ROW_120_2252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12693_ clknet_leaf_31_clk _00285_ net1018 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[6\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_166_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11644_ _05505_ _05523_ vssd1 vssd1 vccd1 vccd1 _05527_ sky130_fd_sc_hd__xor2_1
XANTENNA__08364__A net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_182 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11575_ _05421_ net249 _05424_ vssd1 vssd1 vccd1 vccd1 _05458_ sky130_fd_sc_hd__a21bo_1
Xinput16 DAT_I[22] vssd1 vssd1 vccd1 vccd1 net16 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_92_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput27 DAT_I[3] vssd1 vssd1 vccd1 vccd1 net27 sky130_fd_sc_hd__buf_1
XFILLER_0_91_180 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput38 gpio_in[18] vssd1 vssd1 vccd1 vccd1 net38 sky130_fd_sc_hd__clkbuf_1
XANTENNA__09747__X _04771_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13314_ clknet_leaf_10_clk _00906_ net950 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[25\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_135_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10526_ net1316 net148 net358 vssd1 vssd1 vccd1 vccd1 _00695_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_770 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13245_ clknet_leaf_13_clk _00837_ net953 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[23\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_10457_ net159 net2206 net366 vssd1 vssd1 vccd1 vccd1 _00628_ sky130_fd_sc_hd__mux2_1
XANTENNA__10833__S net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08303__S net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08964__A1_N _02175_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13176_ clknet_leaf_127_clk _00768_ net929 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[21\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_10388_ net1893 net165 net376 vssd1 vssd1 vccd1 vccd1 _00563_ sky130_fd_sc_hd__mux2_1
XANTENNA__06568__A2 net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12753__RESET_B net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12127_ _06008_ _06009_ vssd1 vssd1 vccd1 vccd1 _06010_ sky130_fd_sc_hd__nand2_1
XFILLER_0_165_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12058_ _05909_ _05937_ vssd1 vssd1 vccd1 vccd1 _05941_ sky130_fd_sc_hd__xor2_2
XANTENNA__11313__A2 _05120_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11009_ net1186 _05040_ net589 vssd1 vssd1 vccd1 vccd1 _01125_ sky130_fd_sc_hd__mux2_1
XFILLER_0_177_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09361__C _04420_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_177_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_181_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06740__A2 net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_319 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06550_ top.DUT.register\[13\]\[29\] net776 net653 top.DUT.register\[5\]\[29\] vssd1
+ vssd1 vccd1 vccd1 _01689_ sky130_fd_sc_hd__a22o_1
XFILLER_0_59_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_47_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06481_ net787 _01602_ _01618_ vssd1 vssd1 vccd1 vccd1 _01620_ sky130_fd_sc_hd__and3_2
XANTENNA__09690__A1 top.a1.dataIn\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09690__B2 top.pc\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08220_ _03356_ vssd1 vssd1 vccd1 vccd1 _03357_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_138_2513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08151_ _02944_ net300 vssd1 vssd1 vccd1 vccd1 _03289_ sky130_fd_sc_hd__or2_1
XFILLER_0_43_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09442__A1 _02156_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07102_ _02234_ _02236_ _02238_ _02240_ vssd1 vssd1 vccd1 vccd1 _02241_ sky130_fd_sc_hd__or4_4
XTAP_TAPCELL_ROW_151_2713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07453__B1 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08082_ net276 _03220_ _03217_ vssd1 vssd1 vccd1 vccd1 _03221_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_31_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_99 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07033_ top.DUT.register\[26\]\[20\] net753 net748 top.DUT.register\[17\]\[20\] vssd1
+ vssd1 vccd1 vccd1 _02172_ sky130_fd_sc_hd__a22o_1
XANTENNA__10743__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_675 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_184_3201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_184_3212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11001__B2 top.a1.dataIn\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06559__A2 _01697_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08953__B1 top.ramstore\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08984_ _03832_ _03852_ _03872_ _04058_ vssd1 vssd1 vccd1 vccd1 _04059_ sky130_fd_sc_hd__and4b_1
XANTENNA__06241__B net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1017_A net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_149_2675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07935_ _03073_ vssd1 vssd1 vccd1 vccd1 _03074_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_149_2686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09552__B _04590_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07866_ top.DUT.register\[26\]\[1\] net752 net728 top.DUT.register\[18\]\[1\] vssd1
+ vssd1 vccd1 vccd1 _03005_ sky130_fd_sc_hd__a22o_1
X_09605_ _04638_ _04648_ _04649_ vssd1 vssd1 vccd1 vccd1 _04651_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_162_2875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06817_ top.DUT.register\[30\]\[17\] net759 net710 top.DUT.register\[11\]\[17\] vssd1
+ vssd1 vccd1 vccd1 _01956_ sky130_fd_sc_hd__a22o_1
XFILLER_0_211_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07797_ top.DUT.register\[28\]\[2\] net555 _02935_ vssd1 vssd1 vccd1 vccd1 _02936_
+ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout644_A _01613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_195_403 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06731__A2 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09536_ _04584_ _04585_ vssd1 vssd1 vccd1 vccd1 _04586_ sky130_fd_sc_hd__and2_1
XFILLER_0_211_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06748_ _01880_ _01882_ _01884_ _01886_ vssd1 vssd1 vccd1 vccd1 _01887_ sky130_fd_sc_hd__or4_4
XFILLER_0_210_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13820__1104 vssd1 vssd1 vccd1 vccd1 _13820__1104/HI net1104 sky130_fd_sc_hd__conb_1
XFILLER_0_66_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_195_3374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09467_ top.pc\[23\] _04506_ vssd1 vssd1 vccd1 vccd1 _04521_ sky130_fd_sc_hd__and2_1
XFILLER_0_210_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06679_ top.DUT.register\[18\]\[26\] net729 net720 top.DUT.register\[19\]\[26\] vssd1
+ vssd1 vccd1 vccd1 _01818_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout811_A net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10918__S net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08418_ net1646 net832 net803 _03549_ vssd1 vssd1 vccd1 vccd1 _00025_ sky130_fd_sc_hd__a22o_1
XFILLER_0_136_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07692__B1 net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08184__A _01678_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_175_182 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09398_ _04436_ _04439_ _04441_ vssd1 vssd1 vccd1 vccd1 _04457_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_81_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08349_ net322 _03482_ _03466_ vssd1 vssd1 vccd1 vccd1 _03483_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_80_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_129_Right_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_528 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_78_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_190_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11360_ top.a1.dataIn\[26\] _05238_ vssd1 vssd1 vccd1 vccd1 _05243_ sky130_fd_sc_hd__xor2_2
XANTENNA__07444__B1 net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_375 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout899_X net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06798__A2 net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10311_ net188 net1400 net381 vssd1 vssd1 vccd1 vccd1 _00488_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10653__S net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11291_ net879 _01381_ _05128_ _05180_ vssd1 vssd1 vccd1 vccd1 _05181_ sky130_fd_sc_hd__a31o_1
XFILLER_0_104_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_91_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13030_ clknet_leaf_40_clk _00622_ net1053 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[16\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_91_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10242_ net212 net1945 net389 vssd1 vssd1 vccd1 vccd1 _00421_ sky130_fd_sc_hd__mux2_1
XANTENNA__09736__A2 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_210_3599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08944__B1 _02973_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10173_ net2119 net160 net605 vssd1 vssd1 vccd1 vccd1 _00372_ sky130_fd_sc_hd__mux2_1
XANTENNA__07247__B _02385_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09743__A top.pc\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input38_A gpio_in[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout160 _04906_ vssd1 vssd1 vccd1 vccd1 net160 sky130_fd_sc_hd__clkbuf_2
Xfanout171 _04885_ vssd1 vssd1 vccd1 vccd1 net171 sky130_fd_sc_hd__clkbuf_2
XANTENNA__06970__A2 net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout182 _04858_ vssd1 vssd1 vccd1 vccd1 net182 sky130_fd_sc_hd__clkbuf_2
Xfanout193 _04850_ vssd1 vssd1 vccd1 vccd1 net193 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_89_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_202_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06722__A2 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12814_ clknet_leaf_43_clk _00406_ net1062 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[9\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_158_116 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13794_ clknet_leaf_68_clk _01363_ vssd1 vssd1 vccd1 vccd1 top.pad.button_control.r_counter\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_201_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_114 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12745_ clknet_leaf_21_clk _00337_ net1033 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[7\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_155_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10828__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07683__B1 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_607 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12676_ clknet_leaf_37_clk _00268_ net1051 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[5\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08094__A _02849_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_1944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11627_ _05508_ _05509_ vssd1 vssd1 vccd1 vccd1 _05510_ sky130_fd_sc_hd__nor2_1
XANTENNA__11232__B _01382_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_42_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07435__B1 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08381__X _03514_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11558_ _05415_ _05430_ net249 vssd1 vssd1 vccd1 vccd1 _05441_ sky130_fd_sc_hd__and3_1
XFILLER_0_52_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06789__A2 net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold608 top.DUT.register\[16\]\[17\] vssd1 vssd1 vccd1 vccd1 net1724 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_133_2443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10509_ net1763 net207 net358 vssd1 vssd1 vccd1 vccd1 _00678_ sky130_fd_sc_hd__mux2_1
Xhold619 top.DUT.register\[31\]\[5\] vssd1 vssd1 vccd1 vccd1 net1735 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10563__S net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11489_ _05370_ _05371_ vssd1 vssd1 vccd1 vccd1 _05372_ sky130_fd_sc_hd__nand2_1
XFILLER_0_150_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13228_ clknet_leaf_64_clk _00820_ net1093 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[22\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_176_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13159_ clknet_leaf_5_clk _00751_ net937 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[20\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06961__A2 net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07720_ top.DUT.register\[13\]\[3\] net775 net749 top.DUT.register\[17\]\[3\] vssd1
+ vssd1 vccd1 vccd1 _02859_ sky130_fd_sc_hd__a22o_1
XANTENNA__09372__B _04420_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09360__B1 _04420_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07651_ top.DUT.register\[22\]\[5\] net647 net726 top.DUT.register\[18\]\[5\] _02785_
+ vssd1 vssd1 vccd1 vccd1 _02790_ sky130_fd_sc_hd__a221o_1
XANTENNA__13722__RESET_B net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07910__A1 _02880_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06602_ _01733_ _01740_ vssd1 vssd1 vccd1 vccd1 _01741_ sky130_fd_sc_hd__nor2_1
X_07582_ top.DUT.register\[17\]\[6\] net459 net523 top.DUT.register\[11\]\[6\] _02720_
+ vssd1 vssd1 vccd1 vccd1 _02721_ sky130_fd_sc_hd__a221o_1
XFILLER_0_94_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_177_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09321_ _04380_ _04383_ vssd1 vssd1 vccd1 vccd1 _04384_ sky130_fd_sc_hd__xnor2_1
X_06533_ top.DUT.register\[1\]\[29\] net445 _01669_ _01671_ vssd1 vssd1 vccd1 vccd1
+ _01672_ sky130_fd_sc_hd__a211o_1
XANTENNA__10738__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08466__A2 net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_434 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_672 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_164_119 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09252_ _02329_ _02365_ vssd1 vssd1 vccd1 vccd1 _04319_ sky130_fd_sc_hd__or2_1
XANTENNA__07674__B1 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06464_ _01591_ _01600_ _01602_ vssd1 vssd1 vccd1 vccd1 _01603_ sky130_fd_sc_hd__and3_4
XFILLER_0_185_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08203_ _03167_ _03182_ vssd1 vssd1 vccd1 vccd1 _03341_ sky130_fd_sc_hd__nor2_1
XFILLER_0_44_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09183_ _04239_ _04242_ _04240_ vssd1 vssd1 vccd1 vccd1 _04254_ sky130_fd_sc_hd__a21o_1
X_06395_ net684 _01527_ _01533_ vssd1 vssd1 vccd1 vccd1 _01534_ sky130_fd_sc_hd__and3_1
XANTENNA__06236__B net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout225_A _04805_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08134_ _03270_ _03271_ vssd1 vssd1 vccd1 vccd1 _03272_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_190_3293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08291__X _03427_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08065_ _03196_ _03203_ net311 vssd1 vssd1 vccd1 vccd1 _03204_ sky130_fd_sc_hd__mux2_2
XANTENNA__10473__S net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07016_ _02145_ _02154_ vssd1 vssd1 vccd1 vccd1 _02155_ sky130_fd_sc_hd__nor2_4
XANTENNA__09718__A2 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout594_A _04966_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08926__B1 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_164_2904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08967_ _02131_ net691 net1279 net874 vssd1 vssd1 vccd1 vccd1 _00073_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA_fanout761_A _01617_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout382_X net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout859_A top.ru.next_iready vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07918_ _02678_ _02703_ _03056_ vssd1 vssd1 vccd1 vccd1 _03057_ sky130_fd_sc_hd__a21oi_2
XANTENNA__08179__A _01854_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08898_ net497 _03993_ _04007_ vssd1 vssd1 vccd1 vccd1 _04008_ sky130_fd_sc_hd__o21a_2
XANTENNA__08154__A1 _02498_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_197_3403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07849_ top.DUT.register\[2\]\[0\] net559 net460 top.DUT.register\[17\]\[0\] _02987_
+ vssd1 vssd1 vccd1 vccd1 _02988_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_104_2000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout647_X net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_2011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10860_ net255 net2305 net596 vssd1 vssd1 vccd1 vccd1 _01021_ sky130_fd_sc_hd__mux2_1
XANTENNA__08907__A net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_182_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09519_ net137 _04569_ vssd1 vssd1 vccd1 vccd1 _04570_ sky130_fd_sc_hd__nor2_1
XANTENNA__10648__S net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout814_X net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10791_ net1513 net142 net484 vssd1 vssd1 vccd1 vccd1 _00952_ sky130_fd_sc_hd__mux2_1
XFILLER_0_149_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_242 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12530_ clknet_leaf_25_clk _00122_ net1014 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[1\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_176_491 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12461_ clknet_leaf_106_clk _00056_ net970 vssd1 vssd1 vccd1 vccd1 top.ramstore\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_10_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11412_ top.a1.dataIn\[18\] _05254_ _05285_ vssd1 vssd1 vccd1 vccd1 _05295_ sky130_fd_sc_hd__or3b_1
XFILLER_0_136_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_191_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07417__B1 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12392_ clknet_leaf_95_clk top.ru.next_FetchedInstr\[4\] net981 vssd1 vssd1 vccd1
+ vccd1 top.a1.instruction\[4\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10383__S net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11343_ top.a1.dataIn\[22\] _05211_ _05219_ _05225_ vssd1 vssd1 vccd1 vccd1 _05226_
+ sky130_fd_sc_hd__a31o_1
XANTENNA__06433__Y _01572_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_2173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06162__A net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11274_ top.a1.row1\[114\] _05132_ _05146_ top.a1.row2\[42\] vssd1 vssd1 vccd1 vccd1
+ _05165_ sky130_fd_sc_hd__a22o_1
XFILLER_0_39_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13013_ clknet_leaf_30_clk _00605_ net1019 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[16\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_10225_ net156 net1959 net395 vssd1 vssd1 vccd1 vccd1 _00405_ sky130_fd_sc_hd__mux2_1
X_10156_ net1612 net229 net602 vssd1 vssd1 vccd1 vccd1 _00355_ sky130_fd_sc_hd__mux2_1
XFILLER_0_207_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06943__A2 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold5 top.lcd.cnt_20ms\[17\] vssd1 vssd1 vccd1 vccd1 net1121 sky130_fd_sc_hd__dlygate4sd3_1
X_10087_ net2223 net245 net612 vssd1 vssd1 vccd1 vccd1 _00288_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09342__B1 _04403_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11227__B _01382_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_510 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkload3_A clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08817__A _03909_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10558__S net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13777_ clknet_leaf_99_clk _01348_ vssd1 vssd1 vccd1 vccd1 top.lcd.cnt_500hz\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_44_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10989_ net843 _05024_ _05025_ net849 top.a1.dataIn\[6\] vssd1 vssd1 vccd1 vccd1
+ _05026_ sky130_fd_sc_hd__a32o_1
XANTENNA__11243__A top.lcd.nextState\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_480 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07656__B1 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_631 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12728_ clknet_leaf_125_clk _00320_ net924 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[7\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_787 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_154_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_154_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12659_ clknet_leaf_120_clk _00251_ net932 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[5\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_72_459 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06180_ net2138 _01419_ _01421_ net888 vssd1 vssd1 vccd1 vccd1 _00009_ sky130_fd_sc_hd__a22o_1
XANTENNA__06624__X _01763_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold405 top.DUT.register\[8\]\[21\] vssd1 vssd1 vccd1 vccd1 net1521 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10293__S net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold416 top.DUT.register\[7\]\[10\] vssd1 vssd1 vccd1 vccd1 net1532 sky130_fd_sc_hd__dlygate4sd3_1
Xhold427 top.DUT.register\[15\]\[25\] vssd1 vssd1 vccd1 vccd1 net1543 sky130_fd_sc_hd__dlygate4sd3_1
Xhold438 top.DUT.register\[27\]\[26\] vssd1 vssd1 vccd1 vccd1 net1554 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07168__A _02286_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold449 top.DUT.register\[24\]\[19\] vssd1 vssd1 vccd1 vccd1 net1565 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09870_ top.pc\[25\] _04560_ vssd1 vssd1 vccd1 vccd1 _04881_ sky130_fd_sc_hd__or2_1
Xfanout907 net908 vssd1 vssd1 vccd1 vccd1 net907 sky130_fd_sc_hd__buf_2
Xfanout918 net921 vssd1 vssd1 vccd1 vccd1 net918 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_55_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout929 net931 vssd1 vssd1 vccd1 vccd1 net929 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07187__A2 net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08821_ _01876_ _01918_ vssd1 vssd1 vccd1 vccd1 _03934_ sky130_fd_sc_hd__nor2_1
XANTENNA__09842__B1_N _04855_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1105 top.lcd.cnt_20ms\[0\] vssd1 vssd1 vccd1 vccd1 net2221 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06934__A2 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_146_2634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1116 top.DUT.register\[22\]\[6\] vssd1 vssd1 vccd1 vccd1 net2232 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1127 top.DUT.register\[27\]\[18\] vssd1 vssd1 vccd1 vccd1 net2243 sky130_fd_sc_hd__dlygate4sd3_1
X_08752_ _03853_ _03867_ _03868_ vssd1 vssd1 vccd1 vccd1 _03869_ sky130_fd_sc_hd__or3_2
Xhold1138 top.DUT.register\[2\]\[9\] vssd1 vssd1 vccd1 vccd1 net2254 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1149 top.DUT.register\[1\]\[9\] vssd1 vssd1 vccd1 vccd1 net2265 sky130_fd_sc_hd__dlygate4sd3_1
X_07703_ top.DUT.register\[12\]\[4\] net533 net529 top.DUT.register\[26\]\[4\] vssd1
+ vssd1 vccd1 vccd1 _02842_ sky130_fd_sc_hd__a22o_1
XFILLER_0_136_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_178_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08683_ _03800_ _03801_ _03802_ vssd1 vssd1 vccd1 vccd1 _03803_ sky130_fd_sc_hd__and3_1
XANTENNA__09884__A1 _04151_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout175_A _04876_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_179_3133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07634_ _02763_ _02772_ vssd1 vssd1 vccd1 vccd1 _02773_ sky130_fd_sc_hd__nor2_8
XANTENNA__07895__B1 net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_767 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08727__A net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10468__S net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07565_ _02703_ vssd1 vssd1 vccd1 vccd1 _02704_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout342_A _04992_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_192_203 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_192_3322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11153__A _04658_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09304_ _04355_ _04356_ _04353_ vssd1 vssd1 vccd1 vccd1 _04368_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_192_3333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06516_ _01646_ _01654_ vssd1 vssd1 vccd1 vccd1 _01655_ sky130_fd_sc_hd__nor2_2
XFILLER_0_146_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07647__B1 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07496_ top.DUT.register\[15\]\[14\] net708 net700 top.DUT.register\[31\]\[14\] vssd1
+ vssd1 vccd1 vccd1 _02635_ sky130_fd_sc_hd__a22o_1
XFILLER_0_152_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07111__A2 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold1192_A top.ramload\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09235_ _02497_ _02502_ _04293_ vssd1 vssd1 vccd1 vccd1 _04303_ sky130_fd_sc_hd__o21ba_1
X_06447_ net823 _01585_ vssd1 vssd1 vccd1 vccd1 _01586_ sky130_fd_sc_hd__nor2_2
XFILLER_0_173_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout607_A _04956_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_157_2796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_539 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09166_ _04236_ _04237_ vssd1 vssd1 vccd1 vccd1 _04238_ sky130_fd_sc_hd__or2_1
XANTENNA__09558__A _01722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06378_ net684 _01512_ _01516_ vssd1 vssd1 vccd1 vccd1 _01517_ sky130_fd_sc_hd__and3_1
XFILLER_0_145_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08117_ net319 _03223_ net274 _03255_ _03237_ vssd1 vssd1 vccd1 vccd1 _03256_ sky130_fd_sc_hd__a221o_1
XFILLER_0_9_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09097_ _04167_ _04169_ _04171_ vssd1 vssd1 vccd1 vccd1 _04172_ sky130_fd_sc_hd__or3_4
XFILLER_0_102_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_170_2996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09992__S net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08048_ _03160_ _03164_ vssd1 vssd1 vccd1 vccd1 _03187_ sky130_fd_sc_hd__or2_2
XFILLER_0_141_380 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold950 top.DUT.register\[9\]\[12\] vssd1 vssd1 vccd1 vccd1 net2066 sky130_fd_sc_hd__dlygate4sd3_1
Xhold961 top.DUT.register\[2\]\[29\] vssd1 vssd1 vccd1 vccd1 net2077 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout597_X net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout976_A net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold972 top.DUT.register\[4\]\[3\] vssd1 vssd1 vccd1 vccd1 net2088 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10931__S net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold983 top.DUT.register\[3\]\[4\] vssd1 vssd1 vccd1 vccd1 net2099 sky130_fd_sc_hd__dlygate4sd3_1
Xhold994 top.DUT.register\[21\]\[27\] vssd1 vssd1 vccd1 vccd1 net2110 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07178__A2 net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10010_ net148 net1910 net624 vssd1 vssd1 vccd1 vccd1 _00215_ sky130_fd_sc_hd__mux2_1
XANTENNA__07806__A _02925_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09999_ net184 net1275 net625 vssd1 vssd1 vccd1 vccd1 _00204_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout764_X net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_2092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06925__A2 net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09324__B1 _04386_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11961_ _05817_ _05818_ _05820_ vssd1 vssd1 vccd1 vccd1 _05844_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_86_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_103_Left_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13700_ clknet_leaf_73_clk _01271_ vssd1 vssd1 vccd1 vccd1 net116 sky130_fd_sc_hd__dfxtp_1
X_10912_ net1345 net172 net480 vssd1 vssd1 vccd1 vccd1 _01073_ sky130_fd_sc_hd__mux2_1
XFILLER_0_169_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07886__B1 net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_196_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11892_ _05733_ _05768_ vssd1 vssd1 vccd1 vccd1 _05775_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_168_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07350__A2 net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13631_ clknet_leaf_72_clk _01218_ net1085 vssd1 vssd1 vccd1 vccd1 net58 sky130_fd_sc_hd__dfrtp_1
X_10843_ net1590 net184 net476 vssd1 vssd1 vccd1 vccd1 _01004_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_406 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09627__A1 _04164_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10378__S net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09627__B2 _04658_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13562_ clknet_leaf_105_clk _01149_ net968 vssd1 vssd1 vccd1 vccd1 top.ramload\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_149_480 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10774_ net1216 net197 net484 vssd1 vssd1 vccd1 vccd1 _00935_ sky130_fd_sc_hd__mux2_1
XANTENNA__06157__A top.a1.dataIn\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_181_Right_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12513_ clknet_leaf_82_clk _00105_ net993 vssd1 vssd1 vccd1 vccd1 top.pc\[25\] sky130_fd_sc_hd__dfstp_2
XFILLER_0_136_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13493_ clknet_leaf_32_clk _01085_ net1044 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[31\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_2202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08850__A2 net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_23_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09468__A top.pc\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12444_ clknet_leaf_75_clk _00040_ net1083 vssd1 vssd1 vccd1 vccd1 top.ramaddr\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_152_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08372__A net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_112_Left_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12375_ clknet_leaf_109_clk top.ru.next_FetchedData\[19\] net975 vssd1 vssd1 vccd1
+ vccd1 top.a1.dataIn\[19\] sky130_fd_sc_hd__dfrtp_2
XANTENNA__08602__A2 net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_2402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08091__B net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_97_1898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11326_ top.a1.dataIn\[23\] top.a1.dataIn\[21\] top.a1.dataIn\[20\] top.a1.dataIn\[22\]
+ vssd1 vssd1 vccd1 vccd1 _05209_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_105_594 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11257_ _05129_ _01381_ top.lcd.nextState\[0\] vssd1 vssd1 vccd1 vccd1 _05150_ sky130_fd_sc_hd__and3b_2
XANTENNA__10841__S net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10208_ net221 net1639 net393 vssd1 vssd1 vccd1 vccd1 _00388_ sky130_fd_sc_hd__mux2_1
X_11188_ top.a1.data\[9\] net783 _05033_ vssd1 vssd1 vccd1 vccd1 _05101_ sky130_fd_sc_hd__o21a_1
XFILLER_0_206_112 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06916__A2 net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10139_ net165 net2207 net610 vssd1 vssd1 vccd1 vccd1 _00339_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_128_2364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09490__X _04543_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_121_Left_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_206_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_50_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09866__A1 top.a1.instruction\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_203_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_199_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07877__B1 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07341__A2 net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_141_2564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07451__A _02580_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire408_A net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13829_ net1113 vssd1 vssd1 vccd1 vccd1 gpio_out[28] sky130_fd_sc_hd__buf_2
XANTENNA__10288__S net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07629__B1 net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07350_ top.DUT.register\[22\]\[8\] net578 net563 top.DUT.register\[20\]\[8\] vssd1
+ vssd1 vccd1 vccd1 _02489_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_174_3052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_174_3063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06301_ _01448_ _01457_ _01458_ _01449_ _01455_ vssd1 vssd1 vccd1 vccd1 _00000_ sky130_fd_sc_hd__a32o_1
XFILLER_0_155_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07281_ top.DUT.register\[25\]\[13\] net780 net645 top.DUT.register\[24\]\[13\] _02417_
+ vssd1 vssd1 vccd1 vccd1 _02420_ sky130_fd_sc_hd__a221o_1
XFILLER_0_5_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09020_ _01658_ _03144_ _03411_ vssd1 vssd1 vccd1 vccd1 _04095_ sky130_fd_sc_hd__or3_1
X_06232_ top.ramload\[26\] net858 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedInstr\[26\]
+ sky130_fd_sc_hd__and2_1
XANTENNA__11701__A top.a1.dataIn\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_130_Left_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11189__B1 net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06163_ top.pc\[2\] vssd1 vssd1 vccd1 vccd1 _01406_ sky130_fd_sc_hd__inv_2
XFILLER_0_142_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_57_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold202 top.DUT.register\[12\]\[16\] vssd1 vssd1 vccd1 vccd1 net1318 sky130_fd_sc_hd__dlygate4sd3_1
Xhold213 top.DUT.register\[26\]\[8\] vssd1 vssd1 vccd1 vccd1 net1329 sky130_fd_sc_hd__dlygate4sd3_1
Xhold224 top.DUT.register\[23\]\[22\] vssd1 vssd1 vccd1 vccd1 net1340 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07801__B1 net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold235 top.DUT.register\[28\]\[3\] vssd1 vssd1 vccd1 vccd1 net1351 sky130_fd_sc_hd__dlygate4sd3_1
Xhold246 top.a1.row2\[10\] vssd1 vssd1 vccd1 vccd1 net1362 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_531 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold257 top.DUT.register\[4\]\[28\] vssd1 vssd1 vccd1 vccd1 net1373 sky130_fd_sc_hd__dlygate4sd3_1
Xhold268 top.DUT.register\[13\]\[5\] vssd1 vssd1 vccd1 vccd1 net1384 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10751__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold279 top.DUT.register\[4\]\[14\] vssd1 vssd1 vccd1 vccd1 net1395 sky130_fd_sc_hd__dlygate4sd3_1
X_09922_ net489 _04917_ _04928_ vssd1 vssd1 vccd1 vccd1 _04929_ sky130_fd_sc_hd__and3_4
XANTENNA__06801__Y _01940_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout704 _01642_ vssd1 vssd1 vccd1 vccd1 net704 sky130_fd_sc_hd__clkbuf_8
Xfanout715 _01637_ vssd1 vssd1 vccd1 vccd1 net715 sky130_fd_sc_hd__buf_4
Xfanout726 _01628_ vssd1 vssd1 vccd1 vccd1 net726 sky130_fd_sc_hd__clkbuf_8
Xfanout737 _01626_ vssd1 vssd1 vccd1 vccd1 net737 sky130_fd_sc_hd__buf_4
X_09853_ _04861_ _04863_ _04864_ _04151_ vssd1 vssd1 vccd1 vccd1 _04866_ sky130_fd_sc_hd__a31o_1
Xfanout748 net749 vssd1 vssd1 vccd1 vccd1 net748 sky130_fd_sc_hd__buf_4
XANTENNA_fanout292_A net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06907__A2 _02045_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout759 _01617_ vssd1 vssd1 vccd1 vccd1 net759 sky130_fd_sc_hd__buf_2
X_08804_ _03837_ _03917_ net310 vssd1 vssd1 vccd1 vccd1 _03918_ sky130_fd_sc_hd__mux2_1
X_09784_ net798 _04800_ _04801_ _04803_ vssd1 vssd1 vccd1 vccd1 _04804_ sky130_fd_sc_hd__a211o_1
X_06996_ _02112_ _02132_ vssd1 vssd1 vccd1 vccd1 _02135_ sky130_fd_sc_hd__and2_1
XANTENNA__07580__A2 net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_198_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08735_ _02222_ _03851_ vssd1 vssd1 vccd1 vccd1 _03852_ sky130_fd_sc_hd__xor2_1
XANTENNA_fanout557_A net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08666_ _03782_ _03786_ vssd1 vssd1 vccd1 vccd1 _03787_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_1_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07868__B1 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07617_ top.DUT.register\[14\]\[5\] net584 net555 top.DUT.register\[28\]\[5\] _02755_
+ vssd1 vssd1 vccd1 vccd1 _02756_ sky130_fd_sc_hd__a221o_1
XFILLER_0_95_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10198__S net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09609__A1 net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08597_ _02654_ _03701_ vssd1 vssd1 vccd1 vccd1 _03721_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout345_X net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_159_2825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout724_A _01630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_159_2836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1087_X net1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09987__S net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07548_ top.DUT.register\[15\]\[7\] net706 net698 top.DUT.register\[31\]\[7\] vssd1
+ vssd1 vccd1 vccd1 _02687_ sky130_fd_sc_hd__a22o_1
XFILLER_0_48_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08744__X _03861_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06408__C _01546_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10926__S net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout512_X net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07479_ top.DUT.register\[14\]\[14\] net585 net462 top.DUT.register\[17\]\[14\] _02617_
+ vssd1 vssd1 vccd1 vccd1 _02618_ sky130_fd_sc_hd__a221o_1
XFILLER_0_146_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_256 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09218_ top.pc\[7\] _02729_ _04274_ vssd1 vssd1 vccd1 vccd1 _04287_ sky130_fd_sc_hd__a21bo_1
X_10490_ net1982 net161 net364 vssd1 vssd1 vccd1 vccd1 _00660_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_20_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_347 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09149_ top.pc\[2\] top.pc\[3\] top.pc\[4\] vssd1 vssd1 vccd1 vccd1 _04222_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_32_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09242__C1 net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07399__A2 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08596__A1 net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08596__B2 net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12160_ _06035_ _06041_ top.a1.dataIn\[1\] vssd1 vssd1 vccd1 vccd1 _06043_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_112_2121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_112_2132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11111_ net46 net864 vssd1 vssd1 vccd1 vccd1 _05061_ sky130_fd_sc_hd__and2_1
X_12091_ _05965_ _05972_ vssd1 vssd1 vccd1 vccd1 _05974_ sky130_fd_sc_hd__nand2_1
Xhold780 top.DUT.register\[14\]\[25\] vssd1 vssd1 vccd1 vccd1 net1896 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08348__A1 net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold791 top.DUT.register\[19\]\[7\] vssd1 vssd1 vccd1 vccd1 net1907 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_6_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11042_ net22 net839 net817 net2136 vssd1 vssd1 vccd1 vccd1 _01154_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_207_3549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07571__A2 net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input20_A DAT_I[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12993_ clknet_leaf_18_clk _00585_ net1030 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[15\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_203_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09470__B _04514_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11944_ _05801_ _05826_ vssd1 vssd1 vccd1 vccd1 _05827_ sky130_fd_sc_hd__nand2_1
XFILLER_0_169_542 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07323__A2 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08520__B2 net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11875_ _05740_ _05748_ _05757_ _05742_ vssd1 vssd1 vccd1 vccd1 _05758_ sky130_fd_sc_hd__a22oi_4
XANTENNA__06531__B1 net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_123_2294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_211_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12707__RESET_B net1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10826_ net1769 net265 net474 vssd1 vssd1 vccd1 vccd1 _00987_ sky130_fd_sc_hd__mux2_1
X_13614_ clknet_leaf_91_clk _01201_ net999 vssd1 vssd1 vccd1 vccd1 net71 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_184_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_236 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_184_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10757_ net2019 net153 net420 vssd1 vssd1 vccd1 vccd1 _00918_ sky130_fd_sc_hd__mux2_1
XFILLER_0_165_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13545_ clknet_leaf_102_clk _01132_ net981 vssd1 vssd1 vccd1 vccd1 top.ramload\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10836__S net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_99_1927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_1938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13476_ clknet_leaf_37_clk _01068_ net1052 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[30\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10688_ net1749 net165 net341 vssd1 vssd1 vccd1 vccd1 _00851_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_140_604 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12427_ clknet_leaf_87_clk _00023_ net1004 vssd1 vssd1 vccd1 vccd1 top.ramaddr\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_112_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08587__A1 net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_168_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12358_ clknet_leaf_103_clk top.ru.next_FetchedData\[2\] net981 vssd1 vssd1 vccd1
+ vccd1 top.a1.dataIn\[2\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__08830__A _03370_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06598__B1 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11309_ net1209 net814 _05195_ net1084 vssd1 vssd1 vccd1 vccd1 _01270_ sky130_fd_sc_hd__o211a_1
XANTENNA__10571__S net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12289_ _06104_ net687 _06103_ vssd1 vssd1 vccd1 vccd1 _01347_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_52_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11239__Y _05132_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_184_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06850_ top.DUT.register\[28\]\[19\] net768 net716 top.DUT.register\[27\]\[19\] vssd1
+ vssd1 vccd1 vccd1 _01989_ sky130_fd_sc_hd__a22o_1
XANTENNA__09083__D top.a1.instruction\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06781_ _01918_ _01919_ vssd1 vssd1 vccd1 vccd1 _01920_ sky130_fd_sc_hd__and2b_1
XANTENNA__06770__B1 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11255__X _05148_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08520_ _02476_ net494 _03645_ net428 _03646_ vssd1 vssd1 vccd1 vccd1 _03647_ sky130_fd_sc_hd__a221o_1
XFILLER_0_77_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08511__A1 net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_203_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_194_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08511__B2 _03638_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08451_ _02568_ net431 _03187_ _02570_ vssd1 vssd1 vccd1 vccd1 _03581_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__06522__B1 net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07402_ top.DUT.register\[20\]\[9\] net563 net547 top.DUT.register\[18\]\[9\] vssd1
+ vssd1 vccd1 vccd1 _02541_ sky130_fd_sc_hd__a22o_1
XFILLER_0_9_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08382_ net886 top.pc\[6\] net697 _03514_ vssd1 vssd1 vccd1 vccd1 _03515_ sky130_fd_sc_hd__a22o_1
XFILLER_0_92_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_175_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_72 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07333_ _02463_ _02466_ _02471_ vssd1 vssd1 vccd1 vccd1 _02472_ sky130_fd_sc_hd__or3_4
XFILLER_0_46_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10746__S net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_124_clk clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_124_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_63_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08724__B net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout138_A net139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07264_ top.DUT.register\[12\]\[13\] net533 net458 top.DUT.register\[25\]\[13\] _02402_
+ vssd1 vssd1 vccd1 vccd1 _02403_ sky130_fd_sc_hd__a221o_1
XFILLER_0_155_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_154_2755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09003_ _04077_ _03902_ _04072_ vssd1 vssd1 vccd1 vccd1 _04078_ sky130_fd_sc_hd__or3b_1
XFILLER_0_115_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06215_ top.ramload\[9\] net856 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedInstr\[9\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_54_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07195_ _01389_ _01500_ vssd1 vssd1 vccd1 vccd1 _02334_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout305_A net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06244__B net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1047_A net1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11177__A3 net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09775__B1 net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06146_ top.a1.instruction\[5\] vssd1 vssd1 vccd1 vccd1 _01389_ sky130_fd_sc_hd__inv_2
XFILLER_0_41_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06589__B1 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_187_3254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10481__S net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout501 net502 vssd1 vssd1 vccd1 vccd1 net501 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_6_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09905_ top.a1.instruction\[28\] net487 net402 top.a1.dataIn\[28\] net398 vssd1 vssd1
+ vccd1 vccd1 _04913_ sky130_fd_sc_hd__a221o_1
Xfanout512 _01559_ vssd1 vssd1 vccd1 vccd1 net512 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06260__A top.ramload\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout523 _01554_ vssd1 vssd1 vccd1 vccd1 net523 sky130_fd_sc_hd__clkbuf_8
Xfanout534 _01542_ vssd1 vssd1 vccd1 vccd1 net534 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_6_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout295_X net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout545 net546 vssd1 vssd1 vccd1 vccd1 net545 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout674_A _01597_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout556 net558 vssd1 vssd1 vccd1 vccd1 net556 sky130_fd_sc_hd__clkbuf_8
X_09836_ net2249 net195 net633 vssd1 vssd1 vccd1 vccd1 _00142_ sky130_fd_sc_hd__mux2_1
Xfanout567 _01525_ vssd1 vssd1 vccd1 vccd1 net567 sky130_fd_sc_hd__clkbuf_8
Xfanout578 _01517_ vssd1 vssd1 vccd1 vccd1 net578 sky130_fd_sc_hd__clkbuf_8
Xfanout589 _05003_ vssd1 vssd1 vccd1 vccd1 net589 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07553__A2 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08750__B2 _03854_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout841_A net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06979_ top.DUT.register\[15\]\[23\] net708 net700 top.DUT.register\[31\]\[23\] vssd1
+ vssd1 vccd1 vccd1 _02118_ sky130_fd_sc_hd__a22o_1
X_09767_ net1429 net198 net633 vssd1 vssd1 vccd1 vccd1 _00135_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout462_X net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06761__B1 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout939_A net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08718_ _03303_ _03308_ vssd1 vssd1 vccd1 vccd1 _03836_ sky130_fd_sc_hd__nand2_1
X_09698_ top.a1.dataIn\[3\] _01489_ net798 top.pc\[3\] _04730_ vssd1 vssd1 vccd1 vccd1
+ _04731_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_202_3479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07305__A2 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08649_ _01962_ _02049_ _03768_ vssd1 vssd1 vccd1 vccd1 _03770_ sky130_fd_sc_hd__or3_1
XFILLER_0_68_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06513__B1 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_25_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout727_X net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11660_ _05507_ _05510_ _05515_ _05496_ vssd1 vssd1 vccd1 vccd1 _05543_ sky130_fd_sc_hd__a211o_1
XFILLER_0_95_189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10611_ net188 net1618 net347 vssd1 vssd1 vccd1 vccd1 _00776_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10656__S net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11591_ _05472_ _05473_ vssd1 vssd1 vccd1 vccd1 _05474_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_115_clk clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_115_clk
+ sky130_fd_sc_hd__clkbuf_8
X_13330_ clknet_leaf_31_clk _00922_ net1021 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[26\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_10542_ net1647 net212 _04989_ vssd1 vssd1 vccd1 vccd1 _00709_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13261_ clknet_leaf_42_clk _00853_ net1064 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[23\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06292__A2 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10473_ net1493 net229 net361 vssd1 vssd1 vccd1 vccd1 _00643_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12212_ _06055_ _06056_ _06057_ vssd1 vssd1 vccd1 vccd1 _06058_ sky130_fd_sc_hd__or3_1
XANTENNA__09766__B1 net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13192_ clknet_leaf_8_clk _00784_ net1009 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[21\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_121_136 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08650__A _02049_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_1857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12143_ _06023_ _06024_ _06010_ vssd1 vssd1 vccd1 vccd1 _06026_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10391__S net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07792__A2 net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12074_ _05952_ _05956_ _05931_ vssd1 vssd1 vccd1 vccd1 _05957_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_47_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06170__A top.a1.halfData\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11025_ net4 net838 net816 net1256 vssd1 vssd1 vccd1 vccd1 _01137_ sky130_fd_sc_hd__o22a_1
XANTENNA__08741__A1 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07544__A2 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06752__B1 net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12976_ clknet_leaf_29_clk _00568_ net1017 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[14\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_169_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11927_ _05759_ _05770_ _05775_ _05786_ vssd1 vssd1 vccd1 vccd1 _05810_ sky130_fd_sc_hd__nor4_1
XFILLER_0_169_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11858_ _05705_ _05710_ _05711_ _05719_ vssd1 vssd1 vccd1 vccd1 _05741_ sky130_fd_sc_hd__o31a_1
XFILLER_0_157_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_171_3011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_106_clk clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_106_clk
+ sky130_fd_sc_hd__clkbuf_8
X_10809_ net216 net2212 net599 vssd1 vssd1 vccd1 vccd1 _00970_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_103_1986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10566__S net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11789_ _05659_ _05671_ vssd1 vssd1 vccd1 vccd1 _05672_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_103_1997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13528_ clknet_leaf_92_clk _01115_ net998 vssd1 vssd1 vccd1 vccd1 top.a1.data\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_179_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13459_ clknet_leaf_123_clk _01051_ net927 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[30\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_136_2485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09757__B1 net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput104 net104 vssd1 vssd1 vccd1 vccd1 DAT_O[9] sky130_fd_sc_hd__buf_2
XFILLER_0_2_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput115 net115 vssd1 vssd1 vccd1 vccd1 gpio_out[13] sky130_fd_sc_hd__buf_2
XANTENNA_clkbuf_leaf_71_clk_A clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07951_ _01920_ _03088_ _03089_ vssd1 vssd1 vccd1 vccd1 _03090_ sky130_fd_sc_hd__o21a_1
X_06902_ top.DUT.register\[13\]\[18\] net775 _02040_ vssd1 vssd1 vccd1 vccd1 _02041_
+ sky130_fd_sc_hd__a21o_1
X_07882_ net295 vssd1 vssd1 vccd1 vccd1 _03021_ sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_86_clk_A clknet_4_6__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_182_3173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07535__A2 net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06833_ top.DUT.register\[24\]\[19\] net513 net454 top.DUT.register\[29\]\[19\] _01971_
+ vssd1 vssd1 vccd1 vccd1 _01972_ sky130_fd_sc_hd__a221o_1
X_09621_ top.a1.state\[0\] top.a1.state\[2\] vssd1 vssd1 vccd1 vccd1 _04666_ sky130_fd_sc_hd__nor2_1
XFILLER_0_37_94 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06743__B1 net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09552_ top.pc\[28\] _04590_ vssd1 vssd1 vccd1 vccd1 _04601_ sky130_fd_sc_hd__nand2_1
X_06764_ top.DUT.register\[7\]\[24\] net660 net641 top.DUT.register\[8\]\[24\] vssd1
+ vssd1 vccd1 vccd1 _01903_ sky130_fd_sc_hd__a22o_1
XANTENNA__09288__A2 _02452_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08503_ _03420_ _03630_ net297 vssd1 vssd1 vccd1 vccd1 _03631_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_65_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09483_ net137 _04535_ vssd1 vssd1 vccd1 vccd1 _04536_ sky130_fd_sc_hd__nor2_1
XFILLER_0_144_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_148_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08496__B1 net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06695_ _01833_ vssd1 vssd1 vccd1 vccd1 _01834_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout255_A _04737_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06239__B net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_180 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08434_ _03519_ _03521_ _03517_ vssd1 vssd1 vccd1 vccd1 _03565_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_53_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08294__X _03430_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10984__B net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08365_ net302 _03369_ vssd1 vssd1 vccd1 vccd1 _03498_ sky130_fd_sc_hd__nor2_2
XFILLER_0_19_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10476__S net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_24_clk_A clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07316_ top.DUT.register\[1\]\[12\] net754 net718 top.DUT.register\[19\]\[12\] vssd1
+ vssd1 vccd1 vccd1 _02455_ sky130_fd_sc_hd__a22o_1
XFILLER_0_160_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08296_ net1291 net832 net802 _03431_ vssd1 vssd1 vccd1 vccd1 _00021_ sky130_fd_sc_hd__a22o_1
XANTENNA__07471__A1 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07247_ _02329_ _02385_ vssd1 vssd1 vccd1 vccd1 _02386_ sky130_fd_sc_hd__nor2_1
XFILLER_0_5_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_30_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_39_clk_A clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07178_ top.DUT.register\[17\]\[10\] net459 net455 top.DUT.register\[25\]\[10\] vssd1
+ vssd1 vccd1 vccd1 _02317_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout889_A net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07774__A2 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08971__B2 net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout320 _02830_ vssd1 vssd1 vccd1 vccd1 net320 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_167_2946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_167_2957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06982__B1 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout677_X net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout331 net332 vssd1 vssd1 vccd1 vccd1 net331 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout342 _04992_ vssd1 vssd1 vccd1 vccd1 net342 sky130_fd_sc_hd__buf_8
Xfanout353 _04990_ vssd1 vssd1 vccd1 vccd1 net353 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_204_3508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08469__X _03598_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout364 _04986_ vssd1 vssd1 vccd1 vccd1 net364 sky130_fd_sc_hd__clkbuf_8
Xfanout375 _04981_ vssd1 vssd1 vccd1 vccd1 net375 sky130_fd_sc_hd__buf_6
XANTENNA__07526__A2 net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout386 _04978_ vssd1 vssd1 vccd1 vccd1 net386 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07814__A _02952_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout397 _04753_ vssd1 vssd1 vccd1 vccd1 net397 sky130_fd_sc_hd__buf_2
X_09819_ top.pc\[20\] _04487_ vssd1 vssd1 vccd1 vccd1 _04835_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_107_2053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12830_ clknet_leaf_18_clk _00422_ net1028 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[10\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_158_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12761_ clknet_leaf_14_clk _00353_ net959 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[8\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_201_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_120_2242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11712_ _05593_ _05594_ _05556_ _05582_ vssd1 vssd1 vccd1 vccd1 _05595_ sky130_fd_sc_hd__o2bb2a_2
XTAP_TAPCELL_ROW_120_2253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12692_ clknet_leaf_79_clk _00284_ net1072 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[6\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_139_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_139_578 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11643_ top.a1.dataIn\[11\] _05523_ _05524_ vssd1 vssd1 vccd1 vccd1 _05526_ sky130_fd_sc_hd__or3_1
XFILLER_0_65_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10386__S net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_194 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11574_ _05424_ net249 _05421_ vssd1 vssd1 vccd1 vccd1 _05457_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_181_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput17 DAT_I[23] vssd1 vssd1 vccd1 vccd1 net17 sky130_fd_sc_hd__buf_1
Xinput28 DAT_I[4] vssd1 vssd1 vccd1 vccd1 net28 sky130_fd_sc_hd__buf_1
X_10525_ net1617 net152 net359 vssd1 vssd1 vccd1 vccd1 _00694_ sky130_fd_sc_hd__mux2_1
Xinput39 nrst vssd1 vssd1 vccd1 vccd1 net39 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_91_192 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13313_ clknet_leaf_16_clk _00905_ net963 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[25\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_150_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13244_ clknet_leaf_129_clk _00836_ net910 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[23\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09739__B1 _04752_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09476__A _01585_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10456_ net167 net1834 net366 vssd1 vssd1 vccd1 vccd1 _00627_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10349__A1 _04841_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13175_ clknet_leaf_2_clk _00767_ net918 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[21\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12563__CLK clknet_leaf_120_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10387_ net1896 net168 net373 vssd1 vssd1 vccd1 vccd1 _00562_ sky130_fd_sc_hd__mux2_1
X_12126_ top.a1.dataIn\[2\] _06004_ _06000_ vssd1 vssd1 vccd1 vccd1 _06009_ sky130_fd_sc_hd__o21ai_1
XANTENNA__08962__B2 net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12403__Q top.a1.instruction\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12057_ _05938_ _05939_ vssd1 vssd1 vccd1 vccd1 _05940_ sky130_fd_sc_hd__nor2_1
XFILLER_0_74_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11008_ net843 _05038_ _05039_ net849 top.a1.dataIn\[11\] vssd1 vssd1 vccd1 vccd1
+ _05040_ sky130_fd_sc_hd__a32o_1
XANTENNA__11313__A3 _05148_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06725__B1 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_204_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_204_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12959_ clknet_leaf_24_clk _00551_ net1015 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[14\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_176_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06480_ _01598_ _01601_ vssd1 vssd1 vccd1 vccd1 _01619_ sky130_fd_sc_hd__nor2_4
XTAP_TAPCELL_ROW_47_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07150__B1 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_185_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09690__A2 _01489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_2514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10296__S net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08150_ net300 _03040_ vssd1 vssd1 vccd1 vccd1 _03288_ sky130_fd_sc_hd__and2_1
XFILLER_0_43_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_60_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09442__A2 _04487_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07101_ top.DUT.register\[14\]\[16\] net584 net532 top.DUT.register\[12\]\[16\] _02239_
+ vssd1 vssd1 vccd1 vccd1 _02240_ sky130_fd_sc_hd__a221o_1
X_08081_ _03218_ _03219_ vssd1 vssd1 vccd1 vccd1 _03220_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_151_2714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12906__CLK clknet_leaf_120_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07032_ top.DUT.register\[5\]\[20\] net654 net756 top.DUT.register\[1\]\[20\] _02170_
+ vssd1 vssd1 vccd1 vccd1 _02171_ sky130_fd_sc_hd__a221o_1
XFILLER_0_140_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_141_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_184_3202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_184_3213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07756__A2 net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08953__B2 net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08983_ _03771_ _03790_ _03812_ _04057_ vssd1 vssd1 vccd1 vccd1 _04058_ sky130_fd_sc_hd__and4b_1
XANTENNA__06964__B1 net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07934_ _02614_ _03072_ _03070_ _03059_ vssd1 vssd1 vccd1 vccd1 _03073_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_149_2676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_149_2687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08705__A1 net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07508__A2 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08705__B2 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_208_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07865_ top.DUT.register\[24\]\[1\] net645 net741 top.DUT.register\[12\]\[1\] _03003_
+ vssd1 vssd1 vccd1 vccd1 _03004_ sky130_fd_sc_hd__a221o_1
XANTENNA__06716__B1 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout372_A _04983_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12463__RESET_B net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold1020_A top.ramload\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09604_ _04638_ _04648_ _04649_ vssd1 vssd1 vccd1 vccd1 _04650_ sky130_fd_sc_hd__and3_1
X_06816_ top.DUT.register\[28\]\[17\] net769 net723 top.DUT.register\[29\]\[17\] vssd1
+ vssd1 vccd1 vccd1 _01955_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_162_2876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07796_ top.DUT.register\[15\]\[2\] net679 net675 top.DUT.register\[31\]\[2\] vssd1
+ vssd1 vccd1 vccd1 _02935_ sky130_fd_sc_hd__a22o_1
XFILLER_0_211_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09535_ _04571_ _04572_ _04573_ vssd1 vssd1 vccd1 vccd1 _04585_ sky130_fd_sc_hd__o21a_1
X_06747_ top.DUT.register\[30\]\[24\] net581 net544 top.DUT.register\[16\]\[24\] _01885_
+ vssd1 vssd1 vccd1 vccd1 _01886_ sky130_fd_sc_hd__a221o_1
XFILLER_0_211_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout637_A _01629_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09466_ net901 top.pc\[22\] _04520_ net891 vssd1 vssd1 vccd1 vccd1 _00102_ sky130_fd_sc_hd__o211a_1
XFILLER_0_148_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_195_3364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06678_ top.DUT.register\[20\]\[26\] net666 net740 top.DUT.register\[12\]\[26\] _01816_
+ vssd1 vssd1 vccd1 vccd1 _01817_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_195_3375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07141__B1 net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08417_ net885 top.pc\[7\] net697 _03548_ vssd1 vssd1 vccd1 vccd1 _03549_ sky130_fd_sc_hd__a22o_1
XANTENNA__06495__A2 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09397_ _04454_ _04455_ vssd1 vssd1 vccd1 vccd1 _04456_ sky130_fd_sc_hd__nand2_1
XFILLER_0_148_386 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_340 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout425_X net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_175_194 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09995__S net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08348_ net297 _03481_ _03469_ vssd1 vssd1 vccd1 vccd1 _03482_ sky130_fd_sc_hd__o21a_1
XFILLER_0_191_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08752__X _03869_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10934__S net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08279_ _03187_ _03412_ vssd1 vssd1 vccd1 vccd1 _03415_ sky130_fd_sc_hd__nor2_1
XFILLER_0_34_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_719 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10310_ net196 net1726 net382 vssd1 vssd1 vccd1 vccd1 _00487_ sky130_fd_sc_hd__mux2_1
XANTENNA__07809__A top.a1.instruction\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09296__A top.pc\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07995__A2 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11290_ net882 _05128_ _05136_ _05179_ _05122_ vssd1 vssd1 vccd1 vccd1 _05180_ sky130_fd_sc_hd__a2111o_1
XANTENNA__09197__A1 net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10241_ net220 net2185 net389 vssd1 vssd1 vccd1 vccd1 _00420_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_91_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_210_3589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07747__A2 net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08944__B2 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10172_ net1977 net165 net605 vssd1 vssd1 vccd1 vccd1 _00371_ sky130_fd_sc_hd__mux2_1
XANTENNA__06955__B1 net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09743__B _04172_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout150 _04938_ vssd1 vssd1 vccd1 vccd1 net150 sky130_fd_sc_hd__clkbuf_2
Xfanout161 _04906_ vssd1 vssd1 vccd1 vccd1 net161 sky130_fd_sc_hd__buf_2
Xfanout172 _04876_ vssd1 vssd1 vccd1 vccd1 net172 sky130_fd_sc_hd__buf_2
Xfanout183 _04858_ vssd1 vssd1 vccd1 vccd1 net183 sky130_fd_sc_hd__buf_1
Xfanout194 _04850_ vssd1 vssd1 vccd1 vccd1 net194 sky130_fd_sc_hd__buf_2
XANTENNA__06707__B1 net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11700__B1 top.a1.dataIn\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_231 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07380__B1 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12813_ clknet_leaf_50_clk _00405_ net1057 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[9\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11059__A2 net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13793_ clknet_leaf_68_clk _01362_ vssd1 vssd1 vccd1 vccd1 top.pad.button_control.r_counter\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_158_128 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09121__A1 _02904_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12744_ clknet_leaf_7_clk _00336_ net946 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[7\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_177_Left_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07132__B1 net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06486__A2 top.a1.instruction\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12675_ clknet_leaf_60_clk _00267_ net1089 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[5\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_619 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06166__Y _00016_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_660 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_1945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_13_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11626_ _05447_ _05499_ vssd1 vssd1 vccd1 vccd1 _05509_ sky130_fd_sc_hd__xnor2_2
XANTENNA__11232__C _05123_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08632__B1 net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10844__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11557_ _05430_ net249 vssd1 vssd1 vccd1 vccd1 _05440_ sky130_fd_sc_hd__nand2_1
XFILLER_0_69_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_283 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07986__A2 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_2444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10508_ net1791 net211 net357 vssd1 vssd1 vccd1 vccd1 _00677_ sky130_fd_sc_hd__mux2_1
Xhold609 top.DUT.register\[3\]\[12\] vssd1 vssd1 vccd1 vccd1 net1725 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07719__A _02857_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11488_ _05331_ net273 _05334_ vssd1 vssd1 vccd1 vccd1 _05371_ sky130_fd_sc_hd__a21o_1
X_13227_ clknet_leaf_45_clk _00819_ net1065 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[22\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_10439_ net233 net1580 net365 vssd1 vssd1 vccd1 vccd1 _00610_ sky130_fd_sc_hd__mux2_1
XANTENNA__10145__A top.a1.instruction\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_186_Left_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08935__A1 net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09934__A _04045_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_176_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06910__X _02049_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13158_ clknet_leaf_32_clk _00750_ net1045 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[20\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_209_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06946__B1 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06410__A2 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12109_ _05986_ _05988_ _05991_ _05985_ vssd1 vssd1 vccd1 vccd1 _05992_ sky130_fd_sc_hd__a31o_2
X_13089_ clknet_leaf_16_clk _00681_ net962 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[18\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_192_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09360__A1 _02232_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07650_ _02782_ _02786_ _02787_ _02788_ vssd1 vssd1 vccd1 vccd1 _02789_ sky130_fd_sc_hd__or4_1
XFILLER_0_192_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_189_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08837__X _03950_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_195_Right_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07371__B1 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06601_ _01735_ _01737_ _01739_ vssd1 vssd1 vccd1 vccd1 _01740_ sky130_fd_sc_hd__or3_1
XFILLER_0_177_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07741__X _02880_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07910__A2 _02899_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07581_ top.DUT.register\[6\]\[6\] net567 net527 top.DUT.register\[26\]\[6\] vssd1
+ vssd1 vccd1 vccd1 _02720_ sky130_fd_sc_hd__a22o_1
X_09320_ _04381_ _04382_ vssd1 vssd1 vccd1 vccd1 _04383_ sky130_fd_sc_hd__and2b_1
X_06532_ top.DUT.register\[14\]\[29\] net586 net457 top.DUT.register\[25\]\[29\] _01670_
+ vssd1 vssd1 vccd1 vccd1 _01671_ sky130_fd_sc_hd__a221o_1
XANTENNA__07123__B1 net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09251_ _04313_ _04317_ vssd1 vssd1 vccd1 vccd1 _04318_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_75_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_177_3094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_684 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06463_ top.a1.instruction\[21\] net792 top.a1.instruction\[20\] vssd1 vssd1 vccd1
+ vccd1 _01602_ sky130_fd_sc_hd__and3b_2
XTAP_TAPCELL_ROW_32_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08202_ _02996_ _03043_ vssd1 vssd1 vccd1 vccd1 _03340_ sky130_fd_sc_hd__or2_1
XFILLER_0_7_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09754__A1_N top.a1.dataIn\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09182_ net136 _04252_ vssd1 vssd1 vccd1 vccd1 _04253_ sky130_fd_sc_hd__nor2_1
X_06394_ top.a1.instruction\[17\] top.a1.instruction\[18\] net782 vssd1 vssd1 vccd1
+ vccd1 _01533_ sky130_fd_sc_hd__and3_1
XFILLER_0_55_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_518 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08133_ _02242_ net327 vssd1 vssd1 vccd1 vccd1 _03271_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_190_3294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10754__S net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08623__B1 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09828__B _04499_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_6__f_clk clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_6__leaf_clk sky130_fd_sc_hd__clkbuf_16
XANTENNA_fanout218_A _04814_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07977__A2 net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08064_ _03199_ _03202_ net293 vssd1 vssd1 vccd1 vccd1 _03203_ sky130_fd_sc_hd__mux2_1
XFILLER_0_160_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07015_ _02149_ _02151_ _02153_ vssd1 vssd1 vccd1 vccd1 _02154_ sky130_fd_sc_hd__or3_1
XANTENNA__10981__B2 top.a1.dataIn\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09179__A1 net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12183__B1 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_4__f_clk_X clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06252__B net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06937__B1 net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout587_A net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_164_2905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08966_ net1173 net875 _02218_ _04049_ vssd1 vssd1 vccd1 vccd1 _00072_ sky130_fd_sc_hd__a22o_1
X_07917_ _02678_ _02703_ _03055_ vssd1 vssd1 vccd1 vccd1 _03056_ sky130_fd_sc_hd__o21ba_1
X_08897_ net424 _04006_ _04004_ vssd1 vssd1 vccd1 vccd1 _04007_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout754_A _01620_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_80 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout375_X net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_95_clk clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_95_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_197_3404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07848_ top.DUT.register\[18\]\[0\] net550 net511 top.DUT.register\[24\]\[0\] vssd1
+ vssd1 vccd1 vccd1 _02987_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_104_2001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_162_Right_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_104_2012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout542_X net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout921_A net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10929__S net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_195_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07779_ top.DUT.register\[23\]\[2\] net671 net742 top.DUT.register\[2\]\[2\] vssd1
+ vssd1 vccd1 vccd1 _02918_ sky130_fd_sc_hd__a22o_1
XFILLER_0_78_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_196_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09518_ _04567_ _04568_ vssd1 vssd1 vccd1 vccd1 _04569_ sky130_fd_sc_hd__or2_1
X_10790_ net1364 net150 net485 vssd1 vssd1 vccd1 vccd1 _00951_ sky130_fd_sc_hd__mux2_1
XANTENNA__08195__A net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07114__B1 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08963__A1_N net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_150 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_766 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09449_ net137 _04493_ _04504_ net901 vssd1 vssd1 vccd1 vccd1 _04505_ sky130_fd_sc_hd__o211ai_1
XANTENNA_fanout807_X net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12460_ clknet_leaf_87_clk _00055_ net1006 vssd1 vssd1 vccd1 vccd1 top.ramstore\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_10_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11411_ _01395_ _05285_ _05254_ vssd1 vssd1 vccd1 vccd1 _05294_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_62_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10664__S net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12391_ clknet_leaf_102_clk top.ru.next_FetchedInstr\[3\] net981 vssd1 vssd1 vccd1
+ vccd1 top.a1.instruction\[3\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__11213__A2 net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06714__Y _01853_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11342_ _05211_ _05219_ top.a1.dataIn\[22\] vssd1 vssd1 vccd1 vccd1 _05225_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_61_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07968__A2 net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10972__A1 top.a1.halfData\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_115_2174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06640__A2 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11273_ top.a1.row2\[2\] _05143_ _05162_ _05163_ vssd1 vssd1 vccd1 vccd1 _05164_
+ sky130_fd_sc_hd__a211o_1
XANTENNA__08917__A1 net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12174__B1 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10224_ net159 net1490 net395 vssd1 vssd1 vccd1 vccd1 _00404_ sky130_fd_sc_hd__mux2_1
X_13012_ clknet_leaf_55_clk _00604_ net1031 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[16\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06928__B1 net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10724__A1 net156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10155_ net2276 net232 net602 vssd1 vssd1 vccd1 vccd1 _00354_ sky130_fd_sc_hd__mux2_1
Xhold6 top.a1.dataInTemp\[6\] vssd1 vssd1 vccd1 vccd1 net1122 sky130_fd_sc_hd__dlygate4sd3_1
X_10086_ net2262 net243 net612 vssd1 vssd1 vccd1 vccd1 _00287_ sky130_fd_sc_hd__mux2_1
XANTENNA__08089__B _03040_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_86_clk clknet_4_6__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_86_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__09342__A1 _02580_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_540 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07353__B1 net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_202_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_202_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_159_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10839__S net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08817__B _03929_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12751__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_15__f_clk_X clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13776_ clknet_leaf_99_clk _01347_ vssd1 vssd1 vccd1 vccd1 top.lcd.cnt_500hz\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__07105__B1 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10988_ top.a1.dataInTemp\[6\] net785 vssd1 vssd1 vccd1 vccd1 _05025_ sky130_fd_sc_hd__or2_1
XFILLER_0_85_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11243__B _05128_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12727_ clknet_leaf_128_clk _00319_ net912 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[7\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13173__RESET_B net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09929__A net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12658_ clknet_leaf_23_clk _00250_ net1014 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[5\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_182_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_518 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_142_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11609_ _05461_ _05490_ _05491_ _05456_ vssd1 vssd1 vccd1 vccd1 _05492_ sky130_fd_sc_hd__a22o_1
XANTENNA__10574__S net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12589_ clknet_leaf_43_clk _00181_ net1062 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[2\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_111_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_10_clk clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_10_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_105_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_194_Left_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold406 top.DUT.register\[20\]\[28\] vssd1 vssd1 vccd1 vccd1 net1522 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_187_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xmax_cap125 _05901_ vssd1 vssd1 vccd1 vccd1 net125 sky130_fd_sc_hd__clkbuf_1
Xhold417 top.DUT.register\[17\]\[2\] vssd1 vssd1 vccd1 vccd1 net1533 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10963__A1 top.a1.dataIn\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10963__B2 net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold428 top.DUT.register\[17\]\[1\] vssd1 vssd1 vccd1 vccd1 net1544 sky130_fd_sc_hd__dlygate4sd3_1
Xhold439 top.a1.row2\[26\] vssd1 vssd1 vccd1 vccd1 net1555 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06631__A2 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06919__B1 net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout908 _01405_ vssd1 vssd1 vccd1 vccd1 net908 sky130_fd_sc_hd__clkbuf_2
Xfanout919 net921 vssd1 vssd1 vccd1 vccd1 net919 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_55_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08820_ net1489 net830 net801 _03933_ vssd1 vssd1 vccd1 vccd1 _00043_ sky130_fd_sc_hd__a22o_1
Xclkbuf_4_14__f_clk clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_14__leaf_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__07592__B1 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1106 top.DUT.register\[9\]\[17\] vssd1 vssd1 vccd1 vccd1 net2222 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_146_2635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1117 top.DUT.register\[21\]\[1\] vssd1 vssd1 vccd1 vccd1 net2233 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1128 top.DUT.register\[19\]\[19\] vssd1 vssd1 vccd1 vccd1 net2244 sky130_fd_sc_hd__dlygate4sd3_1
X_08751_ net434 _03861_ _03865_ net424 vssd1 vssd1 vccd1 vccd1 _03868_ sky130_fd_sc_hd__a2bb2o_1
Xhold1139 net124 vssd1 vssd1 vccd1 vccd1 net2255 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_77_clk clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_77_clk
+ sky130_fd_sc_hd__clkbuf_8
X_07702_ top.DUT.register\[13\]\[4\] net464 _02840_ vssd1 vssd1 vccd1 vccd1 _02841_
+ sky130_fd_sc_hd__a21o_1
X_08682_ _03263_ _03791_ _03799_ net435 vssd1 vssd1 vccd1 vccd1 _03802_ sky130_fd_sc_hd__a22oi_1
XANTENNA__07344__B1 net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_179_3134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06698__A2 net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07633_ _02767_ _02769_ _02771_ vssd1 vssd1 vccd1 vccd1 _02772_ sky130_fd_sc_hd__or3_2
XANTENNA__10749__S net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_177_234 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07190__Y _02329_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07564_ net825 _02682_ _02702_ vssd1 vssd1 vccd1 vccd1 _02703_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_0_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_192_3323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_446 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09303_ _04365_ _04366_ vssd1 vssd1 vccd1 vccd1 _04367_ sky130_fd_sc_hd__xnor2_1
X_06515_ _01649_ _01651_ _01653_ vssd1 vssd1 vccd1 vccd1 _01654_ sky130_fd_sc_hd__or3_1
X_07495_ top.DUT.register\[28\]\[14\] net767 net757 top.DUT.register\[1\]\[14\] vssd1
+ vssd1 vccd1 vccd1 _02634_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06247__B net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout335_A net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_3_Right_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06446_ top.a1.instruction\[31\] net804 _01583_ vssd1 vssd1 vccd1 vccd1 _01585_ sky130_fd_sc_hd__o21ai_4
X_09234_ _04298_ _04301_ vssd1 vssd1 vccd1 vccd1 _04302_ sky130_fd_sc_hd__xnor2_1
XANTENNA__08743__A net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_161_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10992__B net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_157_2797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09165_ top.pc\[5\] _04221_ vssd1 vssd1 vccd1 vccd1 _04237_ sky130_fd_sc_hd__nor2_1
XFILLER_0_90_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10484__S net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06870__A2 net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06377_ top.a1.instruction\[18\] net782 top.a1.instruction\[17\] vssd1 vssd1 vccd1
+ vccd1 _01516_ sky130_fd_sc_hd__and3b_2
XANTENNA__09558__B _04605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08116_ _03247_ _03254_ net311 vssd1 vssd1 vccd1 vccd1 _03255_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07359__A _02497_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09096_ _03150_ _04170_ _01389_ _01500_ vssd1 vssd1 vccd1 vccd1 _04171_ sky130_fd_sc_hd__o211a_1
XANTENNA__06263__A top.ramload\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_170_2997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08047_ _03160_ _03164_ vssd1 vssd1 vccd1 vccd1 _03186_ sky130_fd_sc_hd__nor2_1
XANTENNA__06622__A2 net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold940 top.DUT.register\[29\]\[1\] vssd1 vssd1 vccd1 vccd1 net2056 sky130_fd_sc_hd__dlygate4sd3_1
Xhold951 top.pad.button_control.r_counter\[4\] vssd1 vssd1 vccd1 vccd1 net2067 sky130_fd_sc_hd__dlygate4sd3_1
Xhold962 top.DUT.register\[16\]\[12\] vssd1 vssd1 vccd1 vccd1 net2078 sky130_fd_sc_hd__dlygate4sd3_1
Xhold973 top.DUT.register\[14\]\[10\] vssd1 vssd1 vccd1 vccd1 net2089 sky130_fd_sc_hd__dlygate4sd3_1
Xhold984 top.DUT.register\[16\]\[25\] vssd1 vssd1 vccd1 vccd1 net2100 sky130_fd_sc_hd__dlygate4sd3_1
Xhold995 top.DUT.register\[4\]\[15\] vssd1 vssd1 vccd1 vccd1 net2111 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout492_X net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07806__B _02944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09998_ net204 net1418 net624 vssd1 vssd1 vccd1 vccd1 _00203_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_110_2093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_209_3580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08949_ net2236 net877 _02796_ net693 vssd1 vssd1 vccd1 vccd1 _00055_ sky130_fd_sc_hd__a22o_1
XFILLER_0_204_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_68_clk clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_68_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__09324__A1 _02623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout757_X net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12501__Q top.pc\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11960_ _05842_ vssd1 vssd1 vccd1 vccd1 _05843_ sky130_fd_sc_hd__inv_2
XANTENNA__08477__X _03606_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10911_ net1935 net177 net480 vssd1 vssd1 vccd1 vccd1 _01072_ sky130_fd_sc_hd__mux2_1
XANTENNA__10659__S net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11891_ _05725_ _05771_ vssd1 vssd1 vccd1 vccd1 _05774_ sky130_fd_sc_hd__xnor2_1
XANTENNA__08196__Y _03334_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07541__B _02679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13630_ clknet_leaf_72_clk _01217_ net1085 vssd1 vssd1 vccd1 vccd1 net57 sky130_fd_sc_hd__dfrtp_1
X_10842_ net2279 net203 net475 vssd1 vssd1 vccd1 vccd1 _01003_ sky130_fd_sc_hd__mux2_1
XFILLER_0_196_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13561_ clknet_leaf_106_clk _01148_ net968 vssd1 vssd1 vccd1 vccd1 top.ramload\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_183_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10773_ net1942 net210 net484 vssd1 vssd1 vccd1 vccd1 _00934_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12512_ clknet_leaf_82_clk _00104_ net993 vssd1 vssd1 vccd1 vccd1 top.pc\[24\] sky130_fd_sc_hd__dfstp_2
XANTENNA__09749__A top.pc\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13492_ clknet_leaf_55_clk _01084_ net1074 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[31\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_117_2203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_23_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12443_ clknet_leaf_75_clk _00039_ net1083 vssd1 vssd1 vccd1 vccd1 top.ramaddr\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06861__A2 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12374_ clknet_leaf_107_clk top.ru.next_FetchedData\[18\] net971 vssd1 vssd1 vccd1
+ vccd1 top.a1.dataIn\[18\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_34_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_130_2403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06613__A2 net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11325_ top.a1.dataIn\[31\] top.a1.dataIn\[25\] top.a1.dataIn\[24\] top.a1.dataIn\[30\]
+ vssd1 vssd1 vccd1 vccd1 _05208_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_97_1899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11256_ net878 _05130_ _05148_ vssd1 vssd1 vccd1 vccd1 _05149_ sky130_fd_sc_hd__and3_2
XANTENNA__08366__A2 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09563__A1 net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10207_ net227 top.DUT.register\[9\]\[10\] net393 vssd1 vssd1 vccd1 vccd1 _00387_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__09563__B2 net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11187_ net1244 net588 _05098_ _05100_ vssd1 vssd1 vccd1 vccd1 _01243_ sky130_fd_sc_hd__a22o_1
XFILLER_0_206_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08855__A1_N net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10138_ net170 net1712 net607 vssd1 vssd1 vccd1 vccd1 _00338_ sky130_fd_sc_hd__mux2_1
XFILLER_0_206_124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11238__B top.lcd.nextState\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12411__Q top.a1.instruction\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_2365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10069_ net1404 net182 net616 vssd1 vssd1 vccd1 vccd1 _00271_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07326__B1 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10569__S net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_141_2554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_141_2565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13828_ net1112 vssd1 vssd1 vccd1 vccd1 gpio_out[27] sky130_fd_sc_hd__buf_2
XANTENNA__07451__B _02589_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13759_ clknet_leaf_71_clk _01330_ vssd1 vssd1 vccd1 vccd1 top.lcd.currentState\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_174_3053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06300_ _01452_ _01454_ _01456_ vssd1 vssd1 vccd1 vccd1 _01458_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_45_427 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07280_ top.DUT.register\[7\]\[13\] net660 net752 top.DUT.register\[26\]\[13\] _02418_
+ vssd1 vssd1 vccd1 vccd1 _02419_ sky130_fd_sc_hd__a221o_1
XFILLER_0_127_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06231_ top.ramload\[25\] net858 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedInstr\[25\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_122_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06852__A2 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06162_ net1 vssd1 vssd1 vccd1 vccd1 _01405_ sky130_fd_sc_hd__inv_2
XFILLER_0_81_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold203 top.DUT.register\[15\]\[17\] vssd1 vssd1 vccd1 vccd1 net1319 sky130_fd_sc_hd__dlygate4sd3_1
Xhold214 top.DUT.register\[5\]\[31\] vssd1 vssd1 vccd1 vccd1 net1330 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold225 top.DUT.register\[19\]\[17\] vssd1 vssd1 vccd1 vccd1 net1341 sky130_fd_sc_hd__dlygate4sd3_1
Xhold236 top.DUT.register\[26\]\[9\] vssd1 vssd1 vccd1 vccd1 net1352 sky130_fd_sc_hd__dlygate4sd3_1
Xhold247 top.DUT.register\[23\]\[24\] vssd1 vssd1 vccd1 vccd1 net1363 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_543 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold258 top.DUT.register\[20\]\[23\] vssd1 vssd1 vccd1 vccd1 net1374 sky130_fd_sc_hd__dlygate4sd3_1
Xhold269 top.DUT.register\[11\]\[4\] vssd1 vssd1 vccd1 vccd1 net1385 sky130_fd_sc_hd__dlygate4sd3_1
X_09921_ _04923_ _04925_ _04926_ _04927_ vssd1 vssd1 vccd1 vccd1 _04928_ sky130_fd_sc_hd__a211o_1
Xfanout705 _01642_ vssd1 vssd1 vccd1 vccd1 net705 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_1_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout716 net717 vssd1 vssd1 vccd1 vccd1 net716 sky130_fd_sc_hd__buf_4
Xfanout727 _01628_ vssd1 vssd1 vccd1 vccd1 net727 sky130_fd_sc_hd__buf_2
X_09852_ _04863_ _04864_ _04861_ vssd1 vssd1 vccd1 vccd1 _04865_ sky130_fd_sc_hd__a21oi_1
Xfanout738 _01624_ vssd1 vssd1 vccd1 vccd1 net738 sky130_fd_sc_hd__clkbuf_8
Xfanout749 _01622_ vssd1 vssd1 vccd1 vccd1 net749 sky130_fd_sc_hd__buf_4
X_08803_ _03874_ _03915_ net287 vssd1 vssd1 vccd1 vccd1 _03917_ sky130_fd_sc_hd__mux2_1
X_09783_ _04420_ net486 net402 top.a1.dataIn\[16\] net397 vssd1 vssd1 vccd1 vccd1
+ _04803_ sky130_fd_sc_hd__a221o_1
X_06995_ _02133_ vssd1 vssd1 vccd1 vccd1 _02134_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout285_A _03170_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08734_ _03811_ _03850_ _02090_ vssd1 vssd1 vccd1 vccd1 _03851_ sky130_fd_sc_hd__a21oi_2
XANTENNA__08738__A net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07317__B1 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08665_ _03334_ _03771_ _03785_ _03342_ vssd1 vssd1 vccd1 vccd1 _03786_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_1_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10479__S net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout452_A _01561_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08457__B net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07616_ top.DUT.register\[22\]\[5\] net575 net523 top.DUT.register\[11\]\[5\] vssd1
+ vssd1 vccd1 vccd1 _02755_ sky130_fd_sc_hd__a22o_1
X_08596_ net436 _03718_ _03719_ net427 vssd1 vssd1 vccd1 vccd1 _03720_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_159_2826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_159_2837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07547_ top.DUT.register\[20\]\[7\] net663 net702 top.DUT.register\[3\]\[7\] _02683_
+ vssd1 vssd1 vccd1 vccd1 _02686_ sky130_fd_sc_hd__a221o_1
XFILLER_0_119_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_193_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout338_X net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout717_A _01637_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13422__CLK clknet_leaf_40_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07096__A2 net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07478_ top.DUT.register\[30\]\[14\] net581 net513 top.DUT.register\[24\]\[14\] vssd1
+ vssd1 vccd1 vccd1 _02617_ sky130_fd_sc_hd__a22o_1
XFILLER_0_146_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09217_ _04284_ _04285_ vssd1 vssd1 vccd1 vccd1 _04286_ sky130_fd_sc_hd__or2_1
XFILLER_0_106_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_268 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06429_ top.DUT.register\[5\]\[30\] net441 net505 top.DUT.register\[27\]\[30\] vssd1
+ vssd1 vccd1 vccd1 _01568_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout505_X net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09148_ top.pc\[2\] top.pc\[3\] top.pc\[4\] vssd1 vssd1 vccd1 vccd1 _04221_ sky130_fd_sc_hd__and3_1
XFILLER_0_133_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09793__A1 net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13819__A top.lcd.lcd_en vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09079_ top.a1.instruction\[9\] top.a1.instruction\[10\] vssd1 vssd1 vccd1 vccd1
+ _04154_ sky130_fd_sc_hd__nand2_1
XANTENNA__10942__S net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_154 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_2122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08920__B _04027_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11110_ net907 net2289 net862 _05060_ vssd1 vssd1 vccd1 vccd1 _01206_ sky130_fd_sc_hd__a31o_1
XFILLER_0_188_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12090_ _05951_ _05964_ _05968_ _05966_ vssd1 vssd1 vccd1 vccd1 _05973_ sky130_fd_sc_hd__o31a_1
Xhold770 top.DUT.register\[3\]\[7\] vssd1 vssd1 vccd1 vccd1 net1886 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold781 top.DUT.register\[24\]\[14\] vssd1 vssd1 vccd1 vccd1 net1897 sky130_fd_sc_hd__dlygate4sd3_1
X_11041_ net21 net838 net816 top.ramload\[27\] vssd1 vssd1 vccd1 vccd1 _01153_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_9_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold792 top.DUT.register\[11\]\[22\] vssd1 vssd1 vccd1 vccd1 net1908 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09545__A1 net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07020__A2 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_204_628 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07308__B1 net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11104__A1 _01405_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12992_ clknet_leaf_80_clk _00584_ net992 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[15\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09848__A2 _04514_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input13_A DAT_I[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10389__S net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11943_ net128 _05818_ _05798_ _05813_ vssd1 vssd1 vccd1 vccd1 _05826_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_197_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_200_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_169_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_28_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08520__A2 net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11874_ _05747_ _05756_ vssd1 vssd1 vccd1 vccd1 _05757_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_123_2284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_123_2295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_243 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13613_ clknet_leaf_90_clk _01200_ net1002 vssd1 vssd1 vccd1 vccd1 net70 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_211_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10825_ net1670 net267 net475 vssd1 vssd1 vccd1 vccd1 _00986_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_156_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13544_ clknet_leaf_94_clk _01131_ net982 vssd1 vssd1 vccd1 vccd1 top.ramload\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07087__A2 net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10756_ net1579 net158 net420 vssd1 vssd1 vccd1 vccd1 _00917_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_1928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06295__A0 top.lcd.nextState\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_730 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09198__B top.pc\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13475_ clknet_leaf_61_clk _01067_ net1088 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[30\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_600 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10687_ net1932 net169 net339 vssd1 vssd1 vccd1 vccd1 _00850_ sky130_fd_sc_hd__mux2_1
XANTENNA__09766__X _04788_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12426_ clknet_leaf_75_clk _00022_ net1077 vssd1 vssd1 vccd1 vccd1 top.ramaddr\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_140_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_140_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12406__Q top.a1.instruction\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09784__A1 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10852__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12357_ clknet_leaf_95_clk top.ru.next_FetchedData\[1\] net982 vssd1 vssd1 vccd1
+ vccd1 top.a1.dataIn\[1\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__09926__B _04628_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11308_ top.a1.row1\[60\] _05136_ _05194_ net815 vssd1 vssd1 vccd1 vccd1 _05195_
+ sky130_fd_sc_hd__a211o_1
X_12288_ top.lcd.cnt_500hz\[11\] top.lcd.cnt_500hz\[12\] _06100_ vssd1 vssd1 vccd1
+ vccd1 _06104_ sky130_fd_sc_hd__and3_1
XFILLER_0_120_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11239_ _05129_ _05131_ vssd1 vssd1 vccd1 vccd1 _05132_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_52_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07547__B1 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_184_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07011__A2 net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_184_49 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06780_ _01897_ _01917_ vssd1 vssd1 vccd1 vccd1 _01919_ sky130_fd_sc_hd__nand2_1
XFILLER_0_89_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10299__S net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08450_ net324 _03579_ vssd1 vssd1 vccd1 vccd1 _03580_ sky130_fd_sc_hd__nand2_1
X_07401_ top.DUT.register\[3\]\[9\] net551 net439 top.DUT.register\[5\]\[9\] _02539_
+ vssd1 vssd1 vccd1 vccd1 _02540_ sky130_fd_sc_hd__a221o_1
X_08381_ _03512_ _03513_ vssd1 vssd1 vccd1 vccd1 _03514_ sky130_fd_sc_hd__or2_2
XFILLER_0_148_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_175_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10606__A0 net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_163_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07332_ _02468_ _02469_ _02470_ vssd1 vssd1 vccd1 vccd1 _02471_ sky130_fd_sc_hd__or3_1
XFILLER_0_85_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_63_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07263_ top.DUT.register\[28\]\[13\] net556 net548 top.DUT.register\[18\]\[13\] vssd1
+ vssd1 vccd1 vccd1 _02402_ sky130_fd_sc_hd__a22o_1
XFILLER_0_171_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_154_2756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09002_ _04074_ _04076_ vssd1 vssd1 vccd1 vccd1 _04077_ sky130_fd_sc_hd__nand2_1
X_06214_ net1117 net857 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedInstr\[8\] sky130_fd_sc_hd__and2_1
XFILLER_0_26_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_482 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07194_ net894 _02332_ vssd1 vssd1 vccd1 vccd1 _02333_ sky130_fd_sc_hd__nand2_1
XANTENNA__08580__X _03705_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06145_ top.a1.instruction\[3\] vssd1 vssd1 vccd1 vccd1 _01388_ sky130_fd_sc_hd__inv_2
XANTENNA__09775__A1 _03724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10762__S net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_187_3244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_187_3255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09904_ _04909_ _04910_ net798 vssd1 vssd1 vccd1 vccd1 _04912_ sky130_fd_sc_hd__o21ai_1
Xfanout502 _03186_ vssd1 vssd1 vccd1 vccd1 net502 sky130_fd_sc_hd__clkbuf_2
Xfanout513 _01559_ vssd1 vssd1 vccd1 vccd1 net513 sky130_fd_sc_hd__clkbuf_8
Xfanout524 _01554_ vssd1 vssd1 vccd1 vccd1 net524 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06260__B net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout535 _01541_ vssd1 vssd1 vccd1 vccd1 net535 sky130_fd_sc_hd__buf_6
Xfanout546 _01539_ vssd1 vssd1 vccd1 vccd1 net546 sky130_fd_sc_hd__clkbuf_8
XANTENNA__07002__A2 net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input5_A DAT_I[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09835_ _03848_ net405 net489 _04849_ vssd1 vssd1 vccd1 vccd1 _04850_ sky130_fd_sc_hd__o211a_4
Xfanout557 net558 vssd1 vssd1 vccd1 vccd1 net557 sky130_fd_sc_hd__buf_4
Xfanout568 _01525_ vssd1 vssd1 vccd1 vccd1 net568 sky130_fd_sc_hd__buf_4
XANTENNA__13276__RESET_B net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout579 _01514_ vssd1 vssd1 vccd1 vccd1 net579 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout190_X net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout667_A _01599_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08750__A2 net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09766_ _03705_ net404 net490 _04787_ vssd1 vssd1 vccd1 vccd1 _04788_ sky130_fd_sc_hd__o211a_2
X_06978_ top.DUT.register\[23\]\[23\] net672 net779 top.DUT.register\[25\]\[23\] vssd1
+ vssd1 vccd1 vccd1 _02117_ sky130_fd_sc_hd__a22o_1
X_08717_ _03342_ _03834_ vssd1 vssd1 vccd1 vccd1 _03835_ sky130_fd_sc_hd__nor2_1
XFILLER_0_179_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_179_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09697_ net827 _04208_ vssd1 vssd1 vccd1 vccd1 _04730_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_202_3469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout455_X net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09998__S net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08648_ _01962_ _03768_ vssd1 vssd1 vccd1 vccd1 _03769_ sky130_fd_sc_hd__nor2_1
XANTENNA__10002__S net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_194_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_25_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout622_X net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10937__S net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08579_ _03342_ _03685_ _03703_ net496 vssd1 vssd1 vccd1 vccd1 _03704_ sky130_fd_sc_hd__o22a_1
XFILLER_0_154_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09299__A top.pc\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10610_ net197 net2080 net347 vssd1 vssd1 vccd1 vccd1 _00775_ sky130_fd_sc_hd__mux2_1
XANTENNA__08266__A1 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_181_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11590_ _05436_ _05471_ vssd1 vssd1 vccd1 vccd1 _05473_ sky130_fd_sc_hd__nand2_1
XANTENNA__09463__B1 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_147_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10541_ net2211 net219 net354 vssd1 vssd1 vccd1 vccd1 _00708_ sky130_fd_sc_hd__mux2_1
XANTENNA__06816__A2 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11270__B1 _05161_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_279 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13260_ clknet_leaf_47_clk _00852_ net1069 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[23\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_10472_ net1736 net233 net361 vssd1 vssd1 vccd1 vccd1 _00642_ sky130_fd_sc_hd__mux2_1
XFILLER_0_161_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11022__B1 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12211_ top.lcd.cnt_20ms\[15\] top.lcd.cnt_20ms\[14\] top.lcd.cnt_20ms\[17\] top.lcd.cnt_20ms\[16\]
+ vssd1 vssd1 vccd1 vccd1 _06057_ sky130_fd_sc_hd__or4bb_1
XANTENNA__09766__A1 _03705_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10672__S net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13191_ clknet_leaf_6_clk _00783_ net937 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[21\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_103_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07777__B1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_1858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12142_ _06023_ _06024_ vssd1 vssd1 vccd1 vccd1 _06025_ sky130_fd_sc_hd__nand2_1
XANTENNA__07241__A2 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_8_Left_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12073_ _05943_ _05948_ _05955_ _05946_ vssd1 vssd1 vccd1 vccd1 _05956_ sky130_fd_sc_hd__and4bb_1
X_11024_ net3 net841 net818 net2286 vssd1 vssd1 vccd1 vccd1 _01136_ sky130_fd_sc_hd__a22o_1
XANTENNA__09762__A top.pc\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12975_ clknet_leaf_22_clk _00567_ net1033 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[14\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_188_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11926_ _05808_ vssd1 vssd1 vccd1 vccd1 _05809_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07701__B1 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09701__S net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12928__RESET_B net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_184_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11857_ _05726_ _05734_ _05738_ _05722_ vssd1 vssd1 vccd1 vccd1 _05740_ sky130_fd_sc_hd__a211o_2
XANTENNA__10847__S net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_200_675 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10808_ net225 net2219 net601 vssd1 vssd1 vccd1 vccd1 _00969_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_103_1987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_171_3012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11788_ _05641_ _05669_ vssd1 vssd1 vccd1 vccd1 _05671_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_27_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_103_1998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13527_ clknet_leaf_88_clk _01114_ net1001 vssd1 vssd1 vccd1 vccd1 top.a1.data\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06807__A2 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10739_ net1437 net222 net418 vssd1 vssd1 vccd1 vccd1 _00900_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12510__RESET_B net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07480__A2 net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13458_ clknet_leaf_25_clk _01050_ net1012 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[30\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_136_2486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12409_ clknet_leaf_109_clk top.ru.next_FetchedInstr\[21\] net975 vssd1 vssd1 vccd1
+ vccd1 top.a1.instruction\[21\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__10582__S net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13389_ clknet_leaf_43_clk _00981_ net1062 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[27\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
Xoutput105 net105 vssd1 vssd1 vccd1 vccd1 SEL_O[0] sky130_fd_sc_hd__buf_2
XFILLER_0_2_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07768__B1 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput116 net116 vssd1 vssd1 vccd1 vccd1 gpio_out[14] sky130_fd_sc_hd__buf_2
XANTENNA__07232__A2 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_195_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07950_ _01887_ _01896_ _01917_ vssd1 vssd1 vccd1 vccd1 _03089_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_208_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_195_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06901_ top.DUT.register\[26\]\[18\] net752 net724 top.DUT.register\[29\]\[18\] vssd1
+ vssd1 vccd1 vccd1 _02040_ sky130_fd_sc_hd__a22o_1
X_07881_ _03000_ _03019_ net824 vssd1 vssd1 vccd1 vccd1 _03020_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_182_3174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09620_ _04664_ vssd1 vssd1 vccd1 vccd1 _04665_ sky130_fd_sc_hd__inv_2
X_06832_ top.DUT.register\[26\]\[19\] net529 net505 top.DUT.register\[27\]\[19\] vssd1
+ vssd1 vccd1 vccd1 _01971_ sky130_fd_sc_hd__a22o_1
X_09551_ top.pc\[27\] _04577_ _04586_ vssd1 vssd1 vccd1 vccd1 _04600_ sky130_fd_sc_hd__a21o_1
X_06763_ top.DUT.register\[5\]\[24\] net654 net748 top.DUT.register\[17\]\[24\] _01898_
+ vssd1 vssd1 vccd1 vccd1 _01902_ sky130_fd_sc_hd__a221o_1
XFILLER_0_77_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08502_ _03629_ vssd1 vssd1 vccd1 vccd1 _03630_ sky130_fd_sc_hd__inv_2
XFILLER_0_144_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06694_ _01831_ _01832_ vssd1 vssd1 vccd1 vccd1 _01833_ sky130_fd_sc_hd__nand2b_2
XANTENNA__07299__A2 net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09482_ top.pc\[24\] _04521_ vssd1 vssd1 vccd1 vccd1 _04535_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_65_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_144_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08433_ _03263_ _03561_ _03563_ _03557_ vssd1 vssd1 vccd1 vccd1 _03564_ sky130_fd_sc_hd__a211o_1
XANTENNA__10757__S net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_192 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_319 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout150_A _04938_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout248_A _04749_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08364_ net315 _03496_ vssd1 vssd1 vccd1 vccd1 _03497_ sky130_fd_sc_hd__nor2_1
XFILLER_0_46_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_160_51 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07315_ top.DUT.register\[15\]\[12\] net706 net698 top.DUT.register\[31\]\[12\] vssd1
+ vssd1 vccd1 vccd1 _02454_ sky130_fd_sc_hd__a22o_1
XFILLER_0_61_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08295_ net885 top.pc\[3\] net696 _03430_ vssd1 vssd1 vccd1 vccd1 _03431_ sky130_fd_sc_hd__a22o_1
XANTENNA__06255__B net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07246_ _02365_ _02384_ net825 vssd1 vssd1 vccd1 vccd1 _02385_ sky130_fd_sc_hd__mux2_2
XFILLER_0_116_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07471__A2 _02609_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_171_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10492__S net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07177_ top.DUT.register\[18\]\[10\] net547 net447 top.DUT.register\[21\]\[10\] _02315_
+ vssd1 vssd1 vccd1 vccd1 _02316_ sky130_fd_sc_hd__a221o_1
XANTENNA__09566__B _04605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13457__RESET_B net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout310 net314 vssd1 vssd1 vccd1 vccd1 net310 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_167_2947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_167_2958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout321 net323 vssd1 vssd1 vccd1 vccd1 net321 sky130_fd_sc_hd__buf_2
Xfanout332 _02975_ vssd1 vssd1 vccd1 vccd1 net332 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09582__A _01572_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout343 _04992_ vssd1 vssd1 vccd1 vccd1 net343 sky130_fd_sc_hd__buf_4
Xfanout354 _04989_ vssd1 vssd1 vccd1 vccd1 net354 sky130_fd_sc_hd__buf_6
XANTENNA_fanout572_X net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout951_A net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_204_3509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout365 net368 vssd1 vssd1 vccd1 vccd1 net365 sky130_fd_sc_hd__buf_6
Xfanout376 _04981_ vssd1 vssd1 vccd1 vccd1 net376 sky130_fd_sc_hd__buf_4
XANTENNA__08723__A2 net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout387 net388 vssd1 vssd1 vccd1 vccd1 net387 sky130_fd_sc_hd__clkbuf_8
XANTENNA__11617__A top.a1.dataIn\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09818_ top.pc\[20\] _04487_ vssd1 vssd1 vccd1 vccd1 _04834_ sky130_fd_sc_hd__and2_1
Xfanout398 _04753_ vssd1 vssd1 vccd1 vccd1 net398 sky130_fd_sc_hd__dlymetal6s2s_1
X_09749_ top.pc\[13\] _04370_ vssd1 vssd1 vccd1 vccd1 _04772_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_107_2054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout837_X net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12760_ clknet_leaf_127_clk _00352_ net918 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[8\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_96_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11086__A3 net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11711_ top.a1.dataIn\[10\] _05525_ _05550_ vssd1 vssd1 vccd1 vccd1 _05594_ sky130_fd_sc_hd__or3_1
XFILLER_0_84_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_2243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12691_ clknet_leaf_124_clk _00283_ net926 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[6\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10667__S net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11642_ _05523_ _05524_ vssd1 vssd1 vccd1 vccd1 _05525_ sky130_fd_sc_hd__or2_1
XFILLER_0_49_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_154_516 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_324 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11573_ _05454_ _05455_ vssd1 vssd1 vccd1 vccd1 _05456_ sky130_fd_sc_hd__or2_1
XFILLER_0_107_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold996_A top.ramload\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput18 DAT_I[24] vssd1 vssd1 vccd1 vccd1 net18 sky130_fd_sc_hd__buf_1
XANTENNA__07998__B1 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13312_ clknet_leaf_17_clk _00904_ net1032 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[25\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_10524_ net1388 net156 net359 vssd1 vssd1 vccd1 vccd1 _00693_ sky130_fd_sc_hd__mux2_1
XFILLER_0_162_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_238 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput29 DAT_I[5] vssd1 vssd1 vccd1 vccd1 net29 sky130_fd_sc_hd__buf_1
XFILLER_0_122_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13243_ clknet_leaf_125_clk _00835_ net924 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[23\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09739__B2 top.a1.dataIn\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10455_ net170 net2100 net365 vssd1 vssd1 vccd1 vccd1 _00626_ sky130_fd_sc_hd__mux2_1
XANTENNA__09476__B _02111_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13174_ clknet_leaf_4_clk _00766_ net939 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[21\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_10386_ top.DUT.register\[14\]\[24\] net174 net376 vssd1 vssd1 vccd1 vccd1 _00561_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12125_ top.a1.dataIn\[2\] _06000_ _06004_ vssd1 vssd1 vccd1 vccd1 _06008_ sky130_fd_sc_hd__or3_1
XPHY_EDGE_ROW_176_Right_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09492__A _01887_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12056_ _05909_ _05937_ _05918_ vssd1 vssd1 vccd1 vccd1 _05939_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_74_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11007_ top.a1.dataInTemp\[11\] net785 vssd1 vssd1 vccd1 vccd1 _05039_ sky130_fd_sc_hd__or2_1
XANTENNA__11246__B _05118_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_204_266 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12958_ clknet_leaf_54_clk _00550_ net1031 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[14\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_181_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_158_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11909_ _05758_ _05779_ _05782_ _05787_ _05781_ vssd1 vssd1 vccd1 vccd1 _05792_ sky130_fd_sc_hd__a41o_1
XTAP_TAPCELL_ROW_47_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_47_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10577__S net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12889_ clknet_leaf_11_clk _00481_ net951 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[12\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_135_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_2515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07100_ top.DUT.register\[23\]\[16\] net572 net524 top.DUT.register\[11\]\[16\] vssd1
+ vssd1 vccd1 vccd1 _02239_ sky130_fd_sc_hd__a22o_1
XANTENNA__07989__B1 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08080_ _01940_ net328 vssd1 vssd1 vccd1 vccd1 _03219_ sky130_fd_sc_hd__nand2_1
XFILLER_0_82_182 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_151_2704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07453__A2 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_262 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_151_2715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07031_ top.DUT.register\[20\]\[20\] net666 net735 top.DUT.register\[16\]\[20\] vssd1
+ vssd1 vccd1 vccd1 _02170_ sky130_fd_sc_hd__a22o_1
XANTENNA__06661__B1 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06362__Y _01501_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_388 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_184_3203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08982_ _03722_ _03728_ _03748_ _04056_ vssd1 vssd1 vccd1 vccd1 _04057_ sky130_fd_sc_hd__and4_1
XFILLER_0_139_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_143_Right_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07933_ _02656_ _03069_ _03071_ vssd1 vssd1 vccd1 vccd1 _03072_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_149_2677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_149_2688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout198_A _04788_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07864_ top.DUT.register\[2\]\[1\] net744 net732 top.DUT.register\[14\]\[1\] vssd1
+ vssd1 vccd1 vccd1 _03003_ sky130_fd_sc_hd__a22o_1
X_09603_ top.pc\[31\] _04628_ vssd1 vssd1 vccd1 vccd1 _04649_ sky130_fd_sc_hd__xor2_1
X_06815_ top.DUT.register\[20\]\[17\] net664 _01952_ _01953_ vssd1 vssd1 vccd1 vccd1
+ _01954_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_162_2877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07795_ _02927_ _02929_ _02931_ _02933_ vssd1 vssd1 vccd1 vccd1 _02934_ sky130_fd_sc_hd__or4_4
XANTENNA_fanout365_A net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09534_ top.pc\[27\] _04577_ vssd1 vssd1 vccd1 vccd1 _04584_ sky130_fd_sc_hd__xor2_1
X_06746_ top.DUT.register\[28\]\[24\] net557 net548 top.DUT.register\[18\]\[24\] vssd1
+ vssd1 vccd1 vccd1 _01885_ sky130_fd_sc_hd__a22o_1
XANTENNA__08469__B2 net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_455 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10487__S net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09465_ net137 _04508_ _04519_ vssd1 vssd1 vccd1 vccd1 _04520_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_195_3365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06677_ top.DUT.register\[9\]\[26\] net764 net716 top.DUT.register\[27\]\[26\] vssd1
+ vssd1 vccd1 vccd1 _01816_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout532_A _01542_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_195_3376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08416_ net423 _03520_ _03547_ vssd1 vssd1 vccd1 vccd1 _03548_ sky130_fd_sc_hd__a21bo_2
XFILLER_0_171_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07692__A2 net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06266__A top.ramload\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09396_ _02016_ _02025_ _04453_ vssd1 vssd1 vccd1 vccd1 _04455_ sky130_fd_sc_hd__or3_1
XFILLER_0_163_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_148_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_163_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_352 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout320_X net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08347_ net302 _03327_ _03371_ vssd1 vssd1 vccd1 vccd1 _03481_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout418_X net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_89_Left_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07444__A2 net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08278_ _03048_ _03413_ vssd1 vssd1 vccd1 vccd1 _03414_ sky130_fd_sc_hd__xor2_1
XANTENNA__06652__B1 net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout999_A net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07229_ top.DUT.register\[5\]\[10\] net651 net639 top.DUT.register\[8\]\[10\] vssd1
+ vssd1 vccd1 vccd1 _02368_ sky130_fd_sc_hd__a22o_1
XANTENNA__09296__B top.pc\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09864__X _04876_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10240_ net229 net2230 net389 vssd1 vssd1 vccd1 vccd1 _00419_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_91_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06404__B1 net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10171_ net2115 net170 net603 vssd1 vssd1 vccd1 vccd1 _00370_ sky130_fd_sc_hd__mux2_1
XANTENNA__10950__S net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_110_Right_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout140 net141 vssd1 vssd1 vccd1 vccd1 net140 sky130_fd_sc_hd__clkbuf_2
Xfanout151 _04938_ vssd1 vssd1 vccd1 vccd1 net151 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout162 _04906_ vssd1 vssd1 vccd1 vccd1 net162 sky130_fd_sc_hd__buf_1
Xfanout173 _04876_ vssd1 vssd1 vccd1 vccd1 net173 sky130_fd_sc_hd__buf_1
Xfanout184 net187 vssd1 vssd1 vccd1 vccd1 net184 sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_98_Left_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout195 _04850_ vssd1 vssd1 vccd1 vccd1 net195 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_202_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_89_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_202_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_198_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12812_ clknet_leaf_62_clk _00404_ net1089 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[9\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_199_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_198_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13792_ clknet_leaf_68_clk _01361_ vssd1 vssd1 vccd1 vccd1 top.pad.button_control.r_counter\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__09121__A2 _02934_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_70_clk_A clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12743_ clknet_leaf_6_clk _00335_ net944 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[7\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07683__A2 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06176__A top.a1.halfData\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12674_ clknet_leaf_25_clk _00266_ net1012 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[5\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08943__X _04050_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_181_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_166_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06891__B1 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11625_ _05459_ _05490_ vssd1 vssd1 vccd1 vccd1 _05508_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_100_1946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_683 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_85_clk_A clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_42_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11556_ _05432_ _05437_ _05438_ vssd1 vssd1 vccd1 vccd1 _05439_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_52_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07435__A2 net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13379__RESET_B net1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10507_ net1880 net221 net357 vssd1 vssd1 vccd1 vccd1 _00676_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_133_2434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_133_2445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11487_ _05331_ _05334_ net273 vssd1 vssd1 vccd1 vccd1 _05370_ sky130_fd_sc_hd__nand3_1
X_13226_ clknet_leaf_118_clk _00818_ net957 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[22\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_10438_ net238 net1677 net368 vssd1 vssd1 vccd1 vccd1 _00609_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12192__A1 top.a1.dataIn\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13157_ clknet_leaf_35_clk _00749_ net1041 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[20\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09934__B net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10860__S net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10369_ net1640 net247 net373 vssd1 vssd1 vccd1 vccd1 _00544_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12108_ _05990_ _05965_ _05989_ vssd1 vssd1 vccd1 vccd1 _05991_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13088_ clknet_leaf_55_clk _00680_ net1072 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[18\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_23_clk_A clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12039_ _05892_ _05921_ _05901_ vssd1 vssd1 vccd1 vccd1 _05922_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09896__B1 _04904_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_192_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06600_ top.DUT.register\[24\]\[28\] net646 net764 top.DUT.register\[9\]\[28\] _01738_
+ vssd1 vssd1 vccd1 vccd1 _01739_ sky130_fd_sc_hd__a221o_1
X_07580_ top.DUT.register\[22\]\[6\] net575 net447 top.DUT.register\[21\]\[6\] _02718_
+ vssd1 vssd1 vccd1 vccd1 _02719_ sky130_fd_sc_hd__a221o_1
XFILLER_0_149_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08566__A net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_38_clk_A clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06531_ top.DUT.register\[30\]\[29\] net582 net533 top.DUT.register\[12\]\[29\] vssd1
+ vssd1 vccd1 vccd1 _01670_ sky130_fd_sc_hd__a22o_1
XFILLER_0_177_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_628 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07123__A1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12088__A top.a1.dataIn\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08285__B net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08320__B1 _03454_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10100__S net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09250_ _04315_ _04316_ vssd1 vssd1 vccd1 vccd1 _04317_ sky130_fd_sc_hd__nor2_1
X_06462_ _01600_ vssd1 vssd1 vccd1 vccd1 _01601_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_177_3095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07674__A2 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08201_ _03159_ _03182_ vssd1 vssd1 vccd1 vccd1 _03339_ sky130_fd_sc_hd__or2_1
XANTENNA__06882__B1 net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06393_ _01511_ _01512_ _01531_ vssd1 vssd1 vccd1 vccd1 _01532_ sky130_fd_sc_hd__and3_4
X_09181_ top.pc\[6\] _04236_ vssd1 vssd1 vccd1 vccd1 _04252_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_28_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08132_ _02590_ net299 vssd1 vssd1 vccd1 vccd1 _03270_ sky130_fd_sc_hd__nand2_1
XANTENNA__08623__A1 net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_190_3295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08063_ _03200_ _03201_ vssd1 vssd1 vccd1 vccd1 _03202_ sky130_fd_sc_hd__nand2_1
XFILLER_0_113_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07014_ top.DUT.register\[2\]\[20\] net562 net457 top.DUT.register\[25\]\[20\] _02152_
+ vssd1 vssd1 vccd1 vccd1 _02153_ sky130_fd_sc_hd__a221o_1
XFILLER_0_101_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12183__A1 top.a1.row2\[34\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10770__S net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1022_A net1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08965_ net413 net691 net1152 net875 vssd1 vssd1 vccd1 vccd1 _00071_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_164_2906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout482_A _04962_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11167__A net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07916_ _02754_ _03054_ _02750_ vssd1 vssd1 vccd1 vccd1 _03055_ sky130_fd_sc_hd__o21a_1
X_08896_ _03098_ _04005_ vssd1 vssd1 vccd1 vccd1 _04006_ sky130_fd_sc_hd__nor2_1
XANTENNA__12684__RESET_B net1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07847_ top.DUT.register\[10\]\[0\] net519 _02985_ vssd1 vssd1 vccd1 vccd1 _02986_
+ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_197_3405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout747_A _01622_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout368_X net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_2002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_2013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07778_ top.DUT.register\[4\]\[2\] net667 net766 top.DUT.register\[28\]\[2\] _02916_
+ vssd1 vssd1 vccd1 vccd1 _02917_ sky130_fd_sc_hd__a221o_1
X_09517_ top.pc\[26\] _04556_ vssd1 vssd1 vccd1 vccd1 _04568_ sky130_fd_sc_hd__nor2_1
X_06729_ top.DUT.register\[5\]\[25\] net651 net723 top.DUT.register\[29\]\[25\] _01867_
+ vssd1 vssd1 vccd1 vccd1 _01868_ sky130_fd_sc_hd__a221o_1
XFILLER_0_93_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout535_X net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_195_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09448_ net133 _04496_ _04497_ _04503_ net811 vssd1 vssd1 vccd1 vccd1 _04504_ sky130_fd_sc_hd__o32a_1
XANTENNA__10010__S net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_162 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_778 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_163_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06873__B1 net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout702_X net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09379_ _01930_ _01939_ _04438_ vssd1 vssd1 vccd1 vccd1 _04439_ sky130_fd_sc_hd__o21a_1
XFILLER_0_47_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11410_ _01395_ _05285_ vssd1 vssd1 vccd1 vccd1 _05293_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_164_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12390_ clknet_leaf_103_clk top.ru.next_FetchedInstr\[2\] net976 vssd1 vssd1 vccd1
+ vccd1 top.a1.instruction\[2\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__07417__A2 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13472__RESET_B net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11341_ top.a1.dataIn\[19\] _05220_ _05221_ _05222_ vssd1 vssd1 vccd1 vccd1 _05224_
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_104_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08090__A2 _03177_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13401__RESET_B net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_2164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_115_2175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11272_ top.a1.row1\[2\] _05124_ _05125_ top.a1.row1\[18\] vssd1 vssd1 vccd1 vccd1
+ _05163_ sky130_fd_sc_hd__a22o_1
XANTENNA__08378__B1 net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13011_ clknet_leaf_124_clk _00603_ net926 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[16\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_10223_ net167 net1665 net395 vssd1 vssd1 vccd1 vccd1 _00403_ sky130_fd_sc_hd__mux2_1
XANTENNA__10680__S net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09105__A_N _04172_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07050__B1 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10154_ net1468 net235 net603 vssd1 vssd1 vccd1 vccd1 _00353_ sky130_fd_sc_hd__mux2_1
XANTENNA__08003__X _03142_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold7 top.pad.button_control.r_counter\[16\] vssd1 vssd1 vccd1 vccd1 net1123 sky130_fd_sc_hd__dlygate4sd3_1
X_10085_ net2038 net253 net611 vssd1 vssd1 vccd1 vccd1 _00286_ sky130_fd_sc_hd__mux2_1
XANTENNA__09342__A2 _02589_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_18_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_199_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06458__X _01597_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08386__A _02678_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13775_ clknet_leaf_99_clk _01346_ vssd1 vssd1 vccd1 vccd1 top.lcd.cnt_500hz\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_202_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10987_ top.a1.data\[2\] net783 vssd1 vssd1 vccd1 vccd1 _05024_ sky130_fd_sc_hd__or2_1
XFILLER_0_186_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06465__C_N top.a1.instruction\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12726_ clknet_leaf_12_clk _00318_ net942 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[7\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06459__A3 top.a1.instruction\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07656__A2 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12657_ clknet_leaf_112_clk _00249_ net988 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[5\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10855__S net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_603 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11540__A top.a1.dataIn\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_631 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_491 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11608_ _05457_ _05458_ net234 _05476_ _05453_ vssd1 vssd1 vccd1 vccd1 _05491_ sky130_fd_sc_hd__a221o_1
XFILLER_0_155_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_143_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12588_ clknet_leaf_64_clk _00180_ net1092 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[2\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_170_647 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06616__B1 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11539_ _05396_ _05398_ _05365_ vssd1 vssd1 vccd1 vccd1 _05422_ sky130_fd_sc_hd__a21oi_1
Xhold407 top.DUT.register\[20\]\[21\] vssd1 vssd1 vccd1 vccd1 net1523 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold418 top.DUT.register\[31\]\[17\] vssd1 vssd1 vccd1 vccd1 net1534 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_187_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold429 top.DUT.register\[21\]\[23\] vssd1 vssd1 vccd1 vccd1 net1545 sky130_fd_sc_hd__dlygate4sd3_1
X_13209_ clknet_leaf_15_clk _00801_ net959 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[22\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10590__S net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout909 net910 vssd1 vssd1 vccd1 vccd1 net909 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_55_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07041__B1 net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08750_ _02220_ net499 net426 _03854_ _03866_ vssd1 vssd1 vccd1 vccd1 _03867_ sky130_fd_sc_hd__a221o_1
Xhold1107 top.DUT.register\[6\]\[7\] vssd1 vssd1 vccd1 vccd1 net2223 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_146_2636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1118 top.DUT.register\[30\]\[28\] vssd1 vssd1 vccd1 vccd1 net2234 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1129 top.DUT.register\[7\]\[3\] vssd1 vssd1 vccd1 vccd1 net2245 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09680__A net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07701_ top.DUT.register\[15\]\[4\] net681 net677 top.DUT.register\[31\]\[4\] vssd1
+ vssd1 vccd1 vccd1 _02840_ sky130_fd_sc_hd__a22o_1
X_08681_ _02007_ net493 _03792_ _03258_ vssd1 vssd1 vccd1 vccd1 _03801_ sky130_fd_sc_hd__o22a_1
XFILLER_0_45_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_179_3124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07632_ top.DUT.register\[18\]\[5\] net547 net455 top.DUT.register\[25\]\[5\] _02770_
+ vssd1 vssd1 vccd1 vccd1 _02771_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_179_3135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07895__A2 net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_246 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07563_ net809 _02701_ vssd1 vssd1 vccd1 vccd1 _02702_ sky130_fd_sc_hd__or2_1
XFILLER_0_165_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09302_ _04346_ _04347_ _04348_ vssd1 vssd1 vccd1 vccd1 _04366_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_0_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06514_ top.DUT.register\[21\]\[30\] net657 net767 top.DUT.register\[28\]\[30\] _01652_
+ vssd1 vssd1 vccd1 vccd1 _01653_ sky130_fd_sc_hd__a221o_1
XFILLER_0_152_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_192_3324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_458 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08844__A1 _01764_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07647__A2 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07494_ _02623_ _02632_ vssd1 vssd1 vccd1 vccd1 _02633_ sky130_fd_sc_hd__nor2_2
XFILLER_0_186_791 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06855__B1 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09233_ _04299_ _04300_ vssd1 vssd1 vccd1 vccd1 _04301_ sky130_fd_sc_hd__nor2_1
XFILLER_0_61_83 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06445_ top.a1.instruction\[31\] net804 _01583_ vssd1 vssd1 vccd1 vccd1 _01584_ sky130_fd_sc_hd__o21a_2
XANTENNA__10765__S net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout230_A _04763_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_132 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11450__A top.a1.dataIn\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_157_2798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09164_ top.pc\[5\] _04221_ vssd1 vssd1 vccd1 vccd1 _04236_ sky130_fd_sc_hd__and2_1
XFILLER_0_146_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06376_ top.DUT.register\[14\]\[30\] net585 net581 top.DUT.register\[30\]\[30\] vssd1
+ vssd1 vccd1 vccd1 _01515_ sky130_fd_sc_hd__a22o_1
XFILLER_0_44_664 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08115_ _03250_ _03253_ net292 vssd1 vssd1 vccd1 vccd1 _03254_ sky130_fd_sc_hd__mux2_1
XANTENNA__06607__B1 net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_303 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_211_3630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09095_ net894 _01392_ _02345_ vssd1 vssd1 vccd1 vccd1 _04170_ sky130_fd_sc_hd__o21ai_1
XANTENNA__06263__B net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07280__B1 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08046_ _03181_ _03182_ vssd1 vssd1 vccd1 vccd1 _03185_ sky130_fd_sc_hd__or2_4
XTAP_TAPCELL_ROW_170_2998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold930 top.DUT.register\[26\]\[11\] vssd1 vssd1 vccd1 vccd1 net2046 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold941 top.lcd.cnt_20ms\[11\] vssd1 vssd1 vccd1 vccd1 net2057 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_141_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold952 top.DUT.register\[15\]\[10\] vssd1 vssd1 vccd1 vccd1 net2068 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold963 top.DUT.register\[9\]\[6\] vssd1 vssd1 vccd1 vccd1 net2079 sky130_fd_sc_hd__dlygate4sd3_1
Xhold974 top.pad.keyCode\[4\] vssd1 vssd1 vccd1 vccd1 net2090 sky130_fd_sc_hd__dlygate4sd3_1
Xhold985 top.DUT.register\[22\]\[14\] vssd1 vssd1 vccd1 vccd1 net2101 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1025_X net1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold996 top.ramload\[29\] vssd1 vssd1 vccd1 vccd1 net2112 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12865__RESET_B net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07032__B1 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09997_ net215 net1634 net626 vssd1 vssd1 vccd1 vccd1 _00202_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout485_X net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout864_A net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_2094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_209_3581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08948_ _02827_ net691 net1222 net874 vssd1 vssd1 vccd1 vccd1 _00054_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__09324__A2 _02632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout652_X net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08879_ _03988_ _03989_ vssd1 vssd1 vccd1 vccd1 _03990_ sky130_fd_sc_hd__or2_1
XANTENNA__07335__A1 _02443_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10910_ net1354 net183 net479 vssd1 vssd1 vccd1 vccd1 _01071_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_86_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11890_ _05726_ _05771_ _05772_ _05723_ vssd1 vssd1 vccd1 vccd1 _05773_ sky130_fd_sc_hd__a22oi_2
XANTENNA__07886__A2 net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10841_ net1386 net215 net477 vssd1 vssd1 vccd1 vccd1 _01002_ sky130_fd_sc_hd__mux2_1
XANTENNA__07099__B1 net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13560_ clknet_leaf_105_clk _01147_ net968 vssd1 vssd1 vccd1 vccd1 top.ramload\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_17_Left_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10772_ net1869 net211 net482 vssd1 vssd1 vccd1 vccd1 _00933_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12511_ clknet_leaf_78_clk _00103_ net1074 vssd1 vssd1 vccd1 vccd1 top.pc\[23\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__06846__B1 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13491_ clknet_leaf_121_clk _01083_ net934 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[31\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09749__B _04370_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10675__S net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_117_2204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12442_ clknet_leaf_72_clk _00038_ net1080 vssd1 vssd1 vccd1 vccd1 top.ramaddr\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_23_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12373_ clknet_leaf_105_clk top.ru.next_FetchedData\[17\] net971 vssd1 vssd1 vccd1
+ vccd1 top.a1.dataIn\[17\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_50_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_563 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06173__B top.a1.halfData\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11324_ top.a1.dataIn\[25\] top.a1.dataIn\[24\] vssd1 vssd1 vccd1 vccd1 _05207_ sky130_fd_sc_hd__and2_1
XANTENNA__07271__B1 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_26_Left_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11255_ top.lcd.nextState\[3\] _05128_ vssd1 vssd1 vccd1 vccd1 _05148_ sky130_fd_sc_hd__and2b_2
XANTENNA__06460__Y _01599_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07023__B1 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10206_ net233 net1443 net393 vssd1 vssd1 vccd1 vccd1 _00386_ sky130_fd_sc_hd__mux2_1
X_11186_ top.a1.data\[8\] net783 _05031_ vssd1 vssd1 vccd1 vccd1 _05100_ sky130_fd_sc_hd__o21a_1
XFILLER_0_207_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12599__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_207_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10137_ net172 net1808 net609 vssd1 vssd1 vccd1 vccd1 _00337_ sky130_fd_sc_hd__mux2_1
XFILLER_0_206_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_174_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_128_2366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10068_ net1692 net195 net618 vssd1 vssd1 vccd1 vccd1 _00270_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_13_Right_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_203_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07877__A2 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_141_2555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_141_2566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_35_Left_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13827_ net1111 vssd1 vssd1 vccd1 vccd1 gpio_out[26] sky130_fd_sc_hd__buf_2
XANTENNA__07629__A2 net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13758_ clknet_leaf_71_clk _01329_ vssd1 vssd1 vccd1 vccd1 top.lcd.currentState\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__06837__B1 net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_174_3054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12709_ clknet_leaf_34_clk _00301_ net1040 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[6\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_155_430 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10585__S net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13689_ clknet_leaf_71_clk _00001_ vssd1 vssd1 vccd1 vccd1 top.lcd.nextState\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_155_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06230_ top.ramload\[24\] net858 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedInstr\[24\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_72_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_22_Right_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_198_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11189__A2 net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06161_ top.lcd.cnt_500hz\[14\] vssd1 vssd1 vccd1 vccd1 _01404_ sky130_fd_sc_hd__inv_2
XFILLER_0_170_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold204 top.DUT.register\[15\]\[28\] vssd1 vssd1 vccd1 vccd1 net1320 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09675__A top.a1.instruction\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold215 top.DUT.register\[31\]\[22\] vssd1 vssd1 vccd1 vccd1 net1331 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07801__A2 net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_44_Left_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold226 top.DUT.register\[8\]\[5\] vssd1 vssd1 vccd1 vccd1 net1342 sky130_fd_sc_hd__dlygate4sd3_1
Xhold237 top.DUT.register\[15\]\[23\] vssd1 vssd1 vccd1 vccd1 net1353 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold248 top.DUT.register\[26\]\[30\] vssd1 vssd1 vccd1 vccd1 net1364 sky130_fd_sc_hd__dlygate4sd3_1
X_09920_ top.a1.instruction\[29\] net487 net402 top.a1.dataIn\[29\] net398 vssd1 vssd1
+ vccd1 vccd1 _04927_ sky130_fd_sc_hd__a221o_2
XANTENNA__11269__X _05161_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold259 top.DUT.register\[11\]\[19\] vssd1 vssd1 vccd1 vccd1 net1375 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07014__B1 net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout706 _01640_ vssd1 vssd1 vccd1 vccd1 net706 sky130_fd_sc_hd__buf_4
XFILLER_0_1_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09851_ top.pc\[23\] _01584_ vssd1 vssd1 vccd1 vccd1 _04864_ sky130_fd_sc_hd__or2_1
Xfanout717 _01637_ vssd1 vssd1 vccd1 vccd1 net717 sky130_fd_sc_hd__buf_4
XANTENNA__08962__A1_N _02045_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout728 _01628_ vssd1 vssd1 vccd1 vccd1 net728 sky130_fd_sc_hd__clkbuf_8
Xfanout739 _01624_ vssd1 vssd1 vccd1 vccd1 net739 sky130_fd_sc_hd__buf_4
X_08802_ _03915_ vssd1 vssd1 vccd1 vccd1 _03916_ sky130_fd_sc_hd__inv_2
X_09782_ _04149_ _04751_ vssd1 vssd1 vccd1 vccd1 _04802_ sky130_fd_sc_hd__nor2_1
X_06994_ _02112_ _02132_ vssd1 vssd1 vccd1 vccd1 _02133_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_31_Right_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08733_ _02091_ _02177_ vssd1 vssd1 vccd1 vccd1 _03850_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout180_A _04858_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08664_ _02049_ _03783_ vssd1 vssd1 vccd1 vccd1 _03785_ sky130_fd_sc_hd__xor2_1
XPHY_EDGE_ROW_53_Left_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07868__A2 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07615_ _02751_ _02752_ vssd1 vssd1 vccd1 vccd1 _02754_ sky130_fd_sc_hd__nor2_2
X_08595_ _03535_ _03709_ vssd1 vssd1 vccd1 vccd1 _03719_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout445_A net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06258__B net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_159_2827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_159_2838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07546_ top.DUT.register\[16\]\[7\] net734 net710 top.DUT.register\[11\]\[7\] _02684_
+ vssd1 vssd1 vccd1 vccd1 _02685_ sky130_fd_sc_hd__a221o_1
XFILLER_0_76_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_715 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06828__B1 net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_81_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_181_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout612_A _04955_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09490__A1 top.a1.instruction\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07477_ top.DUT.register\[22\]\[14\] net576 net458 top.DUT.register\[25\]\[14\] _02615_
+ vssd1 vssd1 vccd1 vccd1 _02616_ sky130_fd_sc_hd__a221o_1
XFILLER_0_119_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_40_Right_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09216_ top.pc\[8\] _04268_ vssd1 vssd1 vccd1 vccd1 _04285_ sky130_fd_sc_hd__nor2_1
X_06428_ net684 _01518_ _01521_ vssd1 vssd1 vccd1 vccd1 _01567_ sky130_fd_sc_hd__and3_4
XFILLER_0_106_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_496 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09147_ net900 top.pc\[3\] _04209_ _04220_ net890 vssd1 vssd1 vccd1 vccd1 _00083_
+ sky130_fd_sc_hd__o221a_1
X_06359_ net1259 net1119 _01498_ vssd1 vssd1 vccd1 vccd1 _00017_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout400_X net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_62_Left_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07657__X _02796_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07253__B1 net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09078_ top.a1.instruction\[9\] top.a1.instruction\[10\] vssd1 vssd1 vccd1 vccd1
+ _04153_ sky130_fd_sc_hd__and2_2
XANTENNA_fanout981_A net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_2123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08029_ _03160_ _03167_ vssd1 vssd1 vccd1 vccd1 _03168_ sky130_fd_sc_hd__nor2_2
Xhold760 top.DUT.register\[10\]\[8\] vssd1 vssd1 vccd1 vccd1 net1876 sky130_fd_sc_hd__dlygate4sd3_1
Xhold771 top.DUT.register\[25\]\[19\] vssd1 vssd1 vccd1 vccd1 net1887 sky130_fd_sc_hd__dlygate4sd3_1
Xhold782 top.DUT.register\[1\]\[19\] vssd1 vssd1 vccd1 vccd1 net1898 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07005__B1 net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11040_ net20 net841 net818 net2308 vssd1 vssd1 vccd1 vccd1 _01152_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_9_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold793 top.DUT.register\[21\]\[25\] vssd1 vssd1 vccd1 vccd1 net1909 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout867_X net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12512__Q top.pc\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08488__X _03617_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06182__A1_N net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_204_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_71_Left_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12991_ clknet_leaf_19_clk _00583_ net1027 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[15\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_207_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_203_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11942_ _05814_ _05823_ _05824_ vssd1 vssd1 vccd1 vccd1 _05825_ sky130_fd_sc_hd__o21a_1
XFILLER_0_200_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_28_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11873_ _05740_ _05752_ vssd1 vssd1 vccd1 vccd1 _05756_ sky130_fd_sc_hd__and2_1
XANTENNA__06531__A2 net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_2285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_514 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13612_ clknet_leaf_89_clk _01199_ net1003 vssd1 vssd1 vccd1 vccd1 net69 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_123_2296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10824_ net1529 net145 net474 vssd1 vssd1 vccd1 vccd1 _00985_ sky130_fd_sc_hd__mux2_1
XANTENNA__08664__A _02049_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_255 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13543_ clknet_leaf_95_clk _01130_ net981 vssd1 vssd1 vccd1 vccd1 top.ramload\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10755_ net1399 net160 net420 vssd1 vssd1 vccd1 vccd1 _00916_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_603 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_99_1929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13474_ clknet_leaf_9_clk _01066_ net947 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[30\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07492__B1 net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10686_ net1363 net174 net340 vssd1 vssd1 vccd1 vccd1 _00849_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_80_Left_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_180_742 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12425_ clknet_leaf_87_clk _00021_ net1004 vssd1 vssd1 vccd1 vccd1 top.ramaddr\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06471__X _01610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12356_ clknet_leaf_102_clk top.ru.next_FetchedData\[0\] net981 vssd1 vssd1 vccd1
+ vccd1 top.a1.dataIn\[0\] sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_39_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_464 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06598__A2 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12716__RESET_B net1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11307_ _05123_ _05130_ vssd1 vssd1 vccd1 vccd1 _05194_ sky130_fd_sc_hd__and2_1
X_12287_ top.lcd.cnt_500hz\[12\] _06101_ vssd1 vssd1 vccd1 vccd1 _06103_ sky130_fd_sc_hd__or2_1
X_11238_ net881 top.lcd.nextState\[0\] vssd1 vssd1 vccd1 vccd1 _05131_ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_52_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11169_ _01380_ _01418_ _01414_ _01410_ vssd1 vssd1 vccd1 vccd1 _05094_ sky130_fd_sc_hd__o211a_1
XFILLER_0_93_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06770__A2 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_wire413_A _02088_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_203_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_202_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06522__A2 net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07400_ top.DUT.register\[28\]\[9\] net555 net515 top.DUT.register\[7\]\[9\] vssd1
+ vssd1 vccd1 vccd1 _02539_ sky130_fd_sc_hd__a22o_1
XFILLER_0_9_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08380_ _02753_ net432 net426 _03501_ _03491_ vssd1 vssd1 vccd1 vccd1 _03513_ sky130_fd_sc_hd__a221o_1
XFILLER_0_92_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07331_ top.DUT.register\[5\]\[12\] net651 net766 top.DUT.register\[28\]\[12\] vssd1
+ vssd1 vccd1 vccd1 _02470_ sky130_fd_sc_hd__a22o_1
XFILLER_0_128_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12096__A top.a1.dataIn\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09389__B _04438_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_0_clk_X clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_190_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_236 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07483__B1 net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07262_ top.DUT.register\[23\]\[13\] net573 _02400_ vssd1 vssd1 vccd1 vccd1 _02401_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_183_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_450 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09001_ net282 _03381_ _03454_ _04075_ net435 vssd1 vssd1 vccd1 vccd1 _04076_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_171_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_154_2757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06213_ top.ramload\[7\] net856 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedInstr\[7\]
+ sky130_fd_sc_hd__and2_1
XANTENNA__09676__Y _04712_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07193_ _01392_ top.a1.instruction\[14\] vssd1 vssd1 vccd1 vccd1 _02332_ sky130_fd_sc_hd__or2_1
XFILLER_0_26_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07235__B1 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06144_ top.Ren vssd1 vssd1 vccd1 vccd1 _01387_ sky130_fd_sc_hd__inv_2
XANTENNA__09775__A2 net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06589__A2 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07786__A1 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_187_3245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_187_3256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09903_ _04909_ _04910_ vssd1 vssd1 vccd1 vccd1 _04911_ sky130_fd_sc_hd__and2_1
Xfanout503 _01567_ vssd1 vssd1 vccd1 vccd1 net503 sky130_fd_sc_hd__clkbuf_8
Xfanout514 _01559_ vssd1 vssd1 vccd1 vccd1 net514 sky130_fd_sc_hd__clkbuf_4
Xfanout525 net526 vssd1 vssd1 vccd1 vccd1 net525 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_6_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout395_A net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout536 _01541_ vssd1 vssd1 vccd1 vccd1 net536 sky130_fd_sc_hd__buf_4
Xfanout547 net550 vssd1 vssd1 vccd1 vccd1 net547 sky130_fd_sc_hd__clkbuf_8
X_09834_ _04845_ _04846_ _04848_ vssd1 vssd1 vccd1 vccd1 _04849_ sky130_fd_sc_hd__o21ai_1
Xfanout558 _01534_ vssd1 vssd1 vccd1 vccd1 net558 sky130_fd_sc_hd__buf_4
Xfanout569 _01525_ vssd1 vssd1 vccd1 vccd1 net569 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_206_3540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09765_ net799 _04786_ _04782_ vssd1 vssd1 vccd1 vccd1 _04787_ sky130_fd_sc_hd__a21o_1
X_06977_ top.DUT.register\[22\]\[23\] net649 net728 top.DUT.register\[18\]\[23\] _02115_
+ vssd1 vssd1 vccd1 vccd1 _02116_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout562_A _01532_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06761__A2 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08716_ _02092_ _03833_ vssd1 vssd1 vccd1 vccd1 _03834_ sky130_fd_sc_hd__xnor2_1
XANTENNA__11098__A1 net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09696_ net2076 net263 net631 vssd1 vssd1 vccd1 vccd1 _00123_ sky130_fd_sc_hd__mux2_1
XANTENNA__06269__A top.ramload\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08647_ _02266_ _03727_ _03767_ vssd1 vssd1 vccd1 vccd1 _03768_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout350_X net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_520 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06513__A2 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout827_A net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout448_X net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08578_ _03701_ _03702_ vssd1 vssd1 vccd1 vccd1 _03703_ sky130_fd_sc_hd__or2_1
XFILLER_0_166_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07529_ _02661_ _02663_ _02665_ _02667_ vssd1 vssd1 vccd1 vccd1 _02668_ sky130_fd_sc_hd__or4_1
XFILLER_0_76_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout615_X net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10540_ net2074 net230 net354 vssd1 vssd1 vccd1 vccd1 _00707_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10471_ net1833 net235 net361 vssd1 vssd1 vccd1 vccd1 _00641_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_157_Right_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12210_ top.lcd.cnt_20ms\[13\] top.lcd.cnt_20ms\[12\] top.lcd.cnt_20ms\[11\] top.lcd.cnt_20ms\[10\]
+ vssd1 vssd1 vccd1 vccd1 _06056_ sky130_fd_sc_hd__or4bb_1
X_13190_ clknet_leaf_40_clk _00782_ net1053 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[21\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09766__A2 net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_691 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12141_ _06018_ _06019_ vssd1 vssd1 vccd1 vccd1 _06024_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_94_1859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_208_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12072_ _05952_ _05954_ vssd1 vssd1 vccd1 vccd1 _05955_ sky130_fd_sc_hd__and2b_1
Xhold590 top.ramload\[18\] vssd1 vssd1 vccd1 vccd1 net1706 sky130_fd_sc_hd__dlygate4sd3_1
X_11023_ net33 net839 net817 net2072 vssd1 vssd1 vccd1 vccd1 _01135_ sky130_fd_sc_hd__o22a_1
XANTENNA__09762__B _04386_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07834__Y _02973_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07563__A net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06752__A2 net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12974_ clknet_leaf_40_clk _00566_ net1055 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[14\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_2_clk_X clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11925_ _05759_ _05760_ _05782_ vssd1 vssd1 vccd1 vccd1 _05808_ sky130_fd_sc_hd__and3_1
XFILLER_0_86_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_200_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11856_ _05722_ _05735_ vssd1 vssd1 vccd1 vccd1 _05739_ sky130_fd_sc_hd__nor2_1
XFILLER_0_129_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_200_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_184_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10807_ net188 net1756 net599 vssd1 vssd1 vccd1 vccd1 _00968_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_109_Left_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_145_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11787_ _05641_ _05669_ vssd1 vssd1 vccd1 vccd1 _05670_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_184_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_171_3013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_1988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10738_ net1551 net229 net418 vssd1 vssd1 vccd1 vccd1 _00899_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07465__B1 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13526_ clknet_leaf_74_clk top.a1.nextHex\[4\] net1077 vssd1 vssd1 vccd1 vccd1 _01380_
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10863__S net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13457_ clknet_leaf_112_clk _01049_ net988 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[30\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_10669_ net2071 net246 net338 vssd1 vssd1 vccd1 vccd1 _00832_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_124_Right_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_136_2487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12408_ clknet_leaf_109_clk top.ru.next_FetchedInstr\[20\] net975 vssd1 vssd1 vccd1
+ vccd1 top.a1.instruction\[20\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_113_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09757__A2 net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13388_ clknet_leaf_47_clk _00980_ net1093 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[27\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
Xoutput106 net106 vssd1 vssd1 vccd1 vccd1 SEL_O[1] sky130_fd_sc_hd__buf_2
Xoutput117 net117 vssd1 vssd1 vccd1 vccd1 gpio_out[19] sky130_fd_sc_hd__buf_2
X_12339_ net1233 _06134_ _06135_ vssd1 vssd1 vccd1 vccd1 _01366_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_118_Left_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_195_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06900_ top.DUT.register\[4\]\[18\] net669 net653 top.DUT.register\[5\]\[18\] vssd1
+ vssd1 vccd1 vccd1 _02039_ sky130_fd_sc_hd__a22o_1
X_07880_ _03011_ _03018_ vssd1 vssd1 vccd1 vccd1 _03019_ sky130_fd_sc_hd__nor2_4
XTAP_TAPCELL_ROW_182_3175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06831_ top.DUT.register\[25\]\[19\] net457 net509 top.DUT.register\[4\]\[19\] _01969_
+ vssd1 vssd1 vccd1 vccd1 _01970_ sky130_fd_sc_hd__a221o_1
XFILLER_0_208_787 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06743__A2 net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07940__A1 _02007_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09550_ _04597_ _04598_ vssd1 vssd1 vccd1 vccd1 _04599_ sky130_fd_sc_hd__or2_1
X_06762_ top.DUT.register\[23\]\[24\] net674 net716 top.DUT.register\[27\]\[24\] vssd1
+ vssd1 vccd1 vccd1 _01901_ sky130_fd_sc_hd__a22o_1
XANTENNA__10103__S net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08856__X _03968_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08501_ _03541_ _03628_ net313 vssd1 vssd1 vccd1 vccd1 _03629_ sky130_fd_sc_hd__mux2_1
XANTENNA_wire416_X net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09481_ net901 top.pc\[23\] _04534_ net891 vssd1 vssd1 vccd1 vccd1 _00103_ sky130_fd_sc_hd__o211a_1
X_06693_ _01809_ _01830_ vssd1 vssd1 vccd1 vccd1 _01832_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_65_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09693__A1 top.a1.dataIn\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08496__A2 net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08432_ _02524_ net431 net500 _02523_ _03562_ vssd1 vssd1 vccd1 vccd1 _03563_ sky130_fd_sc_hd__a221o_1
XFILLER_0_144_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08363_ _03364_ _03368_ net305 vssd1 vssd1 vccd1 vccd1 _03496_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout143_A _04946_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07314_ _02443_ _02452_ vssd1 vssd1 vccd1 vccd1 _02453_ sky130_fd_sc_hd__nor2_4
XFILLER_0_156_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07456__B1 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_63 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_620 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08294_ net426 _03410_ _03429_ net428 _03425_ vssd1 vssd1 vccd1 vccd1 _03430_ sky130_fd_sc_hd__a221o_2
XFILLER_0_116_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07245_ _02383_ vssd1 vssd1 vccd1 vccd1 _02384_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout310_A net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10773__S net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1052_A net1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11004__A1 top.a1.dataIn\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07176_ top.DUT.register\[8\]\[10\] net539 net519 top.DUT.register\[10\]\[10\] vssd1
+ vssd1 vccd1 vccd1 _02315_ sky130_fd_sc_hd__a22o_1
XFILLER_0_14_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08956__B1 _02472_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout300 net301 vssd1 vssd1 vccd1 vccd1 net300 sky130_fd_sc_hd__buf_2
Xfanout311 net314 vssd1 vssd1 vccd1 vccd1 net311 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_1_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_167_2948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06982__A2 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout322 net323 vssd1 vssd1 vccd1 vccd1 net322 sky130_fd_sc_hd__clkbuf_2
XANTENNA__10361__X _04981_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09582__B _04628_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout333 _03121_ vssd1 vssd1 vccd1 vccd1 net333 sky130_fd_sc_hd__buf_4
Xfanout344 _04992_ vssd1 vssd1 vccd1 vccd1 net344 sky130_fd_sc_hd__buf_8
Xfanout355 net356 vssd1 vssd1 vccd1 vccd1 net355 sky130_fd_sc_hd__clkbuf_8
Xfanout366 net367 vssd1 vssd1 vccd1 vccd1 net366 sky130_fd_sc_hd__clkbuf_8
Xfanout377 net380 vssd1 vssd1 vccd1 vccd1 net377 sky130_fd_sc_hd__buf_8
X_09817_ _04824_ _04827_ _04825_ vssd1 vssd1 vccd1 vccd1 _04833_ sky130_fd_sc_hd__a21o_1
Xfanout388 _04978_ vssd1 vssd1 vccd1 vccd1 net388 sky130_fd_sc_hd__buf_4
XANTENNA_fanout565_X net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout399 net400 vssd1 vssd1 vccd1 vccd1 net399 sky130_fd_sc_hd__buf_2
XANTENNA_fanout944_A net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06734__A2 net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07931__A1 _02580_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09748_ net1457 net212 net631 vssd1 vssd1 vccd1 vccd1 _00133_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_107_2044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_2055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10948__S net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09679_ _02340_ _04177_ vssd1 vssd1 vccd1 vccd1 _04715_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout732_X net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11710_ _05553_ _05581_ _05557_ vssd1 vssd1 vccd1 vccd1 _05593_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_68_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07695__B1 net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12690_ clknet_leaf_24_clk _00282_ net1012 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[6\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_120_2244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11641_ top.a1.dataIn\[12\] _05514_ _05515_ vssd1 vssd1 vccd1 vccd1 _05524_ sky130_fd_sc_hd__and3_1
XFILLER_0_64_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_166_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07447__B1 net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11572_ _05425_ net249 _05428_ vssd1 vssd1 vccd1 vccd1 _05455_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08942__A net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13311_ clknet_leaf_24_clk _00903_ net1013 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[25\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_10523_ net1339 net159 net359 vssd1 vssd1 vccd1 vccd1 _00692_ sky130_fd_sc_hd__mux2_1
Xinput19 DAT_I[25] vssd1 vssd1 vccd1 vccd1 net19 sky130_fd_sc_hd__clkbuf_1
XANTENNA__10683__S net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13242_ clknet_leaf_3_clk _00834_ net917 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[23\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10454_ net173 net2098 net366 vssd1 vssd1 vccd1 vccd1 _00625_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08947__B1 _02878_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_423 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13173_ clknet_leaf_31_clk _00765_ net1020 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[21\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10385_ net2070 net177 net375 vssd1 vssd1 vccd1 vccd1 _00560_ sky130_fd_sc_hd__mux2_1
X_12124_ _06006_ vssd1 vssd1 vccd1 vccd1 _06007_ sky130_fd_sc_hd__inv_2
XFILLER_0_130_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12055_ _05909_ _05918_ _05937_ vssd1 vssd1 vccd1 vccd1 _05938_ sky130_fd_sc_hd__and3_1
XANTENNA__07564__Y _02703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09492__B _01896_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11006_ top.a1.data\[7\] net783 vssd1 vssd1 vccd1 vccd1 _05038_ sky130_fd_sc_hd__or2_1
XANTENNA__06186__A0 net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06725__A2 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11246__C _05120_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_158_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10858__S net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12957_ clknet_leaf_119_clk _00549_ net930 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[14\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06908__Y _02047_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11908_ _05759_ _05786_ _05779_ vssd1 vssd1 vccd1 vccd1 _05791_ sky130_fd_sc_hd__or3b_2
XANTENNA__11482__A1 top.a1.dataIn\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07686__B1 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_47_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12888_ clknet_leaf_125_clk _00480_ net923 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[12\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_47_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07150__A2 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_56 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11839_ _05704_ _05720_ _05721_ vssd1 vssd1 vccd1 vccd1 _05722_ sky130_fd_sc_hd__a21boi_2
XTAP_TAPCELL_ROW_138_2516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07438__B1 net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13509_ clknet_leaf_33_clk _01101_ net1046 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[31\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07739__Y _02878_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10593__S net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_151_2705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_151_2716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07030_ top.DUT.register\[23\]\[20\] net673 _02166_ _02168_ vssd1 vssd1 vccd1 vccd1
+ _02169_ sky130_fd_sc_hd__a211o_1
XFILLER_0_125_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_141_734 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_184_3204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08981_ _04055_ _03703_ _03668_ _03661_ vssd1 vssd1 vccd1 vccd1 _04056_ sky130_fd_sc_hd__and4b_1
XANTENNA__06964__A2 net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07932_ _02623_ _02632_ _02653_ vssd1 vssd1 vccd1 vccd1 _03071_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_149_2678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07863_ top.DUT.register\[10\]\[1\] net772 net708 top.DUT.register\[15\]\[1\] vssd1
+ vssd1 vccd1 vccd1 _03002_ sky130_fd_sc_hd__a22o_1
XANTENNA__06716__A2 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07913__A1 net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06814_ top.DUT.register\[21\]\[17\] net656 net751 top.DUT.register\[26\]\[17\] vssd1
+ vssd1 vccd1 vccd1 _01953_ sky130_fd_sc_hd__a22o_1
X_09602_ _04636_ _04637_ vssd1 vssd1 vccd1 vccd1 _04648_ sky130_fd_sc_hd__nand2b_1
X_07794_ top.DUT.register\[23\]\[2\] net571 net519 top.DUT.register\[10\]\[2\] _02932_
+ vssd1 vssd1 vccd1 vccd1 _02933_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_162_2878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09533_ net900 top.pc\[26\] _04570_ _04583_ net890 vssd1 vssd1 vccd1 vccd1 _00106_
+ sky130_fd_sc_hd__o221a_1
X_06745_ top.DUT.register\[26\]\[24\] net529 net449 top.DUT.register\[21\]\[24\] _01883_
+ vssd1 vssd1 vccd1 vccd1 _01884_ sky130_fd_sc_hd__a221o_1
XANTENNA__09666__A1 top.pc\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10768__S net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout260_A net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout358_A net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09464_ net133 _04513_ _04517_ _04518_ net901 vssd1 vssd1 vccd1 vccd1 _04519_ sky130_fd_sc_hd__o221a_1
XANTENNA__07677__B1 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06676_ top.DUT.register\[26\]\[26\] net753 net748 top.DUT.register\[17\]\[26\] _01814_
+ vssd1 vssd1 vccd1 vccd1 _01815_ sky130_fd_sc_hd__a221o_1
XFILLER_0_78_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_195_3366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13308__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07141__A2 net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_195_3377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08415_ net498 _03523_ _03532_ _03258_ _03546_ vssd1 vssd1 vccd1 vccd1 _03547_ sky130_fd_sc_hd__o221a_1
XFILLER_0_175_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_35_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12819__RESET_B net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09418__A1 net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09395_ _02016_ _02025_ _04453_ vssd1 vssd1 vccd1 vccd1 _04454_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout525_A net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09418__B2 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_175_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06266__B net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08346_ net302 _03327_ vssd1 vssd1 vccd1 vccd1 _03480_ sky130_fd_sc_hd__nor2_1
XFILLER_0_19_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_550 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08277_ _03411_ _03412_ vssd1 vssd1 vccd1 vccd1 _03413_ sky130_fd_sc_hd__and2_2
XTAP_TAPCELL_ROW_78_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12401__RESET_B net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_723 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07228_ top.DUT.register\[7\]\[10\] net659 net742 top.DUT.register\[2\]\[10\] vssd1
+ vssd1 vccd1 vccd1 _02367_ sky130_fd_sc_hd__a22o_1
XFILLER_0_89_80 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10008__S net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07159_ top.DUT.register\[25\]\[11\] net778 net643 top.DUT.register\[24\]\[11\] _02297_
+ vssd1 vssd1 vccd1 vccd1 _02298_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_91_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10170_ net1327 net172 net604 vssd1 vssd1 vccd1 vccd1 _00369_ sky130_fd_sc_hd__mux2_1
XFILLER_0_112_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout682_X net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06955__A2 net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_6_0_clk_X clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout141 net143 vssd1 vssd1 vccd1 vccd1 net141 sky130_fd_sc_hd__clkbuf_2
Xfanout152 _04929_ vssd1 vssd1 vccd1 vccd1 net152 sky130_fd_sc_hd__clkbuf_2
Xfanout174 _04876_ vssd1 vssd1 vccd1 vccd1 net174 sky130_fd_sc_hd__buf_2
XANTENNA__11161__A0 top.a1.row1\[57\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout185 net187 vssd1 vssd1 vccd1 vccd1 net185 sky130_fd_sc_hd__clkbuf_2
XANTENNA__06707__A2 net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout196 _04788_ vssd1 vssd1 vccd1 vccd1 net196 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07380__A2 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12811_ clknet_leaf_48_clk _00403_ net1060 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[9\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10678__S net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13791_ clknet_leaf_68_clk _01360_ vssd1 vssd1 vccd1 vccd1 top.pad.button_control.r_counter\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_96_220 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12742_ clknet_leaf_33_clk _00334_ net1046 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[7\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09121__A3 _02943_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07132__A2 net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_69_Right_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_182_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12673_ clknet_leaf_19_clk _00265_ net1026 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[5\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_528 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11624_ _05503_ _05506_ _05501_ vssd1 vssd1 vccd1 vccd1 _05507_ sky130_fd_sc_hd__a21o_1
XFILLER_0_181_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_1947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08672__A net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11555_ _05394_ _05434_ vssd1 vssd1 vccd1 vccd1 _05438_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_42_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10506_ net1815 net229 net357 vssd1 vssd1 vccd1 vccd1 _00675_ sky130_fd_sc_hd__mux2_1
XFILLER_0_162_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07840__B1 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_2435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11486_ _05367_ _05368_ vssd1 vssd1 vccd1 vccd1 _05369_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_133_2446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13225_ clknet_leaf_52_clk _00817_ net1039 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[22\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_10437_ net245 net2166 net365 vssd1 vssd1 vccd1 vccd1 _00608_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_78_Right_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13156_ clknet_leaf_37_clk _00748_ net1051 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[20\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10368_ net2271 net242 net373 vssd1 vssd1 vccd1 vccd1 _00543_ sky130_fd_sc_hd__mux2_1
XANTENNA__06946__A2 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12107_ _05965_ _05969_ vssd1 vssd1 vccd1 vccd1 _05990_ sky130_fd_sc_hd__xnor2_1
X_13087_ clknet_leaf_20_clk _00679_ net1028 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[18\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12975__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10299_ net259 net2142 net382 vssd1 vssd1 vccd1 vccd1 _00476_ sky130_fd_sc_hd__mux2_1
X_12038_ _05871_ _05910_ vssd1 vssd1 vccd1 vccd1 _05921_ sky130_fd_sc_hd__or2_1
XANTENNA__09896__A1 _04150_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07371__A2 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10588__S net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_87_Right_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06530_ top.DUT.register\[15\]\[29\] net681 net677 top.DUT.register\[31\]\[29\] vssd1
+ vssd1 vccd1 vccd1 _01669_ sky130_fd_sc_hd__a22o_1
XFILLER_0_87_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07123__A2 net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08320__A1 net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08320__B2 net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06461_ top.a1.instruction\[22\] top.a1.instruction\[23\] net792 vssd1 vssd1 vccd1
+ vccd1 _01600_ sky130_fd_sc_hd__and3b_2
XTAP_TAPCELL_ROW_177_3096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08200_ _03159_ _03182_ vssd1 vssd1 vccd1 vccd1 _03338_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_32_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09180_ net900 top.pc\[5\] _04244_ _04251_ net890 vssd1 vssd1 vccd1 vccd1 _00085_
+ sky130_fd_sc_hd__o221a_1
X_06392_ top.a1.instruction\[17\] top.a1.instruction\[18\] net782 vssd1 vssd1 vccd1
+ vccd1 _01531_ sky130_fd_sc_hd__o21ai_4
X_08131_ net1476 net833 _03268_ net803 vssd1 vssd1 vccd1 vccd1 _00018_ sky130_fd_sc_hd__a22o_1
XFILLER_0_71_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_190_3296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08062_ _01853_ net327 vssd1 vssd1 vccd1 vccd1 _03201_ sky130_fd_sc_hd__nand2_1
XFILLER_0_172_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07831__B1 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07013_ top.DUT.register\[23\]\[20\] net574 net509 top.DUT.register\[4\]\[20\] vssd1
+ vssd1 vccd1 vccd1 _02152_ sky130_fd_sc_hd__a22o_1
XFILLER_0_3_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_96_Right_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08638__A1_N _03264_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09677__A_N top.a1.instruction\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12183__A2 net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_72 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06398__B1 net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06937__A2 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08964_ _02175_ net691 net1166 net874 vssd1 vssd1 vccd1 vccd1 _00070_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_164_2907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1015_A net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07915_ _02773_ _02799_ _03053_ vssd1 vssd1 vccd1 vccd1 _03054_ sky130_fd_sc_hd__o21a_1
X_08895_ _01702_ _03097_ vssd1 vssd1 vccd1 vccd1 _04005_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout475_A net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07846_ top.DUT.register\[15\]\[0\] net679 net675 top.DUT.register\[31\]\[0\] vssd1
+ vssd1 vccd1 vccd1 _02985_ sky130_fd_sc_hd__a22o_1
XANTENNA__07898__B1 net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_197_3406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08757__A net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07362__A2 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_2003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07661__A _02773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07777_ top.DUT.register\[25\]\[2\] net779 net722 top.DUT.register\[29\]\[2\] vssd1
+ vssd1 vccd1 vccd1 _02916_ sky130_fd_sc_hd__a22o_1
XANTENNA__10498__S net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06570__B1 net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout642_A _01619_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06728_ top.DUT.register\[15\]\[25\] net706 net698 top.DUT.register\[31\]\[25\] vssd1
+ vssd1 vccd1 vccd1 _01867_ sky130_fd_sc_hd__a22o_1
X_09516_ top.pc\[26\] _04556_ vssd1 vssd1 vccd1 vccd1 _04567_ sky130_fd_sc_hd__and2_1
XFILLER_0_195_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07114__A2 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09447_ _04498_ _04502_ vssd1 vssd1 vccd1 vccd1 _04503_ sky130_fd_sc_hd__xnor2_1
X_06659_ top.DUT.register\[20\]\[26\] net565 net557 top.DUT.register\[28\]\[26\] _01797_
+ vssd1 vssd1 vccd1 vccd1 _01798_ sky130_fd_sc_hd__a221o_1
XFILLER_0_164_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout430_X net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout528_X net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout907_A net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_164_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09378_ net805 _02726_ _04335_ _04437_ vssd1 vssd1 vccd1 vccd1 _04438_ sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_163_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08329_ _03053_ _03462_ vssd1 vssd1 vccd1 vccd1 _03463_ sky130_fd_sc_hd__nand2_1
XFILLER_0_117_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06283__Y _01446_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_163_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11340_ _05221_ _05222_ vssd1 vssd1 vccd1 vccd1 _05223_ sky130_fd_sc_hd__and2_1
XANTENNA__07822__B1 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout897_X net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11271_ top.a1.row1\[10\] _05126_ _05136_ top.a1.row1\[58\] _05153_ vssd1 vssd1 vccd1
+ vccd1 _05162_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_115_2165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_2176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13010_ clknet_leaf_23_clk _00602_ net1015 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[16\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12174__A2 net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10222_ net170 net1812 net393 vssd1 vssd1 vccd1 vccd1 _00402_ sky130_fd_sc_hd__mux2_1
XANTENNA__06928__A2 net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10153_ net1586 net247 net602 vssd1 vssd1 vccd1 vccd1 _00352_ sky130_fd_sc_hd__mux2_1
XANTENNA__10262__A _04155_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input36_A gpio_in[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10084_ net1467 net258 net613 vssd1 vssd1 vccd1 vccd1 _00285_ sky130_fd_sc_hd__mux2_1
Xhold8 top.a1.dataInTemp\[3\] vssd1 vssd1 vccd1 vccd1 net1124 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07889__B1 net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07353__A2 net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_199_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10201__S net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13774_ clknet_leaf_100_clk _01345_ vssd1 vssd1 vccd1 vccd1 top.lcd.cnt_500hz\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_10986_ net1164 _05023_ net589 vssd1 vssd1 vccd1 vccd1 _01119_ sky130_fd_sc_hd__mux2_1
XANTENNA__06187__A net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07105__A2 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12725_ clknet_leaf_31_clk _00317_ net1023 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[7\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12656_ clknet_leaf_29_clk _00248_ net1017 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[4\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_684 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_615 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11607_ net234 _05476_ _05453_ vssd1 vssd1 vccd1 vccd1 _05490_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07289__Y _02428_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12587_ clknet_leaf_45_clk _00179_ net1065 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[2\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09785__X _04805_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11538_ _05419_ _05420_ vssd1 vssd1 vccd1 vccd1 _05421_ sky130_fd_sc_hd__nand2_1
XFILLER_0_111_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold408 top.DUT.register\[2\]\[26\] vssd1 vssd1 vccd1 vccd1 net1524 sky130_fd_sc_hd__dlygate4sd3_1
Xhold419 top.DUT.register\[27\]\[27\] vssd1 vssd1 vccd1 vccd1 net1535 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap127 _05836_ vssd1 vssd1 vccd1 vccd1 net127 sky130_fd_sc_hd__buf_1
XFILLER_0_52_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11469_ _05274_ _05315_ _05345_ vssd1 vssd1 vccd1 vccd1 _05352_ sky130_fd_sc_hd__and3_1
XANTENNA__10871__S net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13208_ clknet_leaf_128_clk _00800_ net912 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[22\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_96_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06919__A2 net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_584 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13139_ clknet_leaf_123_clk _00731_ net927 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[20\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_55_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07592__A2 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13153__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1108 top.DUT.register\[11\]\[1\] vssd1 vssd1 vccd1 vccd1 net2224 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1119 top.DUT.register\[9\]\[22\] vssd1 vssd1 vccd1 vccd1 net2235 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_146_2637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07700_ _02832_ _02834_ _02836_ _02838_ vssd1 vssd1 vccd1 vccd1 _02839_ sky130_fd_sc_hd__or4_4
XFILLER_0_206_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08680_ _02005_ _03185_ _03187_ _02006_ vssd1 vssd1 vccd1 vccd1 _03800_ sky130_fd_sc_hd__o22a_1
XANTENNA__07344__A2 net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07631_ top.DUT.register\[20\]\[5\] net563 net443 top.DUT.register\[1\]\[5\] vssd1
+ vssd1 vccd1 vccd1 _02770_ sky130_fd_sc_hd__a22o_1
XFILLER_0_178_715 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_179_3125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_179_3136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06552__B1 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_177_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07562_ _02693_ _02700_ vssd1 vssd1 vccd1 vccd1 _02701_ sky130_fd_sc_hd__or2_4
XANTENNA__10111__S net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_177_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09301_ _04363_ _04364_ vssd1 vssd1 vccd1 vccd1 _04365_ sky130_fd_sc_hd__or2_1
X_06513_ top.DUT.register\[18\]\[30\] net728 net724 top.DUT.register\[29\]\[30\] vssd1
+ vssd1 vccd1 vccd1 _01652_ sky130_fd_sc_hd__a22o_1
XFILLER_0_193_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_192_3325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07493_ _02625_ _02627_ _02629_ _02631_ vssd1 vssd1 vccd1 vccd1 _02632_ sky130_fd_sc_hd__or4_4
XFILLER_0_152_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09232_ top.pc\[9\] _02502_ vssd1 vssd1 vccd1 vccd1 _04300_ sky130_fd_sc_hd__and2b_1
X_06444_ net805 _01582_ vssd1 vssd1 vccd1 vccd1 _01583_ sky130_fd_sc_hd__or2_2
XFILLER_0_91_716 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_824 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_95 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_144 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_667 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09201__A net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_183 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09163_ _01393_ _04224_ _04234_ _04235_ vssd1 vssd1 vccd1 vccd1 _00084_ sky130_fd_sc_hd__o31a_1
X_06375_ top.a1.instruction\[17\] top.a1.instruction\[18\] net684 _01512_ vssd1 vssd1
+ vccd1 vccd1 _01514_ sky130_fd_sc_hd__and4_4
XFILLER_0_44_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_157_2799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout223_A _04805_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08114_ _03251_ _03252_ vssd1 vssd1 vccd1 vccd1 _03253_ sky130_fd_sc_hd__and2_1
XFILLER_0_32_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_142 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_339 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_462 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09695__X _04729_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_211_3620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09094_ net895 _01478_ _03148_ _04168_ _02337_ vssd1 vssd1 vccd1 vccd1 _04169_ sky130_fd_sc_hd__o311a_1
XTAP_TAPCELL_ROW_211_3631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08045_ _03181_ _03182_ vssd1 vssd1 vccd1 vccd1 _03184_ sky130_fd_sc_hd__nor2_1
XANTENNA__10781__S net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold920 top.DUT.register\[31\]\[8\] vssd1 vssd1 vccd1 vccd1 net2036 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_170_2999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold931 top.DUT.register\[12\]\[9\] vssd1 vssd1 vccd1 vccd1 net2047 sky130_fd_sc_hd__dlygate4sd3_1
Xhold942 top.DUT.register\[3\]\[0\] vssd1 vssd1 vccd1 vccd1 net2058 sky130_fd_sc_hd__dlygate4sd3_1
Xhold953 top.DUT.register\[9\]\[30\] vssd1 vssd1 vccd1 vccd1 net2069 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06560__A _01678_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold964 top.DUT.register\[21\]\[14\] vssd1 vssd1 vccd1 vccd1 net2080 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout592_A _04971_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold975 top.DUT.register\[13\]\[2\] vssd1 vssd1 vccd1 vccd1 net2091 sky130_fd_sc_hd__dlygate4sd3_1
Xhold986 top.DUT.register\[1\]\[22\] vssd1 vssd1 vccd1 vccd1 net2102 sky130_fd_sc_hd__dlygate4sd3_1
Xhold997 top.DUT.register\[12\]\[25\] vssd1 vssd1 vccd1 vccd1 net2113 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_86_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09996_ net223 net1849 net623 vssd1 vssd1 vccd1 vccd1 _00201_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_110_2095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_209_3582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08947_ net1297 net876 _02878_ net693 vssd1 vssd1 vccd1 vccd1 _00053_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout380_X net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout857_A top.ru.next_iready vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout478_X net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_84_clk_A clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09590__B _04620_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08878_ _03969_ _03987_ vssd1 vssd1 vccd1 vccd1 _03989_ sky130_fd_sc_hd__and2_1
XANTENNA__07335__A2 _02452_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07829_ top.DUT.register\[28\]\[0\] net766 net762 top.DUT.register\[9\]\[0\] vssd1
+ vssd1 vccd1 vccd1 _02968_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_86_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06543__B1 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout645_X net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10021__S net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10840_ net1820 net225 net475 vssd1 vssd1 vccd1 vccd1 _01001_ sky130_fd_sc_hd__mux2_1
XANTENNA__08774__X _03890_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_211_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_426 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_99_clk_A clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10771_ net2046 net219 net482 vssd1 vssd1 vccd1 vccd1 _00932_ sky130_fd_sc_hd__mux2_1
XFILLER_0_177_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout812_X net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_623 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11641__A top.a1.dataIn\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12510_ clknet_leaf_78_clk _00102_ net1074 vssd1 vssd1 vccd1 vccd1 top.pc\[22\] sky130_fd_sc_hd__dfrtp_4
X_13490_ clknet_leaf_23_clk _01082_ net1015 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[31\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06735__A _01853_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09111__A top.pc\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_2205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12441_ clknet_leaf_75_clk _00037_ net1081 vssd1 vssd1 vccd1 vccd1 top.ramaddr\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_22_clk_A clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08599__A1 _03342_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08599__B2 net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12372_ clknet_leaf_105_clk top.ru.next_FetchedData\[16\] net973 vssd1 vssd1 vccd1
+ vccd1 top.a1.dataIn\[16\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_90_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06173__C top.a1.halfData\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11323_ top.a1.dataIn\[18\] top.a1.dataIn\[19\] top.a1.dataIn\[17\] top.a1.dataIn\[16\]
+ vssd1 vssd1 vccd1 vccd1 _05206_ sky130_fd_sc_hd__nor4_1
XANTENNA__10691__S net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_37_clk_A clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11254_ top.a1.row2\[16\] _05145_ _05146_ top.a1.row2\[40\] vssd1 vssd1 vccd1 vccd1
+ _05147_ sky130_fd_sc_hd__a22o_1
X_10205_ net237 top.DUT.register\[9\]\[8\] net396 vssd1 vssd1 vccd1 vccd1 _00385_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11185_ net1995 net588 _04668_ vssd1 vssd1 vccd1 vccd1 _01242_ sky130_fd_sc_hd__a21o_1
XANTENNA__09781__A net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10136_ net176 net2097 net608 vssd1 vssd1 vccd1 vccd1 _00336_ sky130_fd_sc_hd__mux2_1
X_10067_ net1343 net202 net618 vssd1 vssd1 vccd1 vccd1 _00269_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_128_2367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07326__A2 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09720__B1 net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_50_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06534__B1 net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_5__f_clk_A clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload1_A clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12504__RESET_B net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_141_2556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13826_ net1110 vssd1 vssd1 vccd1 vccd1 gpio_out[25] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_141_2567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06348__C net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_175_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10866__S net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13757_ clknet_leaf_99_clk _01328_ vssd1 vssd1 vccd1 vccd1 top.lcd.cnt_20ms\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_10969_ net1159 _05010_ net590 vssd1 vssd1 vccd1 vccd1 _01115_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12708_ clknet_leaf_36_clk _00300_ net1051 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[6\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_174_3055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13688_ clknet_leaf_71_clk _00000_ vssd1 vssd1 vccd1 vccd1 top.lcd.nextState\[0\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_31_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12639_ clknet_leaf_19_clk _00231_ net1026 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[4\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_110_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06160_ top.a1.dataIn\[1\] vssd1 vssd1 vccd1 vccd1 _01403_ sky130_fd_sc_hd__inv_2
XFILLER_0_142_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_198_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13519__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_57_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold205 top.DUT.register\[25\]\[9\] vssd1 vssd1 vccd1 vccd1 net1321 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06651__Y _01790_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold216 top.DUT.register\[11\]\[16\] vssd1 vssd1 vccd1 vccd1 net1332 sky130_fd_sc_hd__dlygate4sd3_1
Xhold227 top.DUT.register\[5\]\[20\] vssd1 vssd1 vccd1 vccd1 net1343 sky130_fd_sc_hd__dlygate4sd3_1
Xhold238 top.DUT.register\[30\]\[22\] vssd1 vssd1 vccd1 vccd1 net1354 sky130_fd_sc_hd__dlygate4sd3_1
Xhold249 top.DUT.register\[18\]\[0\] vssd1 vssd1 vccd1 vccd1 net1365 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10106__S net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09850_ top.pc\[23\] _01584_ vssd1 vssd1 vccd1 vccd1 _04863_ sky130_fd_sc_hd__nand2_1
Xfanout707 _01640_ vssd1 vssd1 vccd1 vccd1 net707 sky130_fd_sc_hd__buf_2
Xfanout718 _01635_ vssd1 vssd1 vccd1 vccd1 net718 sky130_fd_sc_hd__clkbuf_8
Xfanout729 _01628_ vssd1 vssd1 vccd1 vccd1 net729 sky130_fd_sc_hd__clkbuf_4
X_08801_ _03300_ _03317_ vssd1 vssd1 vccd1 vccd1 _03915_ sky130_fd_sc_hd__nand2_1
X_06993_ net807 _02131_ net437 vssd1 vssd1 vccd1 vccd1 _02132_ sky130_fd_sc_hd__o21ai_1
X_09781_ net827 _04412_ vssd1 vssd1 vccd1 vccd1 _04801_ sky130_fd_sc_hd__nor2_1
XFILLER_0_147_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06773__B1 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_51 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08732_ net1304 net831 net801 _03849_ vssd1 vssd1 vccd1 vccd1 _00039_ sky130_fd_sc_hd__a22o_1
XANTENNA__07317__A2 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08663_ _03783_ vssd1 vssd1 vccd1 vccd1 _03784_ sky130_fd_sc_hd__inv_2
XANTENNA__08100__A net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06525__B1 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout173_A _04876_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07614_ _02752_ vssd1 vssd1 vccd1 vccd1 _02753_ sky130_fd_sc_hd__inv_2
X_08594_ net320 _03717_ vssd1 vssd1 vccd1 vccd1 _03718_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_68_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_159_2828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07545_ top.DUT.register\[13\]\[7\] net774 net758 top.DUT.register\[30\]\[7\] vssd1
+ vssd1 vccd1 vccd1 _02684_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_127_clk clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_127_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_48_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10776__S net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_138_Right_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout340_A _04993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1082_A net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout438_A _01587_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07476_ top.DUT.register\[8\]\[14\] net541 net510 top.DUT.register\[4\]\[14\] vssd1
+ vssd1 vccd1 vccd1 _02615_ sky130_fd_sc_hd__a22o_1
XFILLER_0_174_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06427_ net683 _01516_ _01523_ vssd1 vssd1 vccd1 vccd1 _01566_ sky130_fd_sc_hd__and3_4
X_09215_ top.pc\[8\] _04268_ vssd1 vssd1 vccd1 vccd1 _04284_ sky130_fd_sc_hd__and2_1
XFILLER_0_106_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_174_795 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout605_A net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_20_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09146_ _01505_ _04218_ _04219_ _04215_ _01393_ vssd1 vssd1 vccd1 vccd1 _04220_ sky130_fd_sc_hd__a311o_1
X_06358_ _01491_ _01495_ _01496_ _01497_ vssd1 vssd1 vccd1 vccd1 _01498_ sky130_fd_sc_hd__or4_1
XANTENNA__13199__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08770__A _03121_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09077_ net894 _01477_ _03156_ vssd1 vssd1 vccd1 vccd1 _04152_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_102_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06289_ _01447_ _01448_ vssd1 vssd1 vccd1 vccd1 _01449_ sky130_fd_sc_hd__nor2_1
XANTENNA__13033__RESET_B net1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_2124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08028_ _03152_ _03158_ vssd1 vssd1 vccd1 vccd1 _03167_ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_96_1890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold750 top.DUT.register\[7\]\[19\] vssd1 vssd1 vccd1 vccd1 net1866 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout974_A net1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout595_X net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold761 top.DUT.register\[27\]\[22\] vssd1 vssd1 vccd1 vccd1 net1877 sky130_fd_sc_hd__dlygate4sd3_1
Xhold772 top.DUT.register\[13\]\[20\] vssd1 vssd1 vccd1 vccd1 net1888 sky130_fd_sc_hd__dlygate4sd3_1
Xhold783 top.DUT.register\[11\]\[27\] vssd1 vssd1 vccd1 vccd1 net1899 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10016__S net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold794 top.DUT.register\[3\]\[30\] vssd1 vssd1 vccd1 vccd1 net1910 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07556__A2 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08753__B2 _03869_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout762_X net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09979_ net690 _04712_ _04949_ vssd1 vssd1 vccd1 vccd1 _04951_ sky130_fd_sc_hd__and3_1
XANTENNA__06764__B1 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12990_ clknet_leaf_21_clk _00582_ net1033 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[15\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07308__A2 net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11104__A3 _01428_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09106__A _04172_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11941_ _05794_ _05822_ _05790_ vssd1 vssd1 vccd1 vccd1 _05824_ sky130_fd_sc_hd__a21o_1
X_11872_ _05753_ _05754_ vssd1 vssd1 vccd1 vccd1 _05755_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_28_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_157_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13611_ clknet_leaf_89_clk _01198_ net1002 vssd1 vssd1 vccd1 vccd1 net68 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_123_2286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10686__S net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_2297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10823_ net140 net1664 net601 vssd1 vssd1 vccd1 vccd1 _00984_ sky130_fd_sc_hd__mux2_1
XFILLER_0_184_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_118_clk clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_118_clk
+ sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_105_Right_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_267 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13542_ clknet_leaf_94_clk _01129_ net982 vssd1 vssd1 vccd1 vccd1 top.ramload\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_10754_ net1454 net164 net420 vssd1 vssd1 vccd1 vccd1 _00915_ sky130_fd_sc_hd__mux2_1
XANTENNA__09481__A2 top.pc\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13803__RESET_B net1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13473_ clknet_leaf_16_clk _01065_ net960 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[30\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_10685_ net1360 net179 net339 vssd1 vssd1 vccd1 vccd1 _00848_ sky130_fd_sc_hd__mux2_1
XFILLER_0_180_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12424_ clknet_leaf_87_clk _00020_ net1004 vssd1 vssd1 vccd1 vccd1 top.ramaddr\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_50_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12355_ clknet_leaf_94_clk top.ru.next_dready net982 vssd1 vssd1 vccd1 vccd1 top.d_ready
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_105_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11306_ net1170 net813 _05193_ net1082 vssd1 vssd1 vccd1 vccd1 _01269_ sky130_fd_sc_hd__o211a_1
X_12286_ top.lcd.cnt_500hz\[11\] _06100_ _06102_ net687 vssd1 vssd1 vccd1 vccd1 _01346_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_120_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11237_ net881 top.lcd.nextState\[0\] vssd1 vssd1 vccd1 vccd1 _05130_ sky130_fd_sc_hd__nor2_2
XANTENNA__11249__C _01382_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07547__A2 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08744__B2 net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11168_ top.a1.row1\[61\] _05085_ _05093_ vssd1 vssd1 vccd1 vccd1 _01231_ sky130_fd_sc_hd__o21a_1
XANTENNA__08398__Y _03530_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06755__B1 net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08839__B _03950_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10119_ net241 net2103 net607 vssd1 vssd1 vccd1 vccd1 _00319_ sky130_fd_sc_hd__mux2_1
X_11099_ net71 net865 vssd1 vssd1 vccd1 vccd1 _05055_ sky130_fd_sc_hd__and2_1
XFILLER_0_158_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13809_ net72 vssd1 vssd1 vccd1 vccd1 net106 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_202_184 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_109_clk clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_109_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__10596__S net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07330_ top.DUT.register\[23\]\[12\] net671 net663 top.DUT.register\[20\]\[12\] vssd1
+ vssd1 vccd1 vccd1 _02469_ sky130_fd_sc_hd__a22o_1
XFILLER_0_45_204 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06375__A top.a1.instruction\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07261_ top.DUT.register\[15\]\[13\] net681 net677 top.DUT.register\[31\]\[13\] vssd1
+ vssd1 vccd1 vccd1 _02400_ sky130_fd_sc_hd__a22o_1
XFILLER_0_45_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08680__B1 _03187_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_568 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09000_ net284 _03332_ _03176_ vssd1 vssd1 vccd1 vccd1 _04075_ sky130_fd_sc_hd__a21oi_1
X_06212_ net1245 net859 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedInstr\[6\] sky130_fd_sc_hd__and2_1
XANTENNA__10328__C net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_3_7_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_3_7_0_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_154_2758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07192_ _01486_ _01588_ vssd1 vssd1 vccd1 vccd1 _02331_ sky130_fd_sc_hd__nor2_1
XFILLER_0_171_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06143_ top.Wen vssd1 vssd1 vccd1 vccd1 _01386_ sky130_fd_sc_hd__inv_2
XFILLER_0_131_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08432__B1 net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_187_3246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07786__A2 _02904_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_187_3257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09902_ _04897_ _04899_ _04898_ vssd1 vssd1 vccd1 vccd1 _04910_ sky130_fd_sc_hd__a21o_1
XFILLER_0_6_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout504 _01567_ vssd1 vssd1 vccd1 vccd1 net504 sky130_fd_sc_hd__clkbuf_4
Xfanout515 _01558_ vssd1 vssd1 vccd1 vccd1 net515 sky130_fd_sc_hd__clkbuf_8
XANTENNA__07493__X _02632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09932__B1 net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout526 _01554_ vssd1 vssd1 vccd1 vccd1 net526 sky130_fd_sc_hd__buf_4
X_09833_ net828 _04493_ _04847_ vssd1 vssd1 vccd1 vccd1 _04848_ sky130_fd_sc_hd__o21ba_1
Xfanout537 net538 vssd1 vssd1 vccd1 vccd1 net537 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_67_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout548 net550 vssd1 vssd1 vccd1 vccd1 net548 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout290_A net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout559 _01532_ vssd1 vssd1 vccd1 vccd1 net559 sky130_fd_sc_hd__clkbuf_8
XANTENNA__06746__B1 net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_207_Right_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_206_3530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout388_A _04978_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_206_3541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09764_ _04783_ _04784_ vssd1 vssd1 vccd1 vccd1 _04786_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_198_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06976_ top.DUT.register\[8\]\[23\] net640 net703 top.DUT.register\[3\]\[23\] vssd1
+ vssd1 vccd1 vccd1 _02115_ sky130_fd_sc_hd__a22o_1
X_08715_ _02156_ _02176_ _03814_ vssd1 vssd1 vccd1 vccd1 _03833_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11175__B net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09695_ _03391_ net403 net488 _04728_ vssd1 vssd1 vccd1 vccd1 _04729_ sky130_fd_sc_hd__o211a_2
XANTENNA_fanout555_A net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06269__B net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08646_ _01963_ _02263_ vssd1 vssd1 vccd1 vccd1 _03767_ sky130_fd_sc_hd__nor2_1
XFILLER_0_194_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_194_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_532 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout722_A _01630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout343_X net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08577_ _02657_ _03700_ vssd1 vssd1 vccd1 vccd1 _03702_ sky130_fd_sc_hd__and2_1
XFILLER_0_193_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07528_ top.DUT.register\[16\]\[7\] net543 net527 top.DUT.register\[26\]\[7\] _02666_
+ vssd1 vssd1 vccd1 vccd1 _02667_ sky130_fd_sc_hd__a221o_1
XFILLER_0_64_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_174_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07459_ top.DUT.register\[10\]\[15\] net771 net731 top.DUT.register\[14\]\[15\] vssd1
+ vssd1 vccd1 vccd1 _02598_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout510_X net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11270__A2 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_272 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout608_X net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_376 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10470_ net1508 net248 net361 vssd1 vssd1 vccd1 vccd1 _00640_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11022__A2 net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09129_ net890 net900 vssd1 vssd1 vccd1 vccd1 _04204_ sky130_fd_sc_hd__and2_1
XANTENNA__07777__A2 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12140_ _06011_ _06021_ _06020_ _06014_ vssd1 vssd1 vccd1 vccd1 _06023_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_94_1849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08974__B2 net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08005__A _03122_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout977_X net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06985__B1 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12523__Q top.a1.halfData\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12071_ _05935_ _05937_ _05930_ vssd1 vssd1 vccd1 vccd1 _05954_ sky130_fd_sc_hd__a21o_1
XFILLER_0_4_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold580 top.DUT.register\[12\]\[17\] vssd1 vssd1 vccd1 vccd1 net1696 sky130_fd_sc_hd__dlygate4sd3_1
Xhold591 top.DUT.register\[17\]\[30\] vssd1 vssd1 vccd1 vccd1 net1707 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08726__A1 net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11022_ net32 net842 net819 net1117 vssd1 vssd1 vccd1 vccd1 _01134_ sky130_fd_sc_hd__a22o_1
XANTENNA__07563__B _02701_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_204_Left_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_125_2326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12973_ clknet_leaf_42_clk _00565_ net1058 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[14\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09687__C1 net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_197_640 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11924_ _05759_ _05760_ vssd1 vssd1 vccd1 vccd1 _05807_ sky130_fd_sc_hd__and2_2
XFILLER_0_59_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07162__B1 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07701__A2 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_196_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11855_ _05677_ _05710_ _05737_ vssd1 vssd1 vccd1 vccd1 _05738_ sky130_fd_sc_hd__or3_1
XANTENNA__06466__Y _01605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_184_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10806_ net196 net1693 net601 vssd1 vssd1 vccd1 vccd1 _00967_ sky130_fd_sc_hd__mux2_1
X_11786_ _05655_ _05656_ _05638_ vssd1 vssd1 vccd1 vccd1 _05669_ sky130_fd_sc_hd__a21oi_4
XANTENNA__09454__A2 _04487_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08961__A1_N _01960_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_200_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_171_3014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_1989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13525_ clknet_leaf_74_clk top.a1.nextHex\[3\] net1077 vssd1 vssd1 vccd1 vccd1 _01379_
+ sky130_fd_sc_hd__dfrtp_1
X_10737_ net1321 _04760_ net418 vssd1 vssd1 vccd1 vccd1 _00898_ sky130_fd_sc_hd__mux2_1
XFILLER_0_165_581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_376 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06482__X _01621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13456_ clknet_leaf_28_clk _01048_ net1011 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[29\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_180_551 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10668_ net2170 net241 net338 vssd1 vssd1 vccd1 vccd1 _00831_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12407_ clknet_leaf_107_clk top.ru.next_FetchedInstr\[19\] net975 vssd1 vssd1 vccd1
+ vccd1 top.a1.instruction\[19\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_3_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_2488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13387_ clknet_leaf_48_clk _00979_ net1059 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[27\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_10599_ net261 net2294 net348 vssd1 vssd1 vccd1 vccd1 _00764_ sky130_fd_sc_hd__mux2_1
XANTENNA__07768__A2 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput107 net107 vssd1 vssd1 vccd1 vccd1 SEL_O[2] sky130_fd_sc_hd__buf_2
XANTENNA__08965__B2 net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput118 net118 vssd1 vssd1 vccd1 vccd1 gpio_out[20] sky130_fd_sc_hd__buf_2
X_12338_ top.pad.button_control.r_counter\[14\] _06134_ net791 vssd1 vssd1 vccd1 vccd1
+ _06135_ sky130_fd_sc_hd__o21ai_1
XANTENNA__06976__B1 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12269_ top.lcd.cnt_500hz\[5\] _06091_ vssd1 vssd1 vccd1 vccd1 _06092_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_195_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10524__A1 net156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06728__B1 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_208_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_182_3176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06830_ top.DUT.register\[30\]\[19\] net582 net553 top.DUT.register\[3\]\[19\] vssd1
+ vssd1 vccd1 vccd1 _01969_ sky130_fd_sc_hd__a22o_1
XFILLER_0_207_254 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10180__A top.a1.instruction\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_208_799 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06761_ top.DUT.register\[11\]\[24\] net713 net705 top.DUT.register\[3\]\[24\] vssd1
+ vssd1 vccd1 vccd1 _01900_ sky130_fd_sc_hd__a22o_1
XFILLER_0_207_298 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08914__A1_N _01659_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08500_ _03575_ _03627_ net293 vssd1 vssd1 vccd1 vccd1 _03628_ sky130_fd_sc_hd__mux2_1
XANTENNA__07760__Y _02899_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06692_ _01809_ _01830_ vssd1 vssd1 vccd1 vccd1 _01831_ sky130_fd_sc_hd__nor2_1
X_09480_ net137 _04523_ _04533_ net901 vssd1 vssd1 vccd1 vccd1 _04534_ sky130_fd_sc_hd__o211ai_1
XANTENNA__07153__B1 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_201_3460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09693__A2 _01489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13725__RESET_B net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_wire409_X net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08431_ _02525_ net492 _03560_ net428 vssd1 vssd1 vccd1 vccd1 _03562_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__06900__B1 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11215__S net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08362_ net283 _03493_ _03494_ net280 _03492_ vssd1 vssd1 vccd1 vccd1 _03495_ sky130_fd_sc_hd__o32a_1
XFILLER_0_74_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_671 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_559 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07313_ _02445_ _02447_ _02449_ _02451_ vssd1 vssd1 vccd1 vccd1 _02452_ sky130_fd_sc_hd__or4_4
X_08293_ net317 _03428_ _03402_ vssd1 vssd1 vccd1 vccd1 _03429_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout136_A net139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07244_ _02376_ _02379_ _02381_ _02382_ vssd1 vssd1 vccd1 vccd1 _02383_ sky130_fd_sc_hd__or4_4
XFILLER_0_116_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_30_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07175_ top.DUT.register\[16\]\[10\] net543 net511 top.DUT.register\[24\]\[10\] _02313_
+ vssd1 vssd1 vccd1 vccd1 _02314_ sky130_fd_sc_hd__a221o_1
XANTENNA__10212__A0 net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1045_A net1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08956__B2 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06967__B1 net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout301 _02974_ vssd1 vssd1 vccd1 vccd1 net301 sky130_fd_sc_hd__buf_2
XANTENNA__08708__A1 net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout312 net314 vssd1 vssd1 vccd1 vccd1 net312 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08708__B2 _03168_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_167_2949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout323 net326 vssd1 vssd1 vccd1 vccd1 net323 sky130_fd_sc_hd__clkbuf_2
Xfanout334 net337 vssd1 vssd1 vccd1 vccd1 net334 sky130_fd_sc_hd__clkbuf_8
XANTENNA__06719__B1 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout672_A _01597_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout345 _04992_ vssd1 vssd1 vccd1 vccd1 net345 sky130_fd_sc_hd__clkbuf_4
Xfanout356 _04989_ vssd1 vssd1 vccd1 vccd1 net356 sky130_fd_sc_hd__buf_6
X_09816_ net1898 net185 net633 vssd1 vssd1 vccd1 vccd1 _00140_ sky130_fd_sc_hd__mux2_1
Xfanout367 net368 vssd1 vssd1 vccd1 vccd1 net367 sky130_fd_sc_hd__buf_6
Xfanout378 net379 vssd1 vssd1 vccd1 vccd1 net378 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout1000_X net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout389 net392 vssd1 vssd1 vccd1 vccd1 net389 sky130_fd_sc_hd__buf_6
XANTENNA__07392__B1 net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07931__A2 _02589_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09747_ _03663_ net403 net488 _04770_ vssd1 vssd1 vccd1 vccd1 _04771_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout460_X net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06959_ top.DUT.register\[3\]\[23\] net552 net546 top.DUT.register\[16\]\[23\] _02097_
+ vssd1 vssd1 vccd1 vccd1 _02098_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_107_2045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout558_X net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_448 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_107_2056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_190_Right_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07144__B1 net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09678_ net689 _04712_ _04713_ vssd1 vssd1 vccd1 vccd1 _04714_ sky130_fd_sc_hd__and3_4
X_08629_ _01962_ _03185_ net499 _01963_ vssd1 vssd1 vccd1 vccd1 _03751_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA_fanout725_X net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_2245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11640_ _05514_ _05515_ top.a1.dataIn\[12\] vssd1 vssd1 vccd1 vccd1 _05523_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_194_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_166_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_181_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11779__B1 top.a1.dataIn\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_194_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_166_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_3_2_0_clk_X clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11571_ _05425_ _05428_ net249 vssd1 vssd1 vccd1 vccd1 _05454_ sky130_fd_sc_hd__and3_1
XANTENNA__08644__B1 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13310_ clknet_leaf_21_clk _00902_ net1034 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[25\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07998__A2 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10522_ net1848 net164 net359 vssd1 vssd1 vccd1 vccd1 _00691_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_150_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13241_ clknet_leaf_13_clk _00833_ net955 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[23\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_10453_ net176 net2171 net367 vssd1 vssd1 vccd1 vccd1 _00624_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08947__B2 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_150_768 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10384_ net1483 net182 net374 vssd1 vssd1 vccd1 vccd1 _00559_ sky130_fd_sc_hd__mux2_1
X_13172_ clknet_leaf_57_clk _00764_ net1076 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[21\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_435 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06958__B1 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12123_ top.a1.dataIn\[2\] _06004_ vssd1 vssd1 vccd1 vccd1 _06006_ sky130_fd_sc_hd__xor2_1
X_12054_ _05928_ _05932_ _05933_ _05934_ _05927_ vssd1 vssd1 vccd1 vccd1 _05937_ sky130_fd_sc_hd__a41o_2
XANTENNA__10506__A1 net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09492__C _04543_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11005_ net1160 _05037_ net589 vssd1 vssd1 vccd1 vccd1 _01124_ sky130_fd_sc_hd__mux2_1
XANTENNA__10204__S net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07383__A0 _02502_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout890 net892 vssd1 vssd1 vccd1 vccd1 net890 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_99_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12956_ clknet_leaf_0_clk _00548_ net915 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[14\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07135__B1 net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11907_ _05758_ _05760_ _05789_ vssd1 vssd1 vccd1 vccd1 _05790_ sky130_fd_sc_hd__a21oi_1
X_12887_ clknet_leaf_129_clk _00479_ net909 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[12\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_47_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06196__Y _01427_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_47_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11838_ _05691_ _05692_ _05695_ _05720_ vssd1 vssd1 vccd1 vccd1 _05721_ sky130_fd_sc_hd__a22o_1
XFILLER_0_114_68 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_2517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10874__S net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11769_ _05606_ _05646_ _05650_ _05648_ vssd1 vssd1 vccd1 vccd1 _05652_ sky130_fd_sc_hd__nor4b_1
XFILLER_0_99_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_40_clk clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_40_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_60_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13508_ clknet_leaf_37_clk _01100_ net1052 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[31\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07989__A2 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_151_2706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10993__B2 top.a1.dataIn\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_151_2717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06661__A2 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13439_ clknet_leaf_19_clk _01031_ net1027 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[29\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_141_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12771__RESET_B net1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_184_3205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07610__A1 _02748_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08980_ _03616_ _03637_ _04054_ _03592_ vssd1 vssd1 vccd1 vccd1 _04055_ sky130_fd_sc_hd__or4b_1
XFILLER_0_121_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07931_ _02580_ _02589_ _02610_ vssd1 vssd1 vccd1 vccd1 _03070_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_149_2679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10114__S net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07862_ top.DUT.register\[20\]\[1\] net665 net717 top.DUT.register\[27\]\[1\] vssd1
+ vssd1 vccd1 vccd1 _03001_ sky130_fd_sc_hd__a22o_1
X_09601_ _04643_ _04645_ _04646_ vssd1 vssd1 vccd1 vccd1 _04647_ sky130_fd_sc_hd__o21a_1
XANTENNA__07913__A2 _02849_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06813_ top.DUT.register\[18\]\[17\] net726 net719 top.DUT.register\[19\]\[17\] vssd1
+ vssd1 vccd1 vccd1 _01952_ sky130_fd_sc_hd__a22o_1
XFILLER_0_155_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07793_ top.DUT.register\[2\]\[2\] net559 net543 top.DUT.register\[16\]\[2\] vssd1
+ vssd1 vccd1 vccd1 _02932_ sky130_fd_sc_hd__a22o_1
XANTENNA__11293__X _05183_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_162_2879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_402 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09532_ _01505_ _04581_ _04582_ _04576_ _01393_ vssd1 vssd1 vccd1 vccd1 _04583_ sky130_fd_sc_hd__a311o_1
X_06744_ top.DUT.register\[8\]\[24\] net541 net517 top.DUT.register\[7\]\[24\] vssd1
+ vssd1 vccd1 vccd1 _01883_ sky130_fd_sc_hd__a22o_1
XANTENNA__09666__A2 _02952_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06675_ top.DUT.register\[1\]\[26\] net756 net733 top.DUT.register\[14\]\[26\] vssd1
+ vssd1 vccd1 vccd1 _01814_ sky130_fd_sc_hd__a22o_1
X_09463_ _04500_ _04515_ _04516_ net811 vssd1 vssd1 vccd1 vccd1 _04518_ sky130_fd_sc_hd__a31o_1
XANTENNA__08874__B1 _03980_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13722__Q top.a1.row2\[40\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout253_A _04741_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_195_3367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08414_ _03260_ _03539_ _03543_ _03169_ _03545_ vssd1 vssd1 vccd1 vccd1 _03546_ sky130_fd_sc_hd__o221a_1
XFILLER_0_59_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_195_3378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09394_ net804 _02679_ _04335_ _04452_ vssd1 vssd1 vccd1 vccd1 _04453_ sky130_fd_sc_hd__o22a_4
XANTENNA__10784__S net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08345_ _02800_ net432 net500 _02801_ _03478_ vssd1 vssd1 vccd1 vccd1 _03479_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout420_A net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_31_clk clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_31_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout518_A _01558_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout139_X net139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08276_ net298 _02899_ vssd1 vssd1 vccd1 vccd1 _03412_ sky130_fd_sc_hd__or2_1
XFILLER_0_144_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_78_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06652__A2 net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07227_ top.DUT.register\[13\]\[10\] net774 net754 top.DUT.register\[1\]\[10\] vssd1
+ vssd1 vccd1 vccd1 _02366_ sky130_fd_sc_hd__a22o_1
XFILLER_0_131_212 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout306_X net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08929__A1 net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1048_X net1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12186__B1 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08929__B2 net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07158_ top.DUT.register\[30\]\[11\] net758 net746 top.DUT.register\[17\]\[11\] vssd1
+ vssd1 vccd1 vccd1 _02297_ sky130_fd_sc_hd__a22o_1
XFILLER_0_14_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_91_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06404__A2 net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07089_ top.DUT.register\[3\]\[16\] net552 net535 top.DUT.register\[19\]\[16\] vssd1
+ vssd1 vccd1 vccd1 _02228_ sky130_fd_sc_hd__a22o_1
XFILLER_0_100_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_98_clk clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_98_clk
+ sky130_fd_sc_hd__clkbuf_8
Xfanout131 _05690_ vssd1 vssd1 vccd1 vccd1 net131 sky130_fd_sc_hd__buf_2
XANTENNA_fanout675_X net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout142 net143 vssd1 vssd1 vccd1 vccd1 net142 sky130_fd_sc_hd__clkbuf_2
Xfanout153 _04929_ vssd1 vssd1 vccd1 vccd1 net153 sky130_fd_sc_hd__buf_1
XANTENNA__10024__S net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout164 net167 vssd1 vssd1 vccd1 vccd1 net164 sky130_fd_sc_hd__clkbuf_2
Xfanout175 _04876_ vssd1 vssd1 vccd1 vccd1 net175 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__07365__B1 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout186 net187 vssd1 vssd1 vccd1 vccd1 net186 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout197 _04788_ vssd1 vssd1 vccd1 vccd1 net197 sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_EDGE_ROW_137_Left_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout842_X net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_199_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12810_ clknet_leaf_118_clk _00402_ net955 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[9\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_13790_ clknet_leaf_68_clk _01359_ vssd1 vssd1 vccd1 vccd1 top.pad.button_control.r_counter\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__07117__B1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_232 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12741_ clknet_leaf_35_clk _00333_ net1041 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[7\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_167_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_276 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12672_ clknet_leaf_113_clk _00264_ net991 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[5\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_13814__1099 vssd1 vssd1 vccd1 vccd1 _13814__1099/HI net1099 sky130_fd_sc_hd__conb_1
XFILLER_0_65_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11623_ top.a1.dataIn\[12\] _05502_ _05504_ vssd1 vssd1 vccd1 vccd1 _05506_ sky130_fd_sc_hd__or3_1
XANTENNA__06891__A2 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_100_1948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_22_clk clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_22_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_92_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11554_ _05435_ _05436_ vssd1 vssd1 vccd1 vccd1 _05437_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_146_Left_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_42_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10505_ net1444 net233 net357 vssd1 vssd1 vccd1 vccd1 _00674_ sky130_fd_sc_hd__mux2_1
XANTENNA__12529__RESET_B net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06643__A2 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_190_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_595 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11485_ _05335_ _05357_ _05340_ vssd1 vssd1 vccd1 vccd1 _05368_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_133_2436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_2447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13224_ clknet_leaf_27_clk _00816_ net1008 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[22\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_10436_ net241 net2296 net365 vssd1 vssd1 vccd1 vccd1 _00607_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13155_ clknet_leaf_60_clk _00747_ net1088 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[20\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_209_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10367_ net1398 net252 net374 vssd1 vssd1 vccd1 vccd1 _00542_ sky130_fd_sc_hd__mux2_1
X_12106_ _05970_ _05972_ _05978_ vssd1 vssd1 vccd1 vccd1 _05989_ sky130_fd_sc_hd__and3b_1
XFILLER_0_209_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10298_ net265 net1955 net381 vssd1 vssd1 vccd1 vccd1 _00475_ sky130_fd_sc_hd__mux2_1
X_13086_ clknet_leaf_18_clk _00678_ net1027 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[18\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_89_clk clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_89_clk
+ sky130_fd_sc_hd__clkbuf_8
X_12037_ _05912_ _05919_ vssd1 vssd1 vccd1 vccd1 _05920_ sky130_fd_sc_hd__nand2b_1
XPHY_EDGE_ROW_155_Left_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11257__C top.lcd.nextState\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07356__B1 net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_68 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13388__RESET_B net1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10869__S net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_192_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07108__B1 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_198_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12939_ clknet_leaf_50_clk _00531_ net1059 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[13\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06460_ _01595_ _01598_ vssd1 vssd1 vccd1 vccd1 _01599_ sky130_fd_sc_hd__nor2_4
XFILLER_0_87_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_177_3097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09678__B _04712_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_408 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06882__A2 net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06391_ top.DUT.register\[20\]\[30\] net565 net464 top.DUT.register\[13\]\[30\] _01526_
+ vssd1 vssd1 vccd1 vccd1 _01530_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_164_Left_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_13_clk clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_13_clk
+ sky130_fd_sc_hd__clkbuf_8
X_08130_ net886 top.ru.state\[0\] net833 vssd1 vssd1 vccd1 vccd1 _03269_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_172_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_172_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_160_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06383__A top.a1.instruction\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_184 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10966__A1 top.a1.halfData\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_190_3297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08061_ _01897_ net299 vssd1 vssd1 vccd1 vccd1 _03200_ sky130_fd_sc_hd__nand2_1
XANTENNA__06634__A2 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10109__S net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07012_ top.DUT.register\[21\]\[20\] net450 net445 top.DUT.register\[1\]\[20\] _02150_
+ vssd1 vssd1 vccd1 vccd1 _02151_ sky130_fd_sc_hd__a221o_1
XANTENNA__12168__B1 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_768 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10192__X _04972_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_84 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07595__B1 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08963_ net414 net691 net1154 net874 vssd1 vssd1 vccd1 vccd1 _00069_ sky130_fd_sc_hd__a2bb2o_1
XPHY_EDGE_ROW_173_Left_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_164_2908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07914_ _02803_ _03052_ vssd1 vssd1 vccd1 vccd1 _03053_ sky130_fd_sc_hd__nand2_1
X_08894_ net435 _03999_ _04003_ net427 _04002_ vssd1 vssd1 vccd1 vccd1 _04004_ sky130_fd_sc_hd__a221o_1
XANTENNA__07347__B1 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1008_A net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07845_ _02977_ _02979_ _02981_ _02983_ vssd1 vssd1 vccd1 vccd1 _02984_ sky130_fd_sc_hd__or4_2
XANTENNA__10779__S net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout370_A net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_197_3407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout468_A net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07661__B _02798_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_196_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_104_2004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07776_ top.DUT.register\[16\]\[2\] net734 _02910_ _02911_ _02914_ vssd1 vssd1 vccd1
+ vccd1 _02915_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_88_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09515_ _04205_ _04559_ _04566_ _04051_ top.pc\[25\] vssd1 vssd1 vccd1 vccd1 _00105_
+ sky130_fd_sc_hd__o32a_1
XFILLER_0_39_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06727_ top.DUT.register\[6\]\[25\] net635 net718 top.DUT.register\[19\]\[25\] _01863_
+ vssd1 vssd1 vccd1 vccd1 _01866_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout635_A _01629_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09869__A top.pc\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09446_ _04500_ _04501_ vssd1 vssd1 vccd1 vccd1 _04502_ sky130_fd_sc_hd__and2_1
XFILLER_0_137_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_182_Left_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06658_ top.DUT.register\[3\]\[26\] net554 net549 top.DUT.register\[18\]\[26\] vssd1
+ vssd1 vccd1 vccd1 _01797_ sky130_fd_sc_hd__a22o_1
XFILLER_0_94_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_149_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_164_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06873__A2 net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09377_ net820 _02774_ vssd1 vssd1 vccd1 vccd1 _04437_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout802_A _03269_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout423_X net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06589_ top.DUT.register\[13\]\[28\] net776 net761 top.DUT.register\[30\]\[28\] vssd1
+ vssd1 vccd1 vccd1 _01728_ sky130_fd_sc_hd__a22o_1
XFILLER_0_148_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_611 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08328_ _02803_ _03052_ vssd1 vssd1 vccd1 vccd1 _03462_ sky130_fd_sc_hd__or2_1
XFILLER_0_151_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08259_ _03393_ _03394_ net312 vssd1 vssd1 vccd1 vccd1 _03395_ sky130_fd_sc_hd__mux2_1
XANTENNA__10019__S net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_519 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11270_ net1157 net814 _05161_ net1003 vssd1 vssd1 vccd1 vccd1 _01265_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_115_2166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_576 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_2177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08378__A2 net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10221_ net175 net2134 net395 vssd1 vssd1 vccd1 vccd1 _00401_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10152_ net2269 net241 net602 vssd1 vssd1 vccd1 vccd1 _00351_ sky130_fd_sc_hd__mux2_1
XANTENNA__09109__A top.pc\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07050__A2 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10083_ net2237 net260 net613 vssd1 vssd1 vccd1 vccd1 _00284_ sky130_fd_sc_hd__mux2_1
Xhold9 top.a1.dataInTemp\[5\] vssd1 vssd1 vccd1 vccd1 net1125 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13481__RESET_B net1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10689__S net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input29_A DAT_I[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13773_ clknet_leaf_100_clk _01344_ vssd1 vssd1 vccd1 vccd1 top.lcd.cnt_500hz\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10985_ net843 _05021_ _05022_ net849 top.a1.dataIn\[5\] vssd1 vssd1 vccd1 vccd1
+ _05023_ sky130_fd_sc_hd__a32o_1
XFILLER_0_85_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12724_ clknet_leaf_79_clk _00316_ net1072 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[7\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_44_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07510__B1 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_194_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06864__A2 net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_182_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12655_ clknet_leaf_22_clk _00247_ net1023 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[4\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06474__Y _01613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11606_ _05485_ _05486_ _05480_ vssd1 vssd1 vccd1 vccd1 _05489_ sky130_fd_sc_hd__a21o_1
XFILLER_0_53_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_791 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12586_ clknet_leaf_118_clk _00178_ net953 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[2\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_142_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_627 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12363__RESET_B net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06616__A2 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11537_ _05361_ _05416_ vssd1 vssd1 vccd1 vccd1 _05420_ sky130_fd_sc_hd__xor2_1
XFILLER_0_151_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold409 top.DUT.register\[20\]\[1\] vssd1 vssd1 vccd1 vccd1 net1525 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06490__X _01629_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06931__A _02069_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11468_ _05322_ _05350_ vssd1 vssd1 vccd1 vccd1 _05351_ sky130_fd_sc_hd__xnor2_1
Xmax_cap128 _05817_ vssd1 vssd1 vccd1 vccd1 net128 sky130_fd_sc_hd__clkbuf_2
X_13207_ clknet_leaf_3_clk _00799_ net919 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[22\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_96_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10419_ net1383 net181 net369 vssd1 vssd1 vccd1 vccd1 _00591_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_790 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11399_ _05279_ _05281_ vssd1 vssd1 vccd1 vccd1 _05282_ sky130_fd_sc_hd__and2b_1
XANTENNA__07577__B1 net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_596 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07041__A2 net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13138_ clknet_leaf_23_clk _00730_ net1021 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[20\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_55_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13069_ clknet_leaf_42_clk _00661_ net1058 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[17\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_2_clk clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_2_clk
+ sky130_fd_sc_hd__clkbuf_8
Xhold1109 top.DUT.register\[21\]\[0\] vssd1 vssd1 vccd1 vccd1 net2225 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07329__B1 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_146_2638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09306__X _04370_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_119_Right_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10599__S net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07630_ top.DUT.register\[10\]\[5\] net519 net439 top.DUT.register\[5\]\[5\] _02768_
+ vssd1 vssd1 vccd1 vccd1 _02769_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_179_3126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_179_3137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_178_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08829__B1 net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07561_ _02695_ _02697_ _02699_ vssd1 vssd1 vccd1 vccd1 _02700_ sky130_fd_sc_hd__or3_1
XFILLER_0_88_574 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09300_ top.pc\[13\] _04352_ vssd1 vssd1 vccd1 vccd1 _04364_ sky130_fd_sc_hd__nor2_1
X_06512_ top.DUT.register\[20\]\[30\] net665 net721 top.DUT.register\[19\]\[30\] _01650_
+ vssd1 vssd1 vccd1 vccd1 _01651_ sky130_fd_sc_hd__a221o_1
XFILLER_0_158_451 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07492_ top.DUT.register\[13\]\[14\] net465 net524 top.DUT.register\[11\]\[14\] _02630_
+ vssd1 vssd1 vccd1 vccd1 _02631_ sky130_fd_sc_hd__a221o_1
XFILLER_0_119_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_192_3326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07501__B1 net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09231_ _02502_ top.pc\[9\] vssd1 vssd1 vccd1 vccd1 _04299_ sky130_fd_sc_hd__and2b_1
XANTENNA__06855__A2 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06443_ top.a1.instruction\[31\] net789 net794 top.a1.instruction\[23\] vssd1 vssd1
+ vccd1 vccd1 _01582_ sky130_fd_sc_hd__a22o_1
XFILLER_0_185_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06374_ top.a1.instruction\[17\] top.a1.instruction\[18\] net683 _01512_ vssd1 vssd1
+ vccd1 vccd1 _01513_ sky130_fd_sc_hd__and4_4
X_09162_ net903 top.pc\[4\] net890 vssd1 vssd1 vccd1 vccd1 _04235_ sky130_fd_sc_hd__o21a_1
XFILLER_0_145_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_290 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08113_ _02544_ net331 vssd1 vssd1 vccd1 vccd1 _03252_ sky130_fd_sc_hd__nand2_1
XFILLER_0_160_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06607__A2 net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_211_3610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09093_ top.a1.instruction\[14\] _01479_ _03150_ _04146_ vssd1 vssd1 vccd1 vccd1
+ _04168_ sky130_fd_sc_hd__a211o_1
XFILLER_0_43_154 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_211_3621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_474 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_211_3632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08044_ _03182_ vssd1 vssd1 vccd1 vccd1 _03183_ sky130_fd_sc_hd__inv_2
XANTENNA__09793__B1_N _04811_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07280__A2 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_170_2989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold910 top.DUT.register\[29\]\[20\] vssd1 vssd1 vccd1 vccd1 net2026 sky130_fd_sc_hd__dlygate4sd3_1
Xhold921 top.DUT.register\[26\]\[22\] vssd1 vssd1 vccd1 vccd1 net2037 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold932 top.DUT.register\[11\]\[7\] vssd1 vssd1 vccd1 vccd1 net2048 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold943 top.DUT.register\[2\]\[0\] vssd1 vssd1 vccd1 vccd1 net2059 sky130_fd_sc_hd__dlygate4sd3_1
Xhold954 top.DUT.register\[14\]\[23\] vssd1 vssd1 vccd1 vccd1 net2070 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07568__B1 net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold965 top.DUT.register\[25\]\[15\] vssd1 vssd1 vccd1 vccd1 net2081 sky130_fd_sc_hd__dlygate4sd3_1
Xhold976 top.DUT.register\[16\]\[20\] vssd1 vssd1 vccd1 vccd1 net2092 sky130_fd_sc_hd__dlygate4sd3_1
Xhold987 top.DUT.register\[7\]\[6\] vssd1 vssd1 vccd1 vccd1 net2103 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07032__A2 net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold998 top.DUT.register\[19\]\[4\] vssd1 vssd1 vccd1 vccd1 net2114 sky130_fd_sc_hd__dlygate4sd3_1
X_09995_ net188 net2006 net626 vssd1 vssd1 vccd1 vccd1 _00200_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout585_A _01513_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08946_ net1247 net873 _02922_ net693 vssd1 vssd1 vccd1 vccd1 _00052_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_110_2096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11116__A1 net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_209_3583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08877_ _03969_ _03987_ vssd1 vssd1 vccd1 vccd1 _03988_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout373_X net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout752_A _01621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10302__S net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07828_ top.DUT.register\[20\]\[0\] net663 _02965_ _02966_ vssd1 vssd1 vccd1 vccd1
+ _02967_ sky130_fd_sc_hd__a211o_1
XFILLER_0_193_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_86_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12815__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_190_Left_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout540_X net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07759_ _02891_ _02893_ _02895_ _02897_ vssd1 vssd1 vccd1 vccd1 _02898_ sky130_fd_sc_hd__or4_4
XFILLER_0_67_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout638_X net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07099__A2 net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09599__A net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_183_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10770_ net1761 net227 net482 vssd1 vssd1 vccd1 vccd1 _00931_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12803__RESET_B net1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09429_ _04482_ _04485_ vssd1 vssd1 vccd1 vccd1 _04486_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_137_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06846__A2 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09111__B _02999_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12440_ clknet_leaf_75_clk _00036_ net1079 vssd1 vssd1 vccd1 vccd1 top.ramaddr\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_191_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_117_2206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_644 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08008__A top.a1.instruction\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12526__Q top.a1.halfData\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08599__A2 _03708_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12371_ clknet_leaf_105_clk top.ru.next_FetchedData\[15\] net972 vssd1 vssd1 vccd1
+ vccd1 top.a1.dataIn\[15\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_50_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11322_ top.a1.dataIn\[31\] top.a1.dataIn\[30\] vssd1 vssd1 vccd1 vccd1 _05205_ sky130_fd_sc_hd__and2_1
XFILLER_0_160_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07271__A2 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11253_ net880 top.lcd.nextState\[0\] _05119_ vssd1 vssd1 vccd1 vccd1 _05146_ sky130_fd_sc_hd__and3_1
XANTENNA__07559__B1 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10204_ net246 net1890 net393 vssd1 vssd1 vccd1 vccd1 _00384_ sky130_fd_sc_hd__mux2_1
XANTENNA__07023__A2 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11184_ _05028_ _05038_ net473 net587 net1158 vssd1 vssd1 vccd1 vccd1 _01241_ sky130_fd_sc_hd__a32o_1
XANTENNA__08771__A2 net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10135_ net181 net1774 net608 vssd1 vssd1 vccd1 vccd1 _00335_ sky130_fd_sc_hd__mux2_1
XANTENNA__08678__A net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10066_ net2147 net186 net618 vssd1 vssd1 vccd1 vccd1 _00268_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_128_2368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08030__X _03169_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09720__A1 _03548_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10212__S net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_50_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_187_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06198__A net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07731__B1 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_202_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13825_ net1109 vssd1 vssd1 vccd1 vccd1 gpio_out[24] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_141_2557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_546 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_141_2568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13756_ clknet_leaf_99_clk _01327_ vssd1 vssd1 vccd1 vccd1 top.lcd.cnt_20ms\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__06485__X _01624_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10968_ top.a1.dataIn\[1\] net850 _05008_ _05009_ vssd1 vssd1 vccd1 vccd1 _05010_
+ sky130_fd_sc_hd__a22o_1
X_12707_ clknet_leaf_60_clk _00299_ net1088 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[6\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06837__A2 net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_174_3056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13687_ clknet_leaf_74_clk _01263_ net1079 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[13\]
+ sky130_fd_sc_hd__dfstp_1
X_10899_ net2293 net219 net478 vssd1 vssd1 vccd1 vccd1 _01060_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_182_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12638_ clknet_leaf_18_clk _00230_ net1031 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[4\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_127_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_143 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10882__S net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12569_ clknet_leaf_14_clk _00161_ net959 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[2\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07798__B1 net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold206 top.DUT.register\[14\]\[15\] vssd1 vssd1 vccd1 vccd1 net1322 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07262__A2 net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold217 top.DUT.register\[4\]\[27\] vssd1 vssd1 vccd1 vccd1 net1333 sky130_fd_sc_hd__dlygate4sd3_1
Xhold228 top.DUT.register\[15\]\[26\] vssd1 vssd1 vccd1 vccd1 net1344 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12177__A2_N _05083_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold239 top.DUT.register\[31\]\[23\] vssd1 vssd1 vccd1 vccd1 net1355 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07014__A2 net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout708 _01640_ vssd1 vssd1 vccd1 vccd1 net708 sky130_fd_sc_hd__clkbuf_8
Xfanout719 _01635_ vssd1 vssd1 vccd1 vccd1 net719 sky130_fd_sc_hd__clkbuf_4
X_08800_ net497 _03913_ vssd1 vssd1 vccd1 vccd1 _03914_ sky130_fd_sc_hd__nor2_1
XANTENNA__13332__RESET_B net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09780_ _04797_ _04798_ vssd1 vssd1 vccd1 vccd1 _04800_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_7_Right_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06992_ _02122_ _02130_ vssd1 vssd1 vccd1 vccd1 _02131_ sky130_fd_sc_hd__nor2_4
XANTENNA__07970__B1 net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08731_ net883 top.pc\[21\] net694 _03848_ vssd1 vssd1 vccd1 vccd1 _03849_ sky130_fd_sc_hd__a22o_1
XFILLER_0_56_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_147_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08662_ _01964_ _03762_ _03077_ vssd1 vssd1 vccd1 vccd1 _03783_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10122__S net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08100__B net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07722__B1 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07613_ _02724_ _02749_ vssd1 vssd1 vccd1 vccd1 _02752_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_1_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08593_ _03542_ _03716_ net297 vssd1 vssd1 vccd1 vccd1 _03717_ sky130_fd_sc_hd__mux2_1
XFILLER_0_178_568 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12988__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07544_ top.DUT.register\[1\]\[7\] net754 net746 top.DUT.register\[17\]\[7\] vssd1
+ vssd1 vccd1 vccd1 _02683_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_159_2829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_159_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_193_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06828__A2 net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11282__B1 _05150_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_81_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07475_ _02612_ _02613_ vssd1 vssd1 vccd1 vccd1 _02614_ sky130_fd_sc_hd__nor2_2
XFILLER_0_48_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout333_A _03121_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1075_A net1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09214_ _04271_ _04282_ _04283_ vssd1 vssd1 vccd1 vccd1 _00087_ sky130_fd_sc_hd__a21oi_1
X_06426_ net683 _01516_ _01527_ vssd1 vssd1 vccd1 vccd1 _01565_ sky130_fd_sc_hd__and3_2
XFILLER_0_91_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09145_ _04195_ _04197_ _04217_ vssd1 vssd1 vccd1 vccd1 _04219_ sky130_fd_sc_hd__a21o_1
X_06357_ top.pad.button_control.r_counter\[1\] top.pad.button_control.r_counter\[4\]
+ top.pad.button_control.r_counter\[3\] _01490_ vssd1 vssd1 vccd1 vccd1 _01497_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_20_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10792__S net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout500_A net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07789__B1 net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_479 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09076_ _01389_ net822 vssd1 vssd1 vccd1 vccd1 _04151_ sky130_fd_sc_hd__nand2_4
XFILLER_0_71_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07253__A2 net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06288_ _01448_ vssd1 vssd1 vccd1 vccd1 _01334_ sky130_fd_sc_hd__inv_2
X_08027_ _03102_ _03145_ _03161_ _03165_ vssd1 vssd1 vccd1 vccd1 _03166_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_96_1880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_96_1891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold740 top.DUT.register\[20\]\[14\] vssd1 vssd1 vccd1 vccd1 net1856 sky130_fd_sc_hd__dlygate4sd3_1
Xhold751 top.DUT.register\[28\]\[26\] vssd1 vssd1 vccd1 vccd1 net1867 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold762 top.DUT.register\[29\]\[17\] vssd1 vssd1 vccd1 vccd1 net1878 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07005__A2 net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold773 top.DUT.register\[12\]\[20\] vssd1 vssd1 vccd1 vccd1 net1889 sky130_fd_sc_hd__dlygate4sd3_1
Xhold784 top.DUT.register\[4\]\[5\] vssd1 vssd1 vccd1 vccd1 net1900 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout490_X net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold795 top.DUT.register\[16\]\[10\] vssd1 vssd1 vccd1 vccd1 net1911 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout967_A net1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13073__RESET_B net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout588_X net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09978_ net690 _04712_ _04949_ vssd1 vssd1 vccd1 vccd1 _04950_ sky130_fd_sc_hd__nand3_1
X_08929_ net324 _03717_ _03877_ net279 vssd1 vssd1 vccd1 vccd1 _04037_ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout755_X net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10032__S net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11940_ _05822_ vssd1 vssd1 vccd1 vccd1 _05823_ sky130_fd_sc_hd__inv_2
XFILLER_0_207_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08910__C1 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout922_X net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11871_ top.a1.dataIn\[5\] _05751_ vssd1 vssd1 vccd1 vccd1 _05754_ sky130_fd_sc_hd__nand2_1
XFILLER_0_211_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13610_ clknet_leaf_89_clk _01197_ net1003 vssd1 vssd1 vccd1 vccd1 net67 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_196_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10822_ net150 net1855 net600 vssd1 vssd1 vccd1 vccd1 _00983_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_123_2287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_123_2298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13541_ clknet_leaf_104_clk _01128_ net973 vssd1 vssd1 vccd1 vccd1 top.ramload\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_149_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10753_ net2261 net170 net421 vssd1 vssd1 vccd1 vccd1 _00914_ sky130_fd_sc_hd__mux2_1
XANTENNA__06819__A2 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13472_ clknet_leaf_115_clk _01064_ net964 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[30\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_192_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_180_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_165_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13143__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10684_ net1340 net183 net338 vssd1 vssd1 vccd1 vccd1 _00847_ sky130_fd_sc_hd__mux2_1
XANTENNA__07492__A2 net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12423_ clknet_leaf_75_clk _00019_ net1077 vssd1 vssd1 vccd1 vccd1 top.ramaddr\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_63_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_766 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12354_ clknet_leaf_111_clk net858 net989 vssd1 vssd1 vccd1 vccd1 top.i_ready sky130_fd_sc_hd__dfrtp_1
XFILLER_0_121_800 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11305_ _05190_ _05192_ _05181_ vssd1 vssd1 vccd1 vccd1 _05193_ sky130_fd_sc_hd__or3b_1
XANTENNA__13293__CLK clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10207__S net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12285_ _06101_ vssd1 vssd1 vccd1 vccd1 _06102_ sky130_fd_sc_hd__inv_2
X_11236_ top.lcd.nextState\[3\] net878 _05128_ vssd1 vssd1 vccd1 vccd1 _05129_ sky130_fd_sc_hd__nand3_1
XFILLER_0_120_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11249__D _05118_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08744__A2 _03534_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11167_ net851 net844 _05002_ _05092_ vssd1 vssd1 vccd1 vccd1 _05093_ sky130_fd_sc_hd__or4_1
X_10118_ net254 net2060 net608 vssd1 vssd1 vccd1 vccd1 _00318_ sky130_fd_sc_hd__mux2_1
X_11098_ net905 net1631 _01428_ _05054_ vssd1 vssd1 vccd1 vccd1 _01200_ sky130_fd_sc_hd__a31o_1
X_10049_ net1850 net265 net615 vssd1 vssd1 vccd1 vccd1 _00251_ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07704__B1 net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_203_631 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10877__S net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_202_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13808_ net72 vssd1 vssd1 vccd1 vccd1 net105 sky130_fd_sc_hd__clkbuf_1
X_13739_ clknet_leaf_96_clk _01310_ vssd1 vssd1 vccd1 vccd1 top.a1.dataInTemp\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10178__A top.a1.instruction\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06375__B top.a1.instruction\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_190_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_251 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07260_ _02392_ _02394_ _02396_ _02398_ vssd1 vssd1 vccd1 vccd1 _02399_ sky130_fd_sc_hd__or4_4
XANTENNA__07483__A2 net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06211_ net1274 net859 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedInstr\[5\] sky130_fd_sc_hd__and2_1
XANTENNA__06691__B1 net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07191_ top.a1.instruction\[28\] net789 net793 top.a1.instruction\[20\] vssd1 vssd1
+ vccd1 vccd1 _02330_ sky130_fd_sc_hd__a22oi_4
XTAP_TAPCELL_ROW_154_2759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_171_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06142_ net888 vssd1 vssd1 vccd1 vccd1 _01385_ sky130_fd_sc_hd__inv_2
XFILLER_0_81_591 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07235__A2 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10184__Y _04964_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_187_3247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10117__S net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_187_3258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09901_ _04907_ _04908_ vssd1 vssd1 vccd1 vccd1 _04909_ sky130_fd_sc_hd__and2_1
XFILLER_0_111_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_98_clk_A clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout505 net506 vssd1 vssd1 vccd1 vccd1 net505 sky130_fd_sc_hd__buf_4
XFILLER_0_111_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08529__A1_N net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout516 _01558_ vssd1 vssd1 vccd1 vccd1 net516 sky130_fd_sc_hd__clkbuf_4
Xfanout527 net530 vssd1 vssd1 vccd1 vccd1 net527 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_6_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09832_ _04499_ net487 net401 top.a1.dataIn\[21\] net397 vssd1 vssd1 vccd1 vccd1
+ _04847_ sky130_fd_sc_hd__a221o_1
XANTENNA__09932__A1 _04027_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_171_Right_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_169_2980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout538 _01541_ vssd1 vssd1 vccd1 vccd1 net538 sky130_fd_sc_hd__buf_4
Xfanout549 net550 vssd1 vssd1 vccd1 vccd1 net549 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_206_3531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09207__A _02678_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_206_3542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09763_ _04784_ _04783_ vssd1 vssd1 vccd1 vccd1 _04785_ sky130_fd_sc_hd__and2b_1
XANTENNA__13725__Q top.a1.row2\[43\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06975_ top.DUT.register\[20\]\[23\] net665 net731 top.DUT.register\[14\]\[23\] _02113_
+ vssd1 vssd1 vccd1 vccd1 _02114_ sky130_fd_sc_hd__a221o_1
XANTENNA__13016__CLK clknet_leaf_128_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_21_clk_A clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08714_ _02092_ _03831_ vssd1 vssd1 vccd1 vccd1 _03832_ sky130_fd_sc_hd__xnor2_1
X_09694_ top.pc\[2\] net799 net407 _04727_ vssd1 vssd1 vccd1 vccd1 _04728_ sky130_fd_sc_hd__a211o_1
XANTENNA__11098__A3 _01428_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08645_ net1708 net833 net803 _03766_ vssd1 vssd1 vccd1 vccd1 _00035_ sky130_fd_sc_hd__a22o_1
XFILLER_0_96_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10787__S net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout450_A _01562_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout548_A net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08257__S net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08576_ _02657_ _03700_ vssd1 vssd1 vccd1 vccd1 _03701_ sky130_fd_sc_hd__nor2_1
XANTENNA_clkbuf_leaf_36_clk_A clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07527_ top.DUT.register\[11\]\[7\] net523 net503 top.DUT.register\[27\]\[7\] vssd1
+ vssd1 vccd1 vccd1 _02666_ sky130_fd_sc_hd__a22o_1
XFILLER_0_76_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_193_357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout715_A _01637_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout336_X net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09877__A top.pc\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07458_ top.DUT.register\[7\]\[15\] net662 net711 top.DUT.register\[11\]\[15\] _02596_
+ vssd1 vssd1 vccd1 vccd1 _02597_ sky130_fd_sc_hd__a221o_1
XFILLER_0_147_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06409_ top.a1.instruction\[19\] _01509_ _01546_ vssd1 vssd1 vccd1 vccd1 _01548_
+ sky130_fd_sc_hd__and3_4
XTAP_TAPCELL_ROW_98_1920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout503_X net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07389_ top.DUT.register\[6\]\[9\] net567 net503 top.DUT.register\[27\]\[9\] vssd1
+ vssd1 vccd1 vccd1 _02528_ sky130_fd_sc_hd__a22o_1
XFILLER_0_91_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09128_ top.pc\[2\] _04183_ _04202_ vssd1 vssd1 vccd1 vccd1 _04203_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_32_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09059_ _03599_ _03817_ _04130_ _04133_ vssd1 vssd1 vccd1 vccd1 _04134_ sky130_fd_sc_hd__or4_1
XFILLER_0_32_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10027__S net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08005__B _03142_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09816__S net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12070_ _05943_ _05948_ _05946_ vssd1 vssd1 vccd1 vccd1 _05953_ sky130_fd_sc_hd__or3b_1
Xhold570 top.DUT.register\[12\]\[19\] vssd1 vssd1 vccd1 vccd1 net1686 sky130_fd_sc_hd__dlygate4sd3_1
Xhold581 top.DUT.register\[9\]\[18\] vssd1 vssd1 vccd1 vccd1 net1697 sky130_fd_sc_hd__dlygate4sd3_1
Xhold592 top.ramaddr\[17\] vssd1 vssd1 vccd1 vccd1 net1708 sky130_fd_sc_hd__dlygate4sd3_1
X_11021_ net31 net838 net816 net2257 vssd1 vssd1 vccd1 vccd1 _01133_ sky130_fd_sc_hd__o22a_1
XANTENNA__09384__C1 net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_109_clk_A clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09117__A _03000_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08021__A _01501_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_125_2316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12972_ clknet_leaf_47_clk _00564_ net1069 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[14\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input11_A DAT_I[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11923_ _05783_ _05791_ vssd1 vssd1 vccd1 vccd1 _05806_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_87_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10697__S net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11854_ _05706_ _05736_ vssd1 vssd1 vccd1 vccd1 _05737_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_129_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_157_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10805_ net209 net1884 net601 vssd1 vssd1 vccd1 vccd1 _00966_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_363 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11785_ _05665_ _05666_ _05661_ vssd1 vssd1 vccd1 vccd1 _05668_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_171_3004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13524_ clknet_leaf_74_clk top.a1.nextHex\[2\] net1077 vssd1 vssd1 vccd1 vccd1 _01378_
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_171_3015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10736_ net1563 net235 net421 vssd1 vssd1 vccd1 vccd1 _00897_ sky130_fd_sc_hd__mux2_1
XANTENNA__07465__A2 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06673__B1 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13455_ clknet_leaf_21_clk _01047_ net1022 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[29\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_10667_ net1843 net253 net338 vssd1 vssd1 vccd1 vccd1 _00830_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_388 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_563 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12406_ clknet_leaf_105_clk top.ru.next_FetchedInstr\[18\] net971 vssd1 vssd1 vccd1
+ vccd1 top.a1.instruction\[18\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__08414__A1 _03260_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_2489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08414__B2 _03169_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13386_ clknet_leaf_117_clk _00978_ net957 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[27\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09611__B1 _04164_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10598_ net265 net1879 net346 vssd1 vssd1 vccd1 vccd1 _00763_ sky130_fd_sc_hd__mux2_1
XFILLER_0_112_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12337_ _06134_ net791 _06133_ vssd1 vssd1 vccd1 vccd1 _01365_ sky130_fd_sc_hd__and3b_1
XFILLER_0_11_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput108 net108 vssd1 vssd1 vccd1 vccd1 SEL_O[3] sky130_fd_sc_hd__buf_2
Xoutput119 net119 vssd1 vssd1 vccd1 vccd1 gpio_out[21] sky130_fd_sc_hd__buf_2
XFILLER_0_11_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12268_ net686 _06090_ _06091_ vssd1 vssd1 vccd1 vccd1 _01339_ sky130_fd_sc_hd__and3_1
X_11219_ _05115_ net1212 net471 vssd1 vssd1 vccd1 vccd1 _01260_ sky130_fd_sc_hd__mux2_1
X_12199_ net1132 _06019_ net688 vssd1 vssd1 vccd1 vccd1 _01306_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput90 net90 vssd1 vssd1 vccd1 vccd1 DAT_O[25] sky130_fd_sc_hd__clkbuf_4
XANTENNA__07246__S net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_182_3177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_266 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06760_ top.DUT.register\[13\]\[24\] net776 net745 top.DUT.register\[2\]\[24\] vssd1
+ vssd1 vccd1 vccd1 _01899_ sky130_fd_sc_hd__a22o_1
X_06691_ net807 _01829_ net437 vssd1 vssd1 vccd1 vccd1 _01830_ sky130_fd_sc_hd__o21a_1
XFILLER_0_203_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_201_3461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08430_ _03537_ _03559_ _03558_ vssd1 vssd1 vccd1 vccd1 _03561_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_65_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10400__S net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08361_ net311 _03356_ vssd1 vssd1 vccd1 vccd1 _03494_ sky130_fd_sc_hd__nor2_1
XFILLER_0_86_683 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07312_ top.DUT.register\[13\]\[12\] net463 net527 top.DUT.register\[26\]\[12\] _02450_
+ vssd1 vssd1 vccd1 vccd1 _02451_ sky130_fd_sc_hd__a221o_1
XANTENNA__09697__A net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08292_ net316 _03427_ _03406_ vssd1 vssd1 vccd1 vccd1 _03428_ sky130_fd_sc_hd__a21o_1
XANTENNA__07456__A2 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_190_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06664__B1 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07243_ top.DUT.register\[4\]\[10\] net667 net726 top.DUT.register\[18\]\[10\] _02368_
+ vssd1 vssd1 vccd1 vccd1 _02382_ sky130_fd_sc_hd__a221o_1
XFILLER_0_128_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_144_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07174_ top.DUT.register\[28\]\[10\] net555 net503 top.DUT.register\[27\]\[10\] vssd1
+ vssd1 vccd1 vccd1 _02313_ sky130_fd_sc_hd__a22o_1
XFILLER_0_103_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08106__A _02453_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1038_A net1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout302 net303 vssd1 vssd1 vccd1 vccd1 net302 sky130_fd_sc_hd__buf_2
XANTENNA_clkbuf_4_7__f_clk_X clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout313 net314 vssd1 vssd1 vccd1 vccd1 net313 sky130_fd_sc_hd__buf_2
Xfanout324 net326 vssd1 vssd1 vccd1 vccd1 net324 sky130_fd_sc_hd__clkbuf_4
Xfanout335 net337 vssd1 vssd1 vccd1 vccd1 net335 sky130_fd_sc_hd__buf_6
Xfanout346 _04991_ vssd1 vssd1 vccd1 vccd1 net346 sky130_fd_sc_hd__clkbuf_8
Xfanout357 net360 vssd1 vssd1 vccd1 vccd1 net357 sky130_fd_sc_hd__buf_6
XANTENNA_input3_A DAT_I[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09815_ _03807_ net405 net489 _04831_ vssd1 vssd1 vccd1 vccd1 _04832_ sky130_fd_sc_hd__o211a_2
Xfanout368 _04985_ vssd1 vssd1 vccd1 vccd1 net368 sky130_fd_sc_hd__buf_4
Xfanout379 net380 vssd1 vssd1 vccd1 vccd1 net379 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout665_A _01605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09746_ top.a1.dataIn\[12\] _04752_ _04754_ _04769_ vssd1 vssd1 vccd1 vccd1 _04770_
+ sky130_fd_sc_hd__a211o_1
X_06958_ top.DUT.register\[19\]\[23\] net536 net508 top.DUT.register\[4\]\[23\] vssd1
+ vssd1 vccd1 vccd1 _02097_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_107_2046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_2057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13832__1116 vssd1 vssd1 vccd1 vccd1 _13832__1116/HI net1116 sky130_fd_sc_hd__conb_1
XFILLER_0_69_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_179_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09677_ top.a1.instruction\[8\] net786 top.a1.instruction\[7\] vssd1 vssd1 vccd1
+ vccd1 _04713_ sky130_fd_sc_hd__and3b_2
X_06889_ top.DUT.register\[22\]\[18\] net649 net732 top.DUT.register\[14\]\[18\] vssd1
+ vssd1 vccd1 vccd1 _02028_ sky130_fd_sc_hd__a22o_1
XFILLER_0_68_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout832_A _01499_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout453_X net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08628_ net317 _03349_ vssd1 vssd1 vccd1 vccd1 _03750_ sky130_fd_sc_hd__nor2_1
XANTENNA__10310__S net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08892__A1 net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07695__A2 net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_2246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11228__B1 _01442_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout620_X net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08559_ _02434_ _03665_ _03063_ vssd1 vssd1 vccd1 vccd1 _03684_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_37_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_59_Left_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout718_X net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_240 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11570_ _05447_ _05452_ vssd1 vssd1 vccd1 vccd1 _05453_ sky130_fd_sc_hd__nor2_1
XANTENNA__07447__A2 net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08644__A1 net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08644__B2 _03765_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06655__B1 net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10521_ net2016 net171 net360 vssd1 vssd1 vccd1 vccd1 _00690_ sky130_fd_sc_hd__mux2_1
X_13240_ clknet_leaf_128_clk _00832_ net913 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[23\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_134_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10452_ net182 net1660 net368 vssd1 vssd1 vccd1 vccd1 _00623_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13171_ clknet_leaf_120_clk _00763_ net933 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[21\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_10383_ net2032 net194 net376 vssd1 vssd1 vccd1 vccd1 _00558_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_594 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12122_ _06004_ vssd1 vssd1 vccd1 vccd1 _06005_ sky130_fd_sc_hd__inv_2
XFILLER_0_103_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_68_Left_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12053_ _05932_ _05935_ vssd1 vssd1 vccd1 vccd1 _05936_ sky130_fd_sc_hd__nand2_1
XFILLER_0_102_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11004_ top.a1.dataIn\[10\] net849 net843 _05036_ vssd1 vssd1 vccd1 vccd1 _05037_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12388__RESET_B net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13331__CLK clknet_leaf_120_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07383__A1 _02521_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout880 net882 vssd1 vssd1 vccd1 vccd1 net880 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07861__Y _03000_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout891 net892 vssd1 vssd1 vccd1 vccd1 net891 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08686__A net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_3_6_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_3_6_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_205_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_189_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12955_ clknet_leaf_120_clk _00547_ net929 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[14\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_11906_ _05758_ _05784_ _05766_ vssd1 vssd1 vccd1 vccd1 _05789_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10220__S net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12886_ clknet_leaf_12_clk _00478_ net942 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[12\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07686__A2 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_655 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06894__B1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11837_ _05698_ _05703_ net130 _05718_ vssd1 vssd1 vccd1 vccd1 _05720_ sky130_fd_sc_hd__a22oi_4
XTAP_TAPCELL_ROW_138_2518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07438__A2 net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11768_ _05606_ _05650_ _05648_ vssd1 vssd1 vccd1 vccd1 _05651_ sky130_fd_sc_hd__or3b_1
XFILLER_0_138_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_60_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13507_ clknet_leaf_57_clk _01099_ net1076 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[31\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10719_ net1426 net176 net337 vssd1 vssd1 vccd1 vccd1 _00880_ sky130_fd_sc_hd__mux2_1
X_11699_ _05553_ _05581_ vssd1 vssd1 vccd1 vccd1 _05582_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_151_2707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13105__RESET_B net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_151_2718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13438_ clknet_leaf_52_clk _01030_ net1037 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[29\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_153_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09596__C1 net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10890__S net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13369_ clknet_leaf_12_clk _00961_ net943 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[27\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_184_3206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07071__B1 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09348__C1 net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07930_ _02434_ _03065_ _03068_ _02478_ _03063_ vssd1 vssd1 vccd1 vccd1 _03069_ sky130_fd_sc_hd__o221a_1
XANTENNA__10191__A top.a1.instruction\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07861_ _02999_ vssd1 vssd1 vccd1 vccd1 _03000_ sky130_fd_sc_hd__inv_2
X_09600_ _04643_ _04645_ net812 vssd1 vssd1 vccd1 vccd1 _04646_ sky130_fd_sc_hd__a21oi_1
X_06812_ top.DUT.register\[23\]\[17\] net672 net777 top.DUT.register\[13\]\[17\] vssd1
+ vssd1 vccd1 vccd1 _01951_ sky130_fd_sc_hd__a22o_1
X_07792_ top.DUT.register\[1\]\[2\] net443 net507 top.DUT.register\[4\]\[2\] _02930_
+ vssd1 vssd1 vccd1 vccd1 _02931_ sky130_fd_sc_hd__a221o_1
XFILLER_0_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_162_2869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09531_ _04561_ _04564_ _04580_ vssd1 vssd1 vccd1 vccd1 _04582_ sky130_fd_sc_hd__a21o_1
X_06743_ top.DUT.register\[9\]\[24\] net468 net458 top.DUT.register\[25\]\[24\] _01881_
+ vssd1 vssd1 vccd1 vccd1 _01882_ sky130_fd_sc_hd__a221o_1
XFILLER_0_78_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_211_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10130__S net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09462_ _04500_ _04516_ _04515_ vssd1 vssd1 vccd1 vccd1 _04517_ sky130_fd_sc_hd__a21oi_1
X_06674_ top.DUT.register\[10\]\[26\] net773 net705 top.DUT.register\[3\]\[26\] vssd1
+ vssd1 vccd1 vccd1 _01813_ sky130_fd_sc_hd__a22o_1
XANTENNA__07677__A2 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08874__B2 _03259_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08413_ net494 _03519_ _03544_ vssd1 vssd1 vccd1 vccd1 _03545_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_195_3368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06885__B1 net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_655 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09393_ net820 _02726_ vssd1 vssd1 vccd1 vccd1 _04452_ sky130_fd_sc_hd__nor2_1
XFILLER_0_93_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_35_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout246_A _04749_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_171_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08344_ _02803_ net492 vssd1 vssd1 vccd1 vccd1 _03478_ sky130_fd_sc_hd__nor2_1
XFILLER_0_176_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06637__B1 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08275_ net298 _02899_ vssd1 vssd1 vccd1 vccd1 _03411_ sky130_fd_sc_hd__nand2_1
XFILLER_0_34_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07226_ net794 _02361_ _02364_ _02330_ net804 vssd1 vssd1 vccd1 vccd1 _02365_ sky130_fd_sc_hd__o32a_1
XFILLER_0_6_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07157_ top.DUT.register\[2\]\[11\] net742 net718 top.DUT.register\[19\]\[11\] _02295_
+ vssd1 vssd1 vccd1 vccd1 _02296_ sky130_fd_sc_hd__a221o_1
XFILLER_0_132_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12899__RESET_B net1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_91_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07062__B1 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07088_ top.DUT.register\[6\]\[16\] net568 net452 top.DUT.register\[29\]\[16\] _02226_
+ vssd1 vssd1 vccd1 vccd1 _02227_ sky130_fd_sc_hd__a221o_1
XANTENNA__10305__S net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_4_1__f_clk clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_1__leaf_clk sky130_fd_sc_hd__clkbuf_16
Xfanout132 net135 vssd1 vssd1 vccd1 vccd1 net132 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08960__A1_N net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout143 _04946_ vssd1 vssd1 vccd1 vccd1 net143 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout154 net155 vssd1 vssd1 vccd1 vccd1 net154 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout570_X net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout165 net166 vssd1 vssd1 vccd1 vccd1 net165 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout668_X net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout176 net179 vssd1 vssd1 vccd1 vccd1 net176 sky130_fd_sc_hd__clkbuf_2
Xfanout187 _04832_ vssd1 vssd1 vccd1 vccd1 net187 sky130_fd_sc_hd__clkbuf_2
Xfanout198 _04788_ vssd1 vssd1 vccd1 vccd1 net198 sky130_fd_sc_hd__buf_2
XFILLER_0_198_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09729_ _03569_ net403 net488 _04756_ vssd1 vssd1 vccd1 vccd1 _04757_ sky130_fd_sc_hd__o211a_2
XANTENNA__08975__A1_N _03141_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12740_ clknet_leaf_37_clk _00332_ net1051 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[7\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10040__S net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06876__B1 net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_139_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12671_ clknet_leaf_10_clk _00263_ net949 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[5\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_96_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_166_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11622_ _05502_ _05504_ vssd1 vssd1 vccd1 vccd1 _05505_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_13_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_1949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06628__B1 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09130__A net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11553_ _05392_ _05400_ vssd1 vssd1 vccd1 vccd1 _05436_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_181_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_42_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10504_ net1669 net235 net357 vssd1 vssd1 vccd1 vccd1 _00673_ sky130_fd_sc_hd__mux2_1
XFILLER_0_162_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_190_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11484_ _05335_ _05340_ _05357_ vssd1 vssd1 vccd1 vccd1 _05367_ sky130_fd_sc_hd__and3_1
XANTENNA__07840__A2 net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_133_2437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13223_ clknet_leaf_5_clk _00815_ net937 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[22\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_133_2448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10435_ net253 net1839 net365 vssd1 vssd1 vccd1 vccd1 _00606_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07585__A _02723_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07053__B1 net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13154_ clknet_leaf_9_clk _00746_ net949 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[20\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_10366_ net1963 net257 net375 vssd1 vssd1 vccd1 vccd1 _00541_ sky130_fd_sc_hd__mux2_1
XFILLER_0_209_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12105_ _05984_ _05987_ vssd1 vssd1 vccd1 vccd1 _05988_ sky130_fd_sc_hd__nor2_1
XANTENNA__10215__S net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13085_ clknet_leaf_119_clk _00677_ net930 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[18\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_10297_ net269 net1721 net382 vssd1 vssd1 vccd1 vccd1 _00474_ sky130_fd_sc_hd__mux2_1
X_12036_ _05914_ _05915_ _05906_ _05908_ vssd1 vssd1 vccd1 vccd1 _05919_ sky130_fd_sc_hd__o211a_2
XANTENNA__08687__Y _03807_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06488__X _01627_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_211 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_144_2599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09024__B _02048_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12938_ clknet_leaf_118_clk _00530_ net954 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[13\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_157_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10885__S net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_185_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12869_ clknet_leaf_33_clk _00461_ net1043 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[11\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_185_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_173_603 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_177_3098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_173_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06390_ top.a1.instruction\[17\] top.a1.instruction\[18\] _01511_ _01523_ vssd1 vssd1
+ vccd1 vccd1 _01529_ sky130_fd_sc_hd__and4_1
XANTENNA__09805__B1 net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_87 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08060_ _03197_ _03198_ vssd1 vssd1 vccd1 vccd1 _03199_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_190_3298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07831__A2 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07011_ top.DUT.register\[20\]\[20\] net565 net549 top.DUT.register\[18\]\[20\] vssd1
+ vssd1 vccd1 vccd1 _02150_ sky130_fd_sc_hd__a22o_1
X_13831__1115 vssd1 vssd1 vccd1 vccd1 _13831__1115/HI net1115 sky130_fd_sc_hd__conb_1
XFILLER_0_141_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06670__Y _01809_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07044__B1 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06398__A2 net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13647__D net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08962_ _02045_ net692 net1134 net875 vssd1 vssd1 vccd1 vccd1 _00068_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__10125__S net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_164_2909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07913_ net318 _02849_ _03051_ vssd1 vssd1 vccd1 vccd1 _03052_ sky130_fd_sc_hd__o21ai_1
X_08893_ net320 _03671_ _03536_ vssd1 vssd1 vccd1 vccd1 _04003_ sky130_fd_sc_hd__o21a_1
XFILLER_0_75_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout196_A _04788_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07844_ top.DUT.register\[9\]\[0\] net467 net530 top.DUT.register\[26\]\[0\] _02982_
+ vssd1 vssd1 vccd1 vccd1 _02983_ sky130_fd_sc_hd__a221o_1
XFILLER_0_166_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07898__A2 net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_197_3408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07775_ top.DUT.register\[5\]\[2\] net651 _02913_ vssd1 vssd1 vccd1 vccd1 _02914_
+ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_104_2005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout363_A net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06570__A2 net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09514_ net133 _04555_ _04564_ _04565_ vssd1 vssd1 vccd1 vccd1 _04566_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__13780__RESET_B net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06726_ top.DUT.register\[8\]\[25\] net639 net734 top.DUT.register\[16\]\[25\] _01864_
+ vssd1 vssd1 vccd1 vccd1 _01865_ sky130_fd_sc_hd__a221o_1
XANTENNA__08847__A1 net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06858__B1 net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09445_ _02070_ _04499_ vssd1 vssd1 vccd1 vccd1 _04501_ sky130_fd_sc_hd__or2_1
X_06657_ top.DUT.register\[29\]\[26\] net454 net450 top.DUT.register\[21\]\[26\] _01795_
+ vssd1 vssd1 vccd1 vccd1 _01796_ sky130_fd_sc_hd__a221o_1
XFILLER_0_176_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10795__S net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09869__B _04560_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout628_A _04948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09376_ _04423_ _04424_ _04421_ vssd1 vssd1 vccd1 vccd1 _04436_ sky130_fd_sc_hd__o21ai_2
X_06588_ top.DUT.register\[8\]\[28\] net642 net729 top.DUT.register\[18\]\[28\] vssd1
+ vssd1 vccd1 vccd1 _01727_ sky130_fd_sc_hd__a22o_1
XFILLER_0_163_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12295__B net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08327_ net1915 net830 net800 _03461_ vssd1 vssd1 vccd1 vccd1 _00022_ sky130_fd_sc_hd__a22o_1
XFILLER_0_164_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_623 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_201_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09885__A net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07283__B1 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08258_ _03275_ _03279_ net293 vssd1 vssd1 vccd1 vccd1 _03394_ sky130_fd_sc_hd__mux2_1
XANTENNA__07822__A2 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_201_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout997_A net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07209_ _01484_ _01487_ _01588_ _02332_ _02338_ vssd1 vssd1 vccd1 vccd1 _02348_ sky130_fd_sc_hd__o221a_1
X_08189_ net288 _03324_ _03326_ vssd1 vssd1 vccd1 vccd1 _03327_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_115_2167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_2178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10220_ net177 net2161 net394 vssd1 vssd1 vccd1 vccd1 _00400_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout785_X net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10151_ net1342 net253 net602 vssd1 vssd1 vccd1 vccd1 _00350_ sky130_fd_sc_hd__mux2_1
XANTENNA__10035__S net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09109__B _02952_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10082_ net2169 net263 net612 vssd1 vssd1 vccd1 vccd1 _00283_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout952_X net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07889__A2 net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06468__B top.a1.instruction\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13772_ clknet_leaf_99_clk _01343_ vssd1 vssd1 vccd1 vccd1 top.lcd.cnt_500hz\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_186_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10984_ top.a1.dataInTemp\[5\] net785 vssd1 vssd1 vccd1 vccd1 _05022_ sky130_fd_sc_hd__or2_1
XANTENNA__06849__B1 net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_186_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_167_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12723_ clknet_leaf_124_clk _00315_ net926 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[7\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_44_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12654_ clknet_leaf_41_clk _00246_ net1056 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[4\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11605_ _05485_ _05486_ _05480_ vssd1 vssd1 vccd1 vccd1 _05488_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_127_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12585_ clknet_leaf_51_clk _00177_ net1035 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[2\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_154_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11536_ top.a1.dataIn\[14\] _05416_ _05417_ vssd1 vssd1 vccd1 vccd1 _05419_ sky130_fd_sc_hd__or3_1
XFILLER_0_108_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07274__B1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11467_ _05319_ _05325_ vssd1 vssd1 vccd1 vccd1 _05350_ sky130_fd_sc_hd__and2_1
Xmax_cap129 _05800_ vssd1 vssd1 vccd1 vccd1 net129 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_150_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07026__B1 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13206_ clknet_leaf_3_clk _00798_ net940 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[22\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_10418_ net1417 net195 net371 vssd1 vssd1 vccd1 vccd1 _00590_ sky130_fd_sc_hd__mux2_1
X_11398_ _05246_ _05250_ _05280_ vssd1 vssd1 vccd1 vccd1 _05281_ sky130_fd_sc_hd__o21ai_1
X_13137_ clknet_leaf_111_clk _00729_ net988 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[20\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_10349_ net1888 _04841_ net378 vssd1 vssd1 vccd1 vccd1 _00525_ sky130_fd_sc_hd__mux2_1
XFILLER_0_209_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09734__S net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13068_ clknet_leaf_63_clk _00660_ net1090 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[17\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_209_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_146_2639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12019_ _05854_ _05878_ vssd1 vssd1 vccd1 vccd1 _05902_ sky130_fd_sc_hd__nand2_1
XFILLER_0_205_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_179_3127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06552__A2 net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_179_3138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07560_ top.DUT.register\[22\]\[7\] net647 net762 top.DUT.register\[9\]\[7\] _02698_
+ vssd1 vssd1 vccd1 vccd1 _02699_ sky130_fd_sc_hd__a221o_1
XFILLER_0_76_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12617__CLK clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06511_ top.DUT.register\[5\]\[30\] net653 net735 top.DUT.register\[16\]\[30\] vssd1
+ vssd1 vccd1 vccd1 _01650_ sky130_fd_sc_hd__a22o_1
XFILLER_0_88_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_186_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07491_ top.DUT.register\[9\]\[14\] net468 net561 top.DUT.register\[2\]\[14\] vssd1
+ vssd1 vccd1 vccd1 _02630_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_192_3327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_463 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09230_ _04287_ _04290_ _04288_ vssd1 vssd1 vccd1 vccd1 _04298_ sky130_fd_sc_hd__a21o_1
XANTENNA__13120__RESET_B net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06442_ net804 net820 vssd1 vssd1 vccd1 vccd1 _01581_ sky130_fd_sc_hd__nand2_1
XFILLER_0_152_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06394__A top.a1.instruction\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09161_ net133 _04229_ _04233_ vssd1 vssd1 vccd1 vccd1 _04234_ sky130_fd_sc_hd__o21ai_1
X_06373_ top.a1.instruction\[15\] top.a1.instruction\[16\] net782 vssd1 vssd1 vccd1
+ vccd1 _01512_ sky130_fd_sc_hd__and3b_2
XFILLER_0_84_792 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_239 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08112_ _02498_ net331 vssd1 vssd1 vccd1 vccd1 _03251_ sky130_fd_sc_hd__or2_1
XANTENNA__09909__S net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07265__B1 net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09092_ _01505_ _04165_ _04166_ vssd1 vssd1 vccd1 vccd1 _04167_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_211_3611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_211_3622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_211_3633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_486 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08043_ _03160_ _03163_ vssd1 vssd1 vccd1 vccd1 _03182_ sky130_fd_sc_hd__nand2_4
XFILLER_0_114_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold900 top.DUT.register\[18\]\[25\] vssd1 vssd1 vccd1 vccd1 net2016 sky130_fd_sc_hd__dlygate4sd3_1
Xhold911 top.pad.keyCode\[0\] vssd1 vssd1 vccd1 vccd1 net2027 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold922 top.DUT.register\[6\]\[5\] vssd1 vssd1 vccd1 vccd1 net2038 sky130_fd_sc_hd__dlygate4sd3_1
Xhold933 top.DUT.register\[13\]\[19\] vssd1 vssd1 vccd1 vccd1 net2049 sky130_fd_sc_hd__dlygate4sd3_1
Xhold944 top.DUT.register\[7\]\[5\] vssd1 vssd1 vccd1 vccd1 net2060 sky130_fd_sc_hd__dlygate4sd3_1
Xhold955 top.DUT.register\[23\]\[7\] vssd1 vssd1 vccd1 vccd1 net2071 sky130_fd_sc_hd__dlygate4sd3_1
Xhold966 top.DUT.register\[1\]\[7\] vssd1 vssd1 vccd1 vccd1 net2082 sky130_fd_sc_hd__dlygate4sd3_1
Xhold977 top.a1.row2\[2\] vssd1 vssd1 vccd1 vccd1 net2093 sky130_fd_sc_hd__dlygate4sd3_1
Xhold988 top.ramload\[31\] vssd1 vssd1 vccd1 vccd1 net2104 sky130_fd_sc_hd__dlygate4sd3_1
X_09994_ net198 net2108 net624 vssd1 vssd1 vccd1 vccd1 _00199_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout1020_A net1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold999 top.DUT.register\[8\]\[25\] vssd1 vssd1 vccd1 vccd1 net2115 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_86_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08945_ _03019_ net691 net1176 net874 vssd1 vssd1 vccd1 vccd1 _00051_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_86_94 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_2097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout480_A _04964_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_209_3584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10324__A0 net156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08876_ _01743_ net501 _03986_ vssd1 vssd1 vccd1 vccd1 _03987_ sky130_fd_sc_hd__a21o_2
XANTENNA__08120__Y _03259_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07827_ top.DUT.register\[4\]\[0\] net667 net774 top.DUT.register\[13\]\[0\] vssd1
+ vssd1 vccd1 vccd1 _02966_ sky130_fd_sc_hd__a22o_1
XFILLER_0_169_706 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06543__A2 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout366_X net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout745_A _01623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07758_ top.DUT.register\[9\]\[3\] net468 net545 top.DUT.register\[16\]\[3\] _02896_
+ vssd1 vssd1 vccd1 vccd1 _02897_ sky130_fd_sc_hd__a221o_1
XFILLER_0_67_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_196_547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06709_ top.DUT.register\[8\]\[25\] net539 net523 top.DUT.register\[11\]\[25\] vssd1
+ vssd1 vccd1 vccd1 _01848_ sky130_fd_sc_hd__a22o_1
XFILLER_0_79_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09599__B _04644_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08296__A2 net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout533_X net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07689_ net807 _02827_ vssd1 vssd1 vccd1 vccd1 _02828_ sky130_fd_sc_hd__or2_1
XFILLER_0_183_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09428_ _04483_ _04484_ vssd1 vssd1 vccd1 vccd1 _04485_ sky130_fd_sc_hd__and2b_1
XFILLER_0_192_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_192_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09359_ net805 _02774_ _04419_ vssd1 vssd1 vccd1 vccd1 _04420_ sky130_fd_sc_hd__a21oi_4
XANTENNA_fanout700_X net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_164_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_2207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08008__B top.a1.instruction\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_656 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07256__B1 net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12370_ clknet_leaf_103_clk top.ru.next_FetchedData\[14\] net974 vssd1 vssd1 vccd1
+ vccd1 top.a1.dataIn\[14\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_34_155 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_185_Right_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11321_ top.a1.dataIn\[26\] top.a1.dataIn\[27\] top.a1.dataIn\[29\] top.a1.dataIn\[28\]
+ vssd1 vssd1 vccd1 vccd1 _05204_ sky130_fd_sc_hd__or4_1
XANTENNA__07008__B1 net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11252_ net878 net880 top.lcd.nextState\[0\] _05118_ vssd1 vssd1 vccd1 vccd1 _05145_
+ sky130_fd_sc_hd__and4_1
XANTENNA__08024__A _03162_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13638__Q top.lcd.nextState\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10203_ net242 net2079 net393 vssd1 vssd1 vccd1 vccd1 _00383_ sky130_fd_sc_hd__mux2_1
X_11183_ net1263 net587 net473 _05099_ vssd1 vssd1 vccd1 vccd1 _01240_ sky130_fd_sc_hd__a22o_1
X_10134_ net193 net1973 net610 vssd1 vssd1 vccd1 vccd1 _00334_ sky130_fd_sc_hd__mux2_1
XANTENNA__08771__A3 _03530_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10065_ net1903 net205 net617 vssd1 vssd1 vccd1 vccd1 _00267_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_128_2369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09720__A2 net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06534__A2 net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06198__B net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13824_ net1108 vssd1 vssd1 vccd1 vccd1 gpio_out[23] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_3_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13830__1114 vssd1 vssd1 vccd1 vccd1 _13830__1114/HI net1114 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_141_2558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09142__X _04216_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13755_ clknet_leaf_99_clk _01326_ vssd1 vssd1 vccd1 vccd1 top.lcd.cnt_20ms\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_10967_ top.a1.halfData\[1\] _04998_ vssd1 vssd1 vccd1 vccd1 _05009_ sky130_fd_sc_hd__or2_1
XANTENNA__09484__A1 top.pc\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12706_ clknet_leaf_9_clk _00298_ net948 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[6\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07495__B1 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10898_ net2199 net227 net478 vssd1 vssd1 vccd1 vccd1 _01059_ sky130_fd_sc_hd__mux2_1
X_13686_ clknet_leaf_89_clk _01262_ net1003 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08161__A1_N net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_174_3057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07103__A _02232_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12717__Q top.DUT.register\[6\]\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_183_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12637_ clknet_leaf_127_clk _00229_ net930 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[4\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12568_ clknet_leaf_128_clk _00160_ net912 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[2\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09787__A2 _04420_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_156_2790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_155 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11519_ _05376_ _05401_ vssd1 vssd1 vccd1 vccd1 _05402_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_152_Right_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12499_ clknet_leaf_82_clk _00091_ net993 vssd1 vssd1 vccd1 vccd1 top.pc\[11\] sky130_fd_sc_hd__dfrtp_2
Xhold207 top.DUT.register\[6\]\[22\] vssd1 vssd1 vccd1 vccd1 net1323 sky130_fd_sc_hd__dlygate4sd3_1
Xhold218 top.DUT.register\[11\]\[25\] vssd1 vssd1 vccd1 vccd1 net1334 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold229 top.DUT.register\[30\]\[24\] vssd1 vssd1 vccd1 vccd1 net1345 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout709 _01640_ vssd1 vssd1 vccd1 vccd1 net709 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_0_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13719__RESET_B net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_13_Left_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06991_ _02125_ _02127_ _02129_ vssd1 vssd1 vccd1 vccd1 _02130_ sky130_fd_sc_hd__or3_1
XANTENNA__06773__A2 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08730_ _03334_ _03832_ _03835_ _03847_ vssd1 vssd1 vccd1 vccd1 _03848_ sky130_fd_sc_hd__a211o_1
XANTENNA__10403__S net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08661_ _03264_ _03772_ _03777_ _03169_ _03781_ vssd1 vssd1 vccd1 vccd1 _03782_ sky130_fd_sc_hd__o221a_1
XANTENNA__06525__A2 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07612_ _02724_ _02749_ vssd1 vssd1 vccd1 vccd1 _02751_ sky130_fd_sc_hd__and2_1
X_08592_ _03628_ _03715_ net313 vssd1 vssd1 vccd1 vccd1 _03716_ sky130_fd_sc_hd__mux2_1
XFILLER_0_163_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07543_ _01580_ _02680_ _02681_ net806 top.a1.instruction\[28\] vssd1 vssd1 vccd1
+ vccd1 _02682_ sky130_fd_sc_hd__a32o_2
XFILLER_0_158_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_22_Left_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07474_ _02590_ _02610_ vssd1 vssd1 vccd1 vccd1 _02613_ sky130_fd_sc_hd__nor2_1
XANTENNA__08109__A _02329_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09213_ net898 top.pc\[7\] net889 vssd1 vssd1 vccd1 vccd1 _04283_ sky130_fd_sc_hd__o21ai_1
X_06425_ net683 _01523_ _01531_ vssd1 vssd1 vccd1 vccd1 _01564_ sky130_fd_sc_hd__and3_4
XANTENNA__09227__A1 net139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_173_263 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_431 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07238__B1 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09144_ _04195_ _04197_ _04217_ vssd1 vssd1 vccd1 vccd1 _04218_ sky130_fd_sc_hd__nand3_1
X_06356_ top.pad.button_control.r_counter\[0\] top.pad.button_control.r_counter\[8\]
+ top.pad.button_control.r_counter\[6\] top.pad.button_control.r_counter\[2\] vssd1
+ vssd1 vccd1 vccd1 _01496_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_20_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09075_ top.a1.instruction\[5\] net820 vssd1 vssd1 vccd1 vccd1 _04150_ sky130_fd_sc_hd__nor2_2
X_06287_ top.lcd.nextState\[5\] net815 net813 top.lcd.currentState\[5\] net1084 vssd1
+ vssd1 vccd1 vccd1 _01448_ sky130_fd_sc_hd__o221ai_4
X_08026_ net333 _03142_ _03158_ _03162_ vssd1 vssd1 vccd1 vccd1 _03165_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_112_2126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold730 top.DUT.register\[4\]\[10\] vssd1 vssd1 vccd1 vccd1 net1846 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_96_1881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_96_1892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold741 top.DUT.register\[25\]\[24\] vssd1 vssd1 vccd1 vccd1 net1857 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12362__Q top.a1.dataIn\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout695_A net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold752 top.DUT.register\[3\]\[8\] vssd1 vssd1 vccd1 vccd1 net1868 sky130_fd_sc_hd__dlygate4sd3_1
Xhold763 top.DUT.register\[21\]\[2\] vssd1 vssd1 vccd1 vccd1 net1879 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_31_Left_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10661__X _04993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold774 top.DUT.register\[9\]\[7\] vssd1 vssd1 vccd1 vccd1 net1890 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold785 top.DUT.register\[27\]\[8\] vssd1 vssd1 vccd1 vccd1 net1901 sky130_fd_sc_hd__dlygate4sd3_1
Xhold796 top.DUT.register\[8\]\[31\] vssd1 vssd1 vccd1 vccd1 net1912 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07410__B1 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09977_ _04155_ _04708_ vssd1 vssd1 vccd1 vccd1 _04949_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout483_X net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout862_A net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06764__A2 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08928_ net313 _03957_ _04035_ net285 vssd1 vssd1 vccd1 vccd1 _04036_ sky130_fd_sc_hd__o211ai_1
XANTENNA__10313__S net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout650_X net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08859_ _03969_ _03970_ net883 top.pc\[27\] vssd1 vssd1 vccd1 vccd1 _03971_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA_fanout748_X net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_207_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11870_ top.a1.dataIn\[5\] _05751_ vssd1 vssd1 vccd1 vccd1 _05753_ sky130_fd_sc_hd__nor2_1
XFILLER_0_211_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10821_ net152 net1790 net600 vssd1 vssd1 vccd1 vccd1 _00982_ sky130_fd_sc_hd__mux2_1
XFILLER_0_157_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_40_Left_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_123_2288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09897__X _04906_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13540_ clknet_leaf_94_clk _01127_ net982 vssd1 vssd1 vccd1 vccd1 top.ramload\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07477__B1 net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10752_ net1857 net173 net419 vssd1 vssd1 vccd1 vccd1 _00913_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08019__A _01589_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13471_ clknet_leaf_24_clk _01063_ net1015 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[30\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_10683_ net1622 net194 net341 vssd1 vssd1 vccd1 vccd1 _00846_ sky130_fd_sc_hd__mux2_1
XFILLER_0_180_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09218__A1 top.pc\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07229__B1 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12422_ clknet_leaf_88_clk _00018_ net1001 vssd1 vssd1 vccd1 vccd1 top.ramaddr\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_124_105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08306__X _03441_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_180_778 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12353_ clknet_leaf_88_clk net1301 net1001 vssd1 vssd1 vccd1 vccd1 top.edg2.flip2
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_133_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_283 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11304_ top.a1.row1\[109\] _05178_ _05191_ _05117_ vssd1 vssd1 vccd1 vccd1 _05192_
+ sky130_fd_sc_hd__a211o_1
X_12284_ top.lcd.cnt_500hz\[11\] _01438_ _06097_ vssd1 vssd1 vccd1 vccd1 _06101_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_39_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11099__B net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11235_ top.lcd.nextState\[5\] top.lcd.nextState\[4\] vssd1 vssd1 vccd1 vccd1 _05128_
+ sky130_fd_sc_hd__nor2_2
XFILLER_0_120_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07401__B1 net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06204__B2 net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11166_ top.a1.row1\[59\] _05092_ _05085_ vssd1 vssd1 vccd1 vccd1 _01230_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_8_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06755__A2 net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10117_ net258 net2005 net609 vssd1 vssd1 vccd1 vccd1 _00317_ sky130_fd_sc_hd__mux2_1
XANTENNA__10223__S net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11097_ net70 net864 vssd1 vssd1 vccd1 vccd1 _05054_ sky130_fd_sc_hd__and2_1
XFILLER_0_89_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10839__A1 net191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10048_ net1679 net268 net617 vssd1 vssd1 vccd1 vccd1 _00250_ sky130_fd_sc_hd__mux2_1
XFILLER_0_203_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold90 _01176_ vssd1 vssd1 vccd1 vccd1 net1206 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_203_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06496__X _01635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13807_ clknet_leaf_69_clk _01376_ net1097 vssd1 vssd1 vccd1 vccd1 top.pad.keyCode\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11999_ _05881_ vssd1 vssd1 vccd1 vccd1 _05882_ sky130_fd_sc_hd__inv_2
XANTENNA__07468__B1 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11264__B2 _01382_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13738_ clknet_leaf_96_clk _01309_ vssd1 vssd1 vccd1 vccd1 top.a1.dataInTemp\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_156_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10893__S net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13669_ clknet_leaf_92_clk _01245_ net996 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[122\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08680__A2 _03185_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_156_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06210_ net1224 net859 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedInstr\[4\] sky130_fd_sc_hd__and2_1
XANTENNA__06691__A1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_154_2749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07190_ _02319_ _02328_ vssd1 vssd1 vccd1 vccd1 _02329_ sky130_fd_sc_hd__nor2_8
XANTENNA__11016__B2 top.ramload\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06141_ net2221 vssd1 vssd1 vccd1 vccd1 _01384_ sky130_fd_sc_hd__inv_2
XANTENNA__10194__A net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09090__C1 _04164_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08432__A2 net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06443__B2 top.a1.instruction\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07640__B1 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_187_3248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09900_ top.pc\[28\] _04605_ vssd1 vssd1 vccd1 vccd1 _04908_ sky130_fd_sc_hd__or2_1
Xfanout506 _01567_ vssd1 vssd1 vccd1 vccd1 net506 sky130_fd_sc_hd__buf_4
XFILLER_0_6_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09831_ _04842_ _04843_ _04844_ _04151_ vssd1 vssd1 vccd1 vccd1 _04846_ sky130_fd_sc_hd__a31o_1
Xfanout517 _01558_ vssd1 vssd1 vccd1 vccd1 net517 sky130_fd_sc_hd__clkbuf_8
XANTENNA__09932__A2 net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_169_2981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout528 net530 vssd1 vssd1 vccd1 vccd1 net528 sky130_fd_sc_hd__clkbuf_8
Xfanout539 _01540_ vssd1 vssd1 vccd1 vccd1 net539 sky130_fd_sc_hd__clkbuf_8
XANTENNA__06746__A2 net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10133__S net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_206_3532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12955__CLK clknet_leaf_120_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09762_ top.pc\[14\] _04386_ vssd1 vssd1 vccd1 vccd1 _04784_ sky130_fd_sc_hd__xnor2_1
X_06974_ top.DUT.register\[7\]\[23\] net660 net747 top.DUT.register\[17\]\[23\] vssd1
+ vssd1 vccd1 vccd1 _02113_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_206_3543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09145__B1 _04217_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08713_ _02178_ _03810_ _02177_ vssd1 vssd1 vccd1 vccd1 _03831_ sky130_fd_sc_hd__a21oi_1
X_09693_ top.a1.dataIn\[2\] _01489_ _01503_ _01406_ vssd1 vssd1 vccd1 vccd1 _04727_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout276_A net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08644_ net885 top.pc\[17\] net696 _03765_ vssd1 vssd1 vccd1 vccd1 _03766_ sky130_fd_sc_hd__a22o_1
XFILLER_0_96_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09223__A _02497_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08575_ _03659_ _03699_ _02431_ vssd1 vssd1 vccd1 vccd1 _03700_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_25_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09448__A1 net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193_303 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout443_A _01564_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09448__B2 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07526_ top.DUT.register\[2\]\[7\] net559 net443 top.DUT.register\[1\]\[7\] _02664_
+ vssd1 vssd1 vccd1 vccd1 _02665_ sky130_fd_sc_hd__a221o_1
XANTENNA__07459__B1 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_190_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_193_369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12357__Q top.a1.dataIn\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_764 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07457_ top.DUT.register\[1\]\[15\] net755 net703 top.DUT.register\[3\]\[15\] vssd1
+ vssd1 vccd1 vccd1 _02596_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout610_A _04956_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_548 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09877__B _04577_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout708_A _01640_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06408_ top.a1.instruction\[19\] net782 _01546_ vssd1 vssd1 vccd1 vccd1 _01547_ sky130_fd_sc_hd__and3b_4
XTAP_TAPCELL_ROW_98_1910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07388_ top.DUT.register\[17\]\[9\] net459 net443 top.DUT.register\[1\]\[9\] _02526_
+ vssd1 vssd1 vccd1 vccd1 _02527_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_98_1921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08126__X _03265_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09127_ _04188_ _04201_ _04198_ _04189_ vssd1 vssd1 vccd1 vccd1 _04202_ sky130_fd_sc_hd__a211o_1
XANTENNA__08959__B1 _02609_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06339_ top.lcd.cnt_500hz\[8\] _01438_ _01482_ top.lcd.cnt_500hz\[11\] top.lcd.cnt_500hz\[12\]
+ vssd1 vssd1 vccd1 vccd1 _01483_ sky130_fd_sc_hd__a311o_1
XANTENNA__10308__S net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_801 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09058_ _03374_ _04063_ _04131_ _04132_ vssd1 vssd1 vccd1 vccd1 _04133_ sky130_fd_sc_hd__or4_1
XFILLER_0_161_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07631__B1 net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_311 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08009_ top.a1.instruction\[22\] top.a1.instruction\[23\] _03146_ _03147_ vssd1 vssd1
+ vccd1 vccd1 _03148_ sky130_fd_sc_hd__or4_2
XANTENNA_fanout698_X net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06985__A2 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold560 top.DUT.register\[29\]\[23\] vssd1 vssd1 vccd1 vccd1 net1676 sky130_fd_sc_hd__dlygate4sd3_1
Xhold571 top.DUT.register\[23\]\[0\] vssd1 vssd1 vccd1 vccd1 net1687 sky130_fd_sc_hd__dlygate4sd3_1
X_11020_ net30 net840 _05044_ net1245 vssd1 vssd1 vccd1 vccd1 _01132_ sky130_fd_sc_hd__o22a_1
Xhold582 top.DUT.register\[17\]\[17\] vssd1 vssd1 vccd1 vccd1 net1698 sky130_fd_sc_hd__dlygate4sd3_1
Xhold593 top.DUT.register\[13\]\[29\] vssd1 vssd1 vccd1 vccd1 net1709 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11191__B1 net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout865_X net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10043__S net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09117__B _03040_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08021__B _03151_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_125_2328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12971_ clknet_leaf_45_clk _00563_ net1068 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[14\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09687__A1 top.a1.dataIn\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11922_ _05799_ net129 _05802_ _05791_ vssd1 vssd1 vccd1 vccd1 _05805_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_87_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07698__B1 net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07162__A2 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_200_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_196_152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11853_ _05716_ _05718_ _05705_ vssd1 vssd1 vccd1 vccd1 _05736_ sky130_fd_sc_hd__a21oi_2
XANTENNA__13651__Q top.a1.row1\[59\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_180 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06476__B _01607_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_640 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10804_ net211 net1819 net598 vssd1 vssd1 vccd1 vccd1 _00965_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11784_ _05665_ _05666_ vssd1 vssd1 vccd1 vccd1 _05667_ sky130_fd_sc_hd__nand2_1
XFILLER_0_95_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_171_3005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13523_ clknet_leaf_88_clk top.a1.nextHex\[1\] net1004 vssd1 vssd1 vccd1 vccd1 top.a1.hexop\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_40_clk_X clknet_leaf_40_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_171_3016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10735_ top.DUT.register\[25\]\[7\] net245 net418 vssd1 vssd1 vccd1 vccd1 _00896_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13454_ clknet_leaf_39_clk _01046_ net1055 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[29\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_180_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10666_ net1520 net257 net340 vssd1 vssd1 vccd1 vccd1 _00829_ sky130_fd_sc_hd__mux2_1
XANTENNA__07870__B1 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_192_391 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12405_ clknet_leaf_105_clk top.ru.next_FetchedInstr\[17\] net971 vssd1 vssd1 vccd1
+ vccd1 top.a1.instruction\[17\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_180_575 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10218__S net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13385_ clknet_leaf_51_clk _00977_ net1056 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[27\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_136_2479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08414__A2 _03539_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09611__A1 top.edg2.flip1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10597_ net267 net2233 net348 vssd1 vssd1 vccd1 vccd1 _00762_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12336_ top.pad.button_control.r_counter\[13\] top.pad.button_control.r_counter\[12\]
+ _06131_ vssd1 vssd1 vccd1 vccd1 _06134_ sky130_fd_sc_hd__and3_1
XFILLER_0_50_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput109 net109 vssd1 vssd1 vccd1 vccd1 STB_O sky130_fd_sc_hd__buf_2
XANTENNA__07622__B1 net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_631 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06976__A2 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12267_ top.lcd.cnt_500hz\[4\] _01436_ vssd1 vssd1 vccd1 vccd1 _06091_ sky130_fd_sc_hd__nand2_1
XFILLER_0_121_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08178__A1 _01764_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11218_ net845 _05102_ vssd1 vssd1 vccd1 vccd1 _05115_ sky130_fd_sc_hd__and2_1
X_12198_ net1122 _06025_ net688 vssd1 vssd1 vccd1 vccd1 _01305_ sky130_fd_sc_hd__mux2_1
Xoutput80 net80 vssd1 vssd1 vccd1 vccd1 DAT_O[16] sky130_fd_sc_hd__clkbuf_4
Xoutput91 net91 vssd1 vssd1 vccd1 vccd1 DAT_O[26] sky130_fd_sc_hd__clkbuf_4
XANTENNA__06728__A2 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_208_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_207_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11149_ _01393_ net810 _05079_ _05080_ net889 vssd1 vssd1 vccd1 vccd1 _01225_ sky130_fd_sc_hd__o311a_1
XTAP_TAPCELL_ROW_182_3178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09742__S net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_207_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10888__S net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06690_ _01821_ _01828_ vssd1 vssd1 vccd1 vccd1 _01829_ sky130_fd_sc_hd__nor2_1
XANTENNA__08350__A1 net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07153__A2 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08350__B2 net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_176_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_65_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_201_3462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13561__Q top.ramload\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06900__A2 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_128_clk_X clknet_leaf_128_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08360_ net305 _03359_ vssd1 vssd1 vccd1 vccd1 _03493_ sky130_fd_sc_hd__nor2_1
XANTENNA__09978__A net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07311_ top.DUT.register\[17\]\[12\] net459 net503 top.DUT.register\[27\]\[12\] vssd1
+ vssd1 vccd1 vccd1 _02450_ sky130_fd_sc_hd__a22o_1
XFILLER_0_128_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08291_ _03407_ _03426_ net302 vssd1 vssd1 vccd1 vccd1 _03427_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07242_ top.DUT.register\[25\]\[10\] net778 net655 top.DUT.register\[21\]\[10\] _02380_
+ vssd1 vssd1 vccd1 vccd1 _02381_ sky130_fd_sc_hd__a221o_1
XFILLER_0_5_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07173_ top.DUT.register\[2\]\[10\] net559 net507 top.DUT.register\[4\]\[10\] _02311_
+ vssd1 vssd1 vccd1 vccd1 _02312_ sky130_fd_sc_hd__a221o_1
XANTENNA__10128__S net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06967__A2 net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_1840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_664 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout303 net307 vssd1 vssd1 vccd1 vccd1 net303 sky130_fd_sc_hd__clkbuf_2
Xfanout314 _02924_ vssd1 vssd1 vccd1 vccd1 net314 sky130_fd_sc_hd__clkbuf_4
Xfanout325 net326 vssd1 vssd1 vccd1 vccd1 net325 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout393_A net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06719__A2 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout336 net337 vssd1 vssd1 vccd1 vccd1 net336 sky130_fd_sc_hd__clkbuf_8
Xfanout347 _04991_ vssd1 vssd1 vccd1 vccd1 net347 sky130_fd_sc_hd__buf_4
X_09814_ _04151_ _04828_ _04830_ vssd1 vssd1 vccd1 vccd1 _04831_ sky130_fd_sc_hd__o21ai_1
XANTENNA_hold1139_A net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout358 net360 vssd1 vssd1 vccd1 vccd1 net358 sky130_fd_sc_hd__buf_6
Xfanout369 net372 vssd1 vssd1 vccd1 vccd1 net369 sky130_fd_sc_hd__buf_6
XANTENNA__07961__A _03099_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07392__A2 net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10798__S net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09745_ net820 _04767_ _04768_ _04345_ net826 vssd1 vssd1 vccd1 vccd1 _04769_ sky130_fd_sc_hd__o32ai_1
XANTENNA_fanout560_A _01532_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06957_ top.DUT.register\[14\]\[23\] net585 net441 top.DUT.register\[5\]\[23\] _02095_
+ vssd1 vssd1 vccd1 vccd1 _02096_ sky130_fd_sc_hd__a221o_1
XANTENNA__09669__B2 _01505_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout279_X net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout658_A _01609_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_2047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_2058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06888_ top.DUT.register\[30\]\[18\] net760 net728 top.DUT.register\[18\]\[18\] vssd1
+ vssd1 vccd1 vccd1 _02027_ sky130_fd_sc_hd__a22o_1
X_09676_ top.a1.instruction\[9\] top.a1.instruction\[10\] net786 vssd1 vssd1 vccd1
+ vccd1 _04712_ sky130_fd_sc_hd__o21ai_4
XANTENNA__07144__A2 net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08627_ net321 _03329_ _03535_ vssd1 vssd1 vccd1 vccd1 _03749_ sky130_fd_sc_hd__a21o_1
XFILLER_0_49_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08892__A2 net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout446_X net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_204_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_120_2247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08558_ net1286 net830 net800 _03683_ vssd1 vssd1 vccd1 vccd1 _00031_ sky130_fd_sc_hd__a22o_1
XFILLER_0_76_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_610 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_829 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07509_ top.DUT.register\[8\]\[14\] net641 net744 top.DUT.register\[2\]\[14\] _02647_
+ vssd1 vssd1 vccd1 vccd1 _02648_ sky130_fd_sc_hd__a221o_1
X_08489_ net886 top.pc\[10\] net697 _03617_ vssd1 vssd1 vccd1 vccd1 _03618_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout613_X net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_252 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06583__Y _01722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09841__A1 _04514_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_1980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10520_ net2226 net172 net359 vssd1 vssd1 vccd1 vccd1 _00689_ sky130_fd_sc_hd__mux2_1
XFILLER_0_162_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07852__B1 net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07201__A net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10451_ net194 net1836 net366 vssd1 vssd1 vccd1 vccd1 _00622_ sky130_fd_sc_hd__mux2_1
XANTENNA__10038__S net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13475__RESET_B net1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07604__B1 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13170_ clknet_leaf_25_clk _00762_ net1012 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[21\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_10382_ net2162 net200 net376 vssd1 vssd1 vccd1 vccd1 _00557_ sky130_fd_sc_hd__mux2_1
XANTENNA__07921__A_N _02544_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12121_ _05994_ _06002_ _06003_ vssd1 vssd1 vccd1 vccd1 _06004_ sky130_fd_sc_hd__a21oi_2
XANTENNA__06958__A2 net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07080__A1 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07855__B _02993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12052_ _05933_ _05934_ vssd1 vssd1 vccd1 vccd1 _05935_ sky130_fd_sc_hd__and2_1
Xhold390 top.DUT.register\[6\]\[20\] vssd1 vssd1 vccd1 vccd1 net1506 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08032__A net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13646__Q top.ru.state\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11164__A0 top.a1.row1\[58\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11003_ top.a1.data\[6\] top.a1.dataInTemp\[10\] net783 vssd1 vssd1 vccd1 vccd1 _05036_
+ sky130_fd_sc_hd__mux2_1
Xfanout870 net871 vssd1 vssd1 vccd1 vccd1 net870 sky130_fd_sc_hd__buf_2
Xfanout881 net882 vssd1 vssd1 vccd1 vccd1 net881 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_205_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout892 top.testpc.en_latched vssd1 vssd1 vccd1 vccd1 net892 sky130_fd_sc_hd__buf_2
XANTENNA__06591__B1 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06758__Y _01897_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10501__S net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_82_clk_A clknet_4_6__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12954_ clknet_leaf_2_clk _00546_ net917 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[14\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1090 top.DUT.register\[16\]\[27\] vssd1 vssd1 vccd1 vccd1 net2206 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07135__A2 net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08332__B2 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11905_ _05758_ _05787_ vssd1 vssd1 vccd1 vccd1 _05788_ sky130_fd_sc_hd__nand2_1
XFILLER_0_197_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12885_ clknet_leaf_31_clk _00477_ net1023 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[12\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_114_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_47_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11836_ net130 _05718_ vssd1 vssd1 vccd1 vccd1 _05719_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_97_clk_A clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_2519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11767_ _05633_ _05649_ vssd1 vssd1 vccd1 vccd1 _05650_ sky130_fd_sc_hd__or2_1
XANTENNA__09832__A1 _04499_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_200 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_520 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13506_ clknet_leaf_11_clk _01098_ net951 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[31\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07843__B1 net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10718_ net2140 net183 net337 vssd1 vssd1 vccd1 vccd1 _00879_ sky130_fd_sc_hd__mux2_1
XFILLER_0_165_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11698_ _05567_ net163 _05575_ _05579_ vssd1 vssd1 vccd1 vccd1 _05581_ sky130_fd_sc_hd__a211o_2
XFILLER_0_36_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_151_2708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13437_ clknet_leaf_119_clk _01029_ net953 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[29\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_20_clk_A clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10649_ net201 net1962 net345 vssd1 vssd1 vccd1 vccd1 _00813_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_153_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13368_ clknet_leaf_128_clk _00960_ net911 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[27\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06949__A2 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12319_ _06122_ _06123_ vssd1 vssd1 vccd1 vccd1 _01358_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_184_3207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13299_ clknet_leaf_122_clk _00891_ net932 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[25\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_35_clk_A clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09038__A _01877_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_166_2940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07860_ net804 _02360_ _02998_ vssd1 vssd1 vccd1 vccd1 _02999_ sky130_fd_sc_hd__o21a_1
XANTENNA__08020__B1 _03152_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06811_ top.DUT.register\[8\]\[17\] net640 _01945_ _01946_ _01949_ vssd1 vssd1 vccd1
+ vccd1 _01950_ sky130_fd_sc_hd__a2111o_1
X_07791_ top.DUT.register\[22\]\[2\] net575 net551 top.DUT.register\[3\]\[2\] vssd1
+ vssd1 vccd1 vccd1 _02930_ sky130_fd_sc_hd__a22o_1
X_09530_ _04561_ _04564_ _04580_ vssd1 vssd1 vccd1 vccd1 _04581_ sky130_fd_sc_hd__nand3_1
X_06742_ top.DUT.register\[22\]\[24\] net576 net510 top.DUT.register\[4\]\[24\] vssd1
+ vssd1 vccd1 vccd1 _01881_ sky130_fd_sc_hd__a22o_1
XANTENNA__12780__RESET_B net1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10411__S net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire414_X net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09461_ _04498_ _04501_ vssd1 vssd1 vccd1 vccd1 _04516_ sky130_fd_sc_hd__nand2_1
X_06673_ top.DUT.register\[15\]\[26\] net709 net701 top.DUT.register\[31\]\[26\] vssd1
+ vssd1 vccd1 vccd1 _01812_ sky130_fd_sc_hd__a22o_1
XFILLER_0_176_612 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08412_ net500 _03517_ _03518_ net432 vssd1 vssd1 vccd1 vccd1 _03544_ sky130_fd_sc_hd__a22o_1
XFILLER_0_65_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09392_ _04447_ _04450_ vssd1 vssd1 vccd1 vccd1 _04451_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_195_3369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_35_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_667 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_191_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08343_ net282 _03476_ vssd1 vssd1 vccd1 vccd1 _03477_ sky130_fd_sc_hd__nor2_1
XFILLER_0_19_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09823__A1 _04487_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_175_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_108_clk_A clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_190_114 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_594 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08274_ net317 _03409_ _03402_ vssd1 vssd1 vccd1 vccd1 _03410_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_46_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07225_ net410 _02363_ vssd1 vssd1 vccd1 vccd1 _02364_ sky130_fd_sc_hd__nor2_1
XFILLER_0_116_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_171_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12186__A2 net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07956__A _01790_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07156_ top.DUT.register\[9\]\[11\] net762 net730 top.DUT.register\[14\]\[11\] vssd1
+ vssd1 vccd1 vccd1 _02295_ sky130_fd_sc_hd__a22o_1
XFILLER_0_30_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_5_Left_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07087_ top.DUT.register\[30\]\[16\] net580 net530 top.DUT.register\[26\]\[16\] vssd1
+ vssd1 vccd1 vccd1 _02226_ sky130_fd_sc_hd__a22o_1
XFILLER_0_100_612 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout396_X net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout775_A net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12370__Q top.a1.dataIn\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout133 net135 vssd1 vssd1 vccd1 vccd1 net133 sky130_fd_sc_hd__clkbuf_4
Xfanout144 net147 vssd1 vssd1 vccd1 vccd1 net144 sky130_fd_sc_hd__buf_2
XFILLER_0_100_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09890__B _04590_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout155 _04929_ vssd1 vssd1 vccd1 vccd1 net155 sky130_fd_sc_hd__clkbuf_2
Xfanout166 net167 vssd1 vssd1 vccd1 vccd1 net166 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07365__A2 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout177 net179 vssd1 vssd1 vccd1 vccd1 net177 sky130_fd_sc_hd__clkbuf_2
Xfanout188 net191 vssd1 vssd1 vccd1 vccd1 net188 sky130_fd_sc_hd__buf_2
XFILLER_0_199_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout199 _04788_ vssd1 vssd1 vccd1 vccd1 net199 sky130_fd_sc_hd__buf_1
XANTENNA__06573__B1 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_29_Right_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout563_X net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07989_ top.DUT.register\[23\]\[31\] net674 net657 top.DUT.register\[21\]\[31\] vssd1
+ vssd1 vccd1 vccd1 _03128_ sky130_fd_sc_hd__a22o_1
XANTENNA__10321__S net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09728_ top.pc\[8\] net799 _04754_ _04755_ vssd1 vssd1 vccd1 vccd1 _04756_ sky130_fd_sc_hd__a211o_1
XFILLER_0_97_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07117__A2 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout730_X net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09659_ _04694_ _04697_ _04698_ vssd1 vssd1 vccd1 vccd1 _04699_ sky130_fd_sc_hd__or3b_1
XANTENNA__08957__A2_N net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout828_X net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_763 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12670_ clknet_leaf_18_clk _00262_ net1030 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[5\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_77_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11621_ top.a1.dataIn\[13\] _05475_ _05476_ vssd1 vssd1 vccd1 vccd1 _05504_ sky130_fd_sc_hd__and3_1
XFILLER_0_194_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09814__A1 _04151_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_100_1939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_181_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09130__B net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11552_ _05391_ _05433_ vssd1 vssd1 vccd1 vccd1 _05435_ sky130_fd_sc_hd__xor2_1
XPHY_EDGE_ROW_38_Right_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10503_ net1408 net247 net357 vssd1 vssd1 vccd1 vccd1 _00672_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_42_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11483_ _05360_ _05365_ vssd1 vssd1 vccd1 vccd1 _05366_ sky130_fd_sc_hd__nor2_1
XFILLER_0_135_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_150_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_133_2438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13222_ clknet_leaf_39_clk _00814_ net1055 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[22\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_10434_ net256 net1609 net366 vssd1 vssd1 vccd1 vccd1 _00605_ sky130_fd_sc_hd__mux2_1
XANTENNA__13179__CLK clknet_leaf_120_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13153_ clknet_leaf_16_clk _00745_ net962 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[20\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_10365_ net1606 net261 net375 vssd1 vssd1 vccd1 vccd1 _00540_ sky130_fd_sc_hd__mux2_1
XANTENNA__08033__Y _03172_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12104_ _05975_ _05978_ _05973_ vssd1 vssd1 vccd1 vccd1 _05987_ sky130_fd_sc_hd__a21oi_1
X_13084_ clknet_leaf_0_clk _00676_ net915 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[18\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_209_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10296_ net145 net1461 net381 vssd1 vssd1 vccd1 vccd1 _00473_ sky130_fd_sc_hd__mux2_1
X_12035_ _05882_ _05916_ vssd1 vssd1 vccd1 vccd1 _05918_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_47_Right_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07356__A2 net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08553__B2 net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_148_2670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06564__B1 net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10231__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_236 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07108__A2 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12937_ clknet_leaf_51_clk _00529_ net1056 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[13\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12868_ clknet_leaf_36_clk _00460_ net1042 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[11\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_199_Right_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_177_3099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11819_ _05700_ _05701_ vssd1 vssd1 vccd1 vccd1 _05702_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_32_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09805__A1 _03787_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_56_Right_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12799_ clknet_leaf_20_clk _00391_ net1028 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[9\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07816__B1 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_153_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_190_3299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07010_ top.DUT.register\[9\]\[20\] net469 _02146_ _02148_ vssd1 vssd1 vccd1 vccd1
+ _02149_ sky130_fd_sc_hd__a211o_1
XANTENNA__12168__A2 net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_180_180 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11298__A _05182_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10406__S net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07595__A2 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08961_ _01960_ net691 net1139 net874 vssd1 vssd1 vccd1 vccd1 _00067_ sky130_fd_sc_hd__a2bb2o_1
XPHY_EDGE_ROW_65_Right_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_209_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07912_ _03050_ _02852_ vssd1 vssd1 vccd1 vccd1 _03051_ sky130_fd_sc_hd__nand2b_1
X_08892_ net284 net429 _03470_ _04001_ vssd1 vssd1 vccd1 vccd1 _04002_ sky130_fd_sc_hd__a31o_1
XANTENNA__12961__RESET_B net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_54 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07347__A2 net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09741__B1 net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07843_ top.DUT.register\[6\]\[0\] net567 net503 top.DUT.register\[27\]\[0\] vssd1
+ vssd1 vccd1 vccd1 _02982_ sky130_fd_sc_hd__a22o_1
XFILLER_0_75_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06555__B1 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_87_Left_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout189_A net191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10141__S net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07774_ top.DUT.register\[24\]\[2\] net643 net710 top.DUT.register\[11\]\[2\] _02912_
+ vssd1 vssd1 vccd1 vccd1 _02913_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_104_2006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09513_ _04544_ _04548_ _04563_ net811 vssd1 vssd1 vccd1 vccd1 _04565_ sky130_fd_sc_hd__a31oi_1
X_06725_ top.DUT.register\[1\]\[25\] net754 net727 top.DUT.register\[18\]\[25\] vssd1
+ vssd1 vccd1 vccd1 _01864_ sky130_fd_sc_hd__a22o_1
XFILLER_0_189_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout356_A _04989_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06656_ top.DUT.register\[14\]\[26\] net586 net569 top.DUT.register\[6\]\[26\] vssd1
+ vssd1 vccd1 vccd1 _01795_ sky130_fd_sc_hd__a22o_1
X_09444_ _02070_ _04499_ vssd1 vssd1 vccd1 vccd1 _04500_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_166_Right_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_74_Right_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06587_ top.DUT.register\[5\]\[28\] net654 net745 top.DUT.register\[2\]\[28\] _01725_
+ vssd1 vssd1 vccd1 vccd1 _01726_ sky130_fd_sc_hd__a221o_1
XANTENNA__09257__C1 net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09375_ _04433_ _04434_ vssd1 vssd1 vccd1 vccd1 _04435_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout523_A _01554_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08326_ net884 top.pc\[4\] net695 _03460_ vssd1 vssd1 vccd1 vccd1 _03461_ sky130_fd_sc_hd__a22o_1
XFILLER_0_62_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_163_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12365__Q top.a1.dataIn\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08257_ _03272_ _03312_ net277 vssd1 vssd1 vccd1 vccd1 _03393_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07208_ top.a1.instruction\[5\] _01473_ _01480_ _02346_ _01476_ vssd1 vssd1 vccd1
+ vccd1 _02347_ sky130_fd_sc_hd__a32o_1
Xclkbuf_3_5_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_3_5_0_clk sky130_fd_sc_hd__clkbuf_8
X_08188_ net288 _03122_ vssd1 vssd1 vccd1 vccd1 _03326_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_115_2168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07139_ top.DUT.register\[22\]\[11\] net575 _02277_ vssd1 vssd1 vccd1 vccd1 _02278_
+ sky130_fd_sc_hd__a21o_1
XANTENNA__10316__S net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_83_Right_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10150_ net1891 net255 net604 vssd1 vssd1 vccd1 vccd1 _00349_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout680_X net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06794__B1 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout778_X net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10081_ net2035 net267 net613 vssd1 vssd1 vccd1 vccd1 _00282_ sky130_fd_sc_hd__mux2_1
XANTENNA__08535__B2 net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06546__B1 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10051__S net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13771_ clknet_leaf_100_clk _01342_ vssd1 vssd1 vccd1 vccd1 top.lcd.cnt_500hz\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_97_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10983_ top.a1.data\[1\] net784 vssd1 vssd1 vccd1 vccd1 _05021_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_92_Right_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12722_ clknet_leaf_23_clk _00314_ net1014 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[7\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_44_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09141__A net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07510__A2 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_133_Right_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12653_ clknet_leaf_42_clk _00245_ net1064 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[4\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_195_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_139_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11604_ _05485_ _05486_ vssd1 vssd1 vccd1 vccd1 _05487_ sky130_fd_sc_hd__and2_1
XFILLER_0_53_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12584_ clknet_leaf_27_clk _00176_ net1008 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[2\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11535_ _05416_ _05417_ vssd1 vssd1 vccd1 vccd1 _05418_ sky130_fd_sc_hd__or2_1
XANTENNA__08191__S net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11466_ _05335_ _05341_ _05347_ vssd1 vssd1 vccd1 vccd1 _05349_ sky130_fd_sc_hd__a21o_1
XFILLER_0_33_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13205_ clknet_leaf_30_clk _00797_ net1019 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[22\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_111_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10417_ net1632 _04841_ net371 vssd1 vssd1 vccd1 vccd1 _00589_ sky130_fd_sc_hd__mux2_1
XANTENNA__10226__S net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11397_ top.a1.dataIn\[27\] _05269_ _05240_ vssd1 vssd1 vccd1 vccd1 _05280_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_96_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07577__A2 net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08774__A1 net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13136_ clknet_leaf_28_clk _00728_ net1010 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[19\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_10348_ net2049 net187 net378 vssd1 vssd1 vccd1 vccd1 _00524_ sky130_fd_sc_hd__mux2_1
XANTENNA__06785__B1 net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08849__A2_N net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13067_ clknet_leaf_46_clk _00659_ net1068 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[17\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10279_ net1332 net224 net386 vssd1 vssd1 vccd1 vccd1 _00457_ sky130_fd_sc_hd__mux2_1
XANTENNA__06499__X _01638_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_800 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07329__A2 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_146_2629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12018_ _05893_ _05894_ _05895_ _05900_ vssd1 vssd1 vccd1 vccd1 _05901_ sky130_fd_sc_hd__nor4_1
XANTENNA__06537__B1 net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_179_3128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10896__S net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08829__A2 net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06510_ top.DUT.register\[31\]\[30\] net700 _01648_ _01641_ vssd1 vssd1 vccd1 vccd1
+ _01649_ sky130_fd_sc_hd__a211o_1
X_07490_ top.DUT.register\[16\]\[14\] net545 net504 top.DUT.register\[27\]\[14\] _02628_
+ vssd1 vssd1 vccd1 vccd1 _02629_ sky130_fd_sc_hd__a221o_1
XFILLER_0_0_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07501__A2 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_192_3328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06441_ net806 net821 vssd1 vssd1 vccd1 vccd1 _01580_ sky130_fd_sc_hd__nor2_1
XFILLER_0_158_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_100_Right_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06394__B top.a1.instruction\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10628__C net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09160_ net811 _04231_ _04232_ vssd1 vssd1 vccd1 vccd1 _04233_ sky130_fd_sc_hd__or3b_1
X_06372_ top.a1.instruction\[19\] net782 vssd1 vssd1 vccd1 vccd1 _01511_ sky130_fd_sc_hd__nand2_1
XFILLER_0_28_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08111_ _03248_ _03249_ vssd1 vssd1 vccd1 vccd1 _03250_ sky130_fd_sc_hd__and2_1
XFILLER_0_71_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09091_ net894 net893 _01475_ _01488_ _04152_ vssd1 vssd1 vccd1 vccd1 _04166_ sky130_fd_sc_hd__o32a_1
XFILLER_0_44_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_211_3612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_211_3623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08042_ _03152_ _03158_ vssd1 vssd1 vccd1 vccd1 _03181_ sky130_fd_sc_hd__nand2_2
XFILLER_0_114_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_153_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold901 top.DUT.register\[1\]\[25\] vssd1 vssd1 vccd1 vccd1 net2017 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold912 top.DUT.register\[19\]\[1\] vssd1 vssd1 vccd1 vccd1 net2028 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08214__B1 net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold923 top.DUT.register\[21\]\[9\] vssd1 vssd1 vccd1 vccd1 net2039 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10136__S net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold934 top.DUT.register\[9\]\[14\] vssd1 vssd1 vccd1 vccd1 net2050 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08974__A1_N _01655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold945 top.DUT.register\[2\]\[2\] vssd1 vssd1 vccd1 vccd1 net2061 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07568__A2 net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold956 top.ramload\[9\] vssd1 vssd1 vccd1 vccd1 net2072 sky130_fd_sc_hd__dlygate4sd3_1
Xhold967 top.DUT.register\[9\]\[0\] vssd1 vssd1 vccd1 vccd1 net2083 sky130_fd_sc_hd__dlygate4sd3_1
Xhold978 top.DUT.register\[27\]\[19\] vssd1 vssd1 vccd1 vccd1 net2094 sky130_fd_sc_hd__dlygate4sd3_1
Xhold989 top.DUT.register\[29\]\[25\] vssd1 vssd1 vccd1 vccd1 net2105 sky130_fd_sc_hd__dlygate4sd3_1
X_09993_ net209 net2063 net624 vssd1 vssd1 vccd1 vccd1 _00198_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08944_ net1276 net876 _02973_ net693 vssd1 vssd1 vccd1 vccd1 _00050_ sky130_fd_sc_hd__a22o_1
XANTENNA__12351__S _00016_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_95_Left_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_209_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1013_A net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_209_3574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11116__A3 net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_2098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_209_3585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08875_ _03334_ _03975_ _03982_ net424 _03985_ vssd1 vssd1 vccd1 vccd1 _03986_ sky130_fd_sc_hd__a221o_1
XANTENNA__06528__B1 net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07826_ top.DUT.register\[1\]\[0\] net754 net718 top.DUT.register\[19\]\[0\] vssd1
+ vssd1 vccd1 vccd1 _02965_ sky130_fd_sc_hd__a22o_1
XANTENNA__07017__Y _02156_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_169_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_196_515 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout640_A _01619_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07757_ top.DUT.register\[6\]\[3\] net569 net556 top.DUT.register\[28\]\[3\] vssd1
+ vssd1 vccd1 vccd1 _02896_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout359_X net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout738_A _01624_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_420 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06708_ top.DUT.register\[17\]\[25\] net459 _01844_ _01846_ vssd1 vssd1 vccd1 vccd1
+ _01847_ sky130_fd_sc_hd__a211o_1
XFILLER_0_94_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07688_ _02813_ _02817_ _02826_ vssd1 vssd1 vccd1 vccd1 _02827_ sky130_fd_sc_hd__nor3_4
XFILLER_0_177_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13248__RESET_B net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09427_ top.pc\[20\] _04471_ vssd1 vssd1 vccd1 vccd1 _04484_ sky130_fd_sc_hd__or2_1
XFILLER_0_137_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06639_ top.DUT.register\[1\]\[27\] net756 _01776_ _01777_ vssd1 vssd1 vccd1 vccd1
+ _01778_ sky130_fd_sc_hd__a211o_1
XFILLER_0_177_795 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout905_A _01405_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06700__B1 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout526_X net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_191_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09358_ net822 _02805_ _04335_ vssd1 vssd1 vccd1 vccd1 _04419_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_164_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_2208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08309_ net321 _03441_ _03442_ _03437_ vssd1 vssd1 vccd1 vccd1 _03444_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_23_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09289_ _04352_ _02453_ vssd1 vssd1 vccd1 vccd1 _04354_ sky130_fd_sc_hd__and2b_1
XFILLER_0_105_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_167 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11320_ top.a1.dataIn\[0\] _04658_ net850 _05203_ vssd1 vssd1 vccd1 vccd1 _01273_
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_105_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_342 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11251_ top.a1.row2\[24\] _05142_ _05143_ top.a1.row2\[0\] _05141_ vssd1 vssd1 vccd1
+ vccd1 _05144_ sky130_fd_sc_hd__a221o_1
XANTENNA__08205__B1 net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07559__A2 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10202_ net254 net1425 net393 vssd1 vssd1 vccd1 vccd1 _00382_ sky130_fd_sc_hd__mux2_1
X_11182_ top.a1.data\[6\] net783 _05025_ vssd1 vssd1 vccd1 vccd1 _05099_ sky130_fd_sc_hd__o21a_1
X_10133_ net200 net2180 net610 vssd1 vssd1 vccd1 vccd1 _00333_ sky130_fd_sc_hd__mux2_1
XANTENNA__09705__B1 net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input34_A en vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10064_ net1801 net218 net617 vssd1 vssd1 vccd1 vccd1 _00266_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_202_Right_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_128_2359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06479__B top.a1.instruction\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_307 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13367__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07731__A2 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13823_ net1107 vssd1 vssd1 vccd1 vccd1 gpio_out[18] sky130_fd_sc_hd__buf_2
XFILLER_0_106_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_141_2559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13754_ clknet_leaf_99_clk _01325_ vssd1 vssd1 vccd1 vccd1 top.lcd.cnt_20ms\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_10966_ top.a1.halfData\[1\] _04667_ _05007_ net844 vssd1 vssd1 vccd1 vccd1 _05008_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09484__A2 _04514_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12705_ clknet_leaf_16_clk _00297_ net959 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[6\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_168_795 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13685_ clknet_leaf_92_clk _01261_ net997 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_10897_ net1694 net233 net478 vssd1 vssd1 vccd1 vccd1 _01058_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_174_3058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12636_ clknet_leaf_0_clk _00228_ net915 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[4\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_183_787 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12567_ clknet_leaf_2_clk _00159_ net914 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[2\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_156_2780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_156_2791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07798__A2 net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11518_ _05396_ _05398_ _05374_ vssd1 vssd1 vccd1 vccd1 _05401_ sky130_fd_sc_hd__a21o_1
XFILLER_0_53_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12498_ clknet_leaf_94_clk _00090_ net994 vssd1 vssd1 vccd1 vccd1 top.pc\[10\] sky130_fd_sc_hd__dfrtp_2
Xhold208 top.DUT.register\[10\]\[28\] vssd1 vssd1 vccd1 vccd1 net1324 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold219 top.ramaddr\[30\] vssd1 vssd1 vccd1 vccd1 net1335 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_151_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11449_ _05287_ net278 _05297_ vssd1 vssd1 vccd1 vccd1 _05332_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_21_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12553__RESET_B net1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13119_ clknet_leaf_10_clk _00711_ net950 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[19\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_06990_ top.DUT.register\[21\]\[23\] net656 net723 top.DUT.register\[29\]\[23\] _02128_
+ vssd1 vssd1 vccd1 vccd1 _02129_ sky130_fd_sc_hd__a221o_1
XANTENNA__11295__B _05123_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07970__A2 net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13564__Q top.ramload\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08660_ _02049_ net493 _03778_ _03258_ _03780_ vssd1 vssd1 vccd1 vccd1 _03781_ sky130_fd_sc_hd__o221a_1
XANTENNA__07183__B1 net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07722__A2 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07611_ _02723_ _02749_ vssd1 vssd1 vccd1 vccd1 _02750_ sky130_fd_sc_hd__or2_1
X_08591_ _03674_ _03714_ net289 vssd1 vssd1 vccd1 vccd1 _03715_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_85_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07542_ top.a1.instruction\[28\] _01508_ net411 vssd1 vssd1 vccd1 vccd1 _02681_ sky130_fd_sc_hd__a21o_1
XFILLER_0_88_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_158_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07473_ _02611_ vssd1 vssd1 vccd1 vccd1 _02612_ sky130_fd_sc_hd__inv_2
XFILLER_0_186_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09212_ net132 _04275_ _04279_ _04281_ net899 vssd1 vssd1 vccd1 vccd1 _04282_ sky130_fd_sc_hd__o221a_1
X_06424_ top.DUT.register\[29\]\[30\] net453 net449 top.DUT.register\[21\]\[30\] _01560_
+ vssd1 vssd1 vccd1 vccd1 _01563_ sky130_fd_sc_hd__a221o_1
XFILLER_0_118_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06355_ top.pad.button_control.r_counter\[16\] top.pad.button_control.r_counter\[15\]
+ vssd1 vssd1 vccd1 vccd1 _01495_ sky130_fd_sc_hd__nand2_1
XFILLER_0_173_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09143_ _02857_ _02889_ _02898_ _04216_ vssd1 vssd1 vccd1 vccd1 _04217_ sky130_fd_sc_hd__o31ai_2
XFILLER_0_44_443 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout221_A _04766_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout319_A _02830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07789__A2 net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09074_ _02342_ _04148_ vssd1 vssd1 vccd1 vccd1 _04149_ sky130_fd_sc_hd__nand2b_2
XANTENNA__11171__A1_N top.a1.halfData\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06286_ _01332_ _01333_ vssd1 vssd1 vccd1 vccd1 _01447_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_16_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08025_ _01589_ _03152_ _03157_ vssd1 vssd1 vccd1 vccd1 _03164_ sky130_fd_sc_hd__or3_2
Xhold720 top.DUT.register\[16\]\[21\] vssd1 vssd1 vccd1 vccd1 net1836 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_112_2127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold731 top.DUT.register\[20\]\[27\] vssd1 vssd1 vccd1 vccd1 net1847 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_96_1882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold742 top.DUT.register\[4\]\[11\] vssd1 vssd1 vccd1 vccd1 net1858 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_96_1893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold753 top.DUT.register\[26\]\[12\] vssd1 vssd1 vccd1 vccd1 net1869 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09508__X _04560_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold764 top.DUT.register\[18\]\[11\] vssd1 vssd1 vccd1 vccd1 net1880 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_682 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06749__B1 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold775 top.DUT.register\[8\]\[4\] vssd1 vssd1 vccd1 vccd1 net1891 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout688_A _06049_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold786 top.DUT.register\[9\]\[31\] vssd1 vssd1 vccd1 vccd1 net1902 sky130_fd_sc_hd__dlygate4sd3_1
Xhold797 top.DUT.register\[3\]\[31\] vssd1 vssd1 vccd1 vccd1 net1913 sky130_fd_sc_hd__dlygate4sd3_1
X_09976_ net2218 net140 net629 vssd1 vssd1 vccd1 vccd1 _00184_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout1016_X net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08927_ net277 _03995_ _04034_ net307 vssd1 vssd1 vccd1 vccd1 _04035_ sky130_fd_sc_hd__a211o_1
XANTENNA__12298__A1 net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09163__A1 _01393_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout476_X net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_207_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08858_ _03951_ _03968_ net695 vssd1 vssd1 vccd1 vccd1 _03970_ sky130_fd_sc_hd__a21bo_1
XPHY_EDGE_ROW_179_Left_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07174__B1 net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08795__A _03909_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07809_ top.a1.instruction\[8\] _01474_ vssd1 vssd1 vccd1 vccd1 _02948_ sky130_fd_sc_hd__and2_1
XANTENNA__06921__B1 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08789_ _01920_ net495 _03883_ _03903_ vssd1 vssd1 vccd1 vccd1 _03904_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout643_X net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10820_ net157 net1765 net600 vssd1 vssd1 vccd1 vccd1 _00981_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_28_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_211_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_123_2289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout810_X net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10751_ net1469 net179 net419 vssd1 vssd1 vccd1 vccd1 _00912_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_579 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout908_X net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08019__B _03157_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13470_ clknet_leaf_54_clk _01062_ net1032 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[30\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_10682_ net1253 net202 net341 vssd1 vssd1 vccd1 vccd1 _00845_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_590 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_478 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_404 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12421_ clknet_leaf_68_clk _00017_ vssd1 vssd1 vccd1 vccd1 top.pad.button_control.debounce
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_125_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_180_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11013__X _05044_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12352_ clknet_leaf_70_clk top.edg2.button_i net1086 vssd1 vssd1 vccd1 vccd1 top.edg2.flip1
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__06988__B1 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13649__Q top.a1.row1\[57\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11303_ top.a1.row1\[13\] _05123_ _05131_ _05136_ top.a1.row1\[61\] vssd1 vssd1 vccd1
+ vccd1 _05191_ sky130_fd_sc_hd__a32o_1
XFILLER_0_132_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12283_ _06100_ net687 _06099_ vssd1 vssd1 vccd1 vccd1 _01345_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_39_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08729__A1 net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08729__B2 net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11234_ top.a1.row1\[16\] _05125_ _05126_ top.a1.row1\[8\] vssd1 vssd1 vccd1 vccd1
+ _05127_ sky130_fd_sc_hd__a22o_1
XFILLER_0_120_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_8_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10504__S net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11165_ _01379_ _01418_ _01410_ vssd1 vssd1 vccd1 vccd1 _05092_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_52_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10116_ net260 net2245 net609 vssd1 vssd1 vccd1 vccd1 _00316_ sky130_fd_sc_hd__mux2_1
X_11096_ net908 net1646 net863 _05053_ vssd1 vssd1 vccd1 vccd1 _01199_ sky130_fd_sc_hd__a31o_1
XANTENNA__08976__Y _04051_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10047_ net1357 net144 net615 vssd1 vssd1 vccd1 vccd1 _00249_ sky130_fd_sc_hd__mux2_1
XANTENNA__07880__Y _03019_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold80 net116 vssd1 vssd1 vccd1 vccd1 net1196 sky130_fd_sc_hd__dlygate4sd3_1
Xhold91 top.ramstore\[7\] vssd1 vssd1 vccd1 vccd1 net1207 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07704__A2 net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06912__B1 net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13806_ clknet_leaf_69_clk _01375_ net1097 vssd1 vssd1 vccd1 vccd1 top.pad.keyCode\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_67_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11998_ _05862_ net126 _05880_ vssd1 vssd1 vccd1 vccd1 _05881_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_187_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13737_ clknet_leaf_95_clk _01308_ vssd1 vssd1 vccd1 vccd1 top.a1.dataInTemp\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_10949_ net1944 net155 net592 vssd1 vssd1 vccd1 vccd1 _01110_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_158_2820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09032__C _03187_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_70_clk clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_70_clk
+ sky130_fd_sc_hd__clkbuf_8
X_13668_ clknet_leaf_91_clk _01244_ net996 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[121\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_80_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12619_ clknet_leaf_50_clk _00211_ net1059 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[3\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08417__B1 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06691__A2 _01829_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13599_ clknet_leaf_65_clk net1230 net1095 vssd1 vssd1 vccd1 vccd1 net91 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_143_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06140_ top.lcd.cnt_20ms\[6\] vssd1 vssd1 vccd1 vccd1 _01383_ sky130_fd_sc_hd__inv_2
XANTENNA__08968__B2 net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09090__B1 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13559__Q top.ramload\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10775__A1 net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06979__B1 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06443__A2 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_187_3249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07784__A net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout507 _01565_ vssd1 vssd1 vccd1 vccd1 net507 sky130_fd_sc_hd__clkbuf_8
X_09830_ _04843_ _04844_ _04842_ vssd1 vssd1 vccd1 vccd1 _04845_ sky130_fd_sc_hd__a21oi_1
Xfanout518 _01558_ vssd1 vssd1 vccd1 vccd1 net518 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10414__S net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout529 net530 vssd1 vssd1 vccd1 vccd1 net529 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_169_2982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09761_ top.pc\[13\] _04370_ _04774_ vssd1 vssd1 vccd1 vccd1 _04783_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_206_3533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06973_ _02111_ vssd1 vssd1 vccd1 vccd1 _02112_ sky130_fd_sc_hd__inv_2
X_08712_ net1703 net831 net801 _03830_ vssd1 vssd1 vccd1 vccd1 _00038_ sky130_fd_sc_hd__a22o_1
X_09692_ net1389 net268 net633 vssd1 vssd1 vccd1 vccd1 _00122_ sky130_fd_sc_hd__mux2_1
XANTENNA__07156__B1 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09504__A top.pc\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08643_ _03753_ _03760_ _03764_ vssd1 vssd1 vccd1 vccd1 _03765_ sky130_fd_sc_hd__or3_2
XANTENNA_fanout171_A _04885_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout269_A _04726_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09223__B _02502_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_194_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08574_ _02433_ _02474_ vssd1 vssd1 vccd1 vccd1 _03699_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_25_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_178_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07525_ top.DUT.register\[20\]\[7\] net563 net547 top.DUT.register\[18\]\[7\] vssd1
+ vssd1 vccd1 vccd1 _02664_ sky130_fd_sc_hd__a22o_1
XFILLER_0_193_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_193_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_61_clk clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_61_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout436_A _03168_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_592 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07456_ top.DUT.register\[17\]\[15\] net747 net739 top.DUT.register\[12\]\[15\] vssd1
+ vssd1 vccd1 vccd1 _02595_ sky130_fd_sc_hd__a22o_1
XANTENNA__08407__X _03539_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06407_ top.a1.instruction\[17\] top.a1.instruction\[18\] _01518_ vssd1 vssd1 vccd1
+ vccd1 _01546_ sky130_fd_sc_hd__and3_1
XFILLER_0_107_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_162_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_1911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_240 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07387_ top.DUT.register\[19\]\[9\] net536 net456 top.DUT.register\[25\]\[9\] vssd1
+ vssd1 vccd1 vccd1 _02526_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout603_A _04957_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_1922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08959__A1 top.ramstore\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_199_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09126_ _04199_ _04200_ vssd1 vssd1 vccd1 vccd1 _04201_ sky130_fd_sc_hd__nand2_1
XFILLER_0_72_571 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08959__B2 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06338_ top.lcd.cnt_500hz\[5\] top.lcd.cnt_500hz\[4\] top.lcd.cnt_500hz\[7\] top.lcd.cnt_500hz\[6\]
+ vssd1 vssd1 vccd1 vccd1 _01482_ sky130_fd_sc_hd__or4_1
XANTENNA__12373__Q top.a1.dataIn\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09057_ _03121_ _03264_ _03737_ _03881_ vssd1 vssd1 vccd1 vccd1 _04132_ sky130_fd_sc_hd__or4_1
X_06269_ top.ramload\[30\] net853 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedData\[30\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_102_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_660 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08008_ top.a1.instruction\[24\] top.a1.instruction\[25\] top.a1.instruction\[26\]
+ top.a1.instruction\[27\] vssd1 vssd1 vccd1 vccd1 _03147_ sky130_fd_sc_hd__or4_1
XANTENNA__09908__B1 net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold550 top.DUT.register\[19\]\[23\] vssd1 vssd1 vccd1 vccd1 net1666 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout593_X net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold561 top.DUT.register\[16\]\[8\] vssd1 vssd1 vccd1 vccd1 net1677 sky130_fd_sc_hd__dlygate4sd3_1
Xhold572 top.DUT.register\[8\]\[22\] vssd1 vssd1 vccd1 vccd1 net1688 sky130_fd_sc_hd__dlygate4sd3_1
Xhold583 top.DUT.register\[26\]\[25\] vssd1 vssd1 vccd1 vccd1 net1699 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09384__A1 net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10324__S net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold594 top.DUT.register\[10\]\[30\] vssd1 vssd1 vccd1 vccd1 net1710 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09959_ net1904 net199 net629 vssd1 vssd1 vccd1 vccd1 _00167_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout760_X net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout858_X net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12970_ clknet_leaf_120_clk _00562_ net933 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[14\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_99_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_125_2318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09687__A2 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11921_ _05803_ vssd1 vssd1 vccd1 vccd1 _05804_ sky130_fd_sc_hd__inv_2
XANTENNA__09414__A _01983_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_169_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11852_ _05726_ _05734_ vssd1 vssd1 vccd1 vccd1 _05735_ sky130_fd_sc_hd__and2_1
XFILLER_0_196_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10803_ net221 net1956 net598 vssd1 vssd1 vccd1 vccd1 _00964_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_192 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11783_ _05624_ _05662_ vssd1 vssd1 vccd1 vccd1 _05666_ sky130_fd_sc_hd__xnor2_1
Xclkbuf_leaf_52_clk clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_52_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_184_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13522_ clknet_leaf_74_clk top.a1.nextHex\[0\] net1077 vssd1 vssd1 vccd1 vccd1 _01377_
+ sky130_fd_sc_hd__dfrtp_1
X_10734_ net2251 net243 net418 vssd1 vssd1 vccd1 vccd1 _00895_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_171_3006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_171_3017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13453_ clknet_leaf_44_clk _01045_ net1063 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[29\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06673__A2 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10665_ net1870 net261 net340 vssd1 vssd1 vccd1 vccd1 _00828_ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12404_ clknet_leaf_105_clk top.ru.next_FetchedInstr\[16\] net969 vssd1 vssd1 vccd1
+ vccd1 top.a1.instruction\[16\] sky130_fd_sc_hd__dfrtp_4
X_13384_ clknet_leaf_27_clk _00976_ net1010 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[27\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10596_ net144 net2225 net346 vssd1 vssd1 vccd1 vccd1 _00761_ sky130_fd_sc_hd__mux2_1
XFILLER_0_180_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12335_ top.pad.button_control.r_counter\[12\] _06131_ top.pad.button_control.r_counter\[13\]
+ vssd1 vssd1 vccd1 vccd1 _06133_ sky130_fd_sc_hd__a21o_1
XFILLER_0_121_643 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12266_ top.lcd.cnt_500hz\[4\] _01436_ vssd1 vssd1 vccd1 vccd1 _06090_ sky130_fd_sc_hd__or2_1
X_11217_ _05114_ net1272 net471 vssd1 vssd1 vccd1 vccd1 _01259_ sky130_fd_sc_hd__mux2_1
XFILLER_0_208_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10234__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_208_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12197_ net1125 _06034_ _06049_ vssd1 vssd1 vccd1 vccd1 _01304_ sky130_fd_sc_hd__mux2_1
Xoutput70 net70 vssd1 vssd1 vccd1 vccd1 ADR_O[8] sky130_fd_sc_hd__buf_2
XFILLER_0_120_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput81 net81 vssd1 vssd1 vccd1 vccd1 DAT_O[17] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_208_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput92 net92 vssd1 vssd1 vccd1 vccd1 DAT_O[27] sky130_fd_sc_hd__clkbuf_4
X_11148_ _01388_ net898 _01503_ top.pc\[0\] vssd1 vssd1 vccd1 vccd1 _05080_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_182_3179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11079_ net96 net872 net836 net1136 vssd1 vssd1 vccd1 vccd1 _01190_ sky130_fd_sc_hd__a22o_1
XANTENNA__07138__B1 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_188_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_201_3463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09978__B _04712_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_43_clk clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_43_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__10445__A0 net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_175_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_376 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07310_ top.DUT.register\[9\]\[12\] net467 net555 top.DUT.register\[28\]\[12\] _02448_
+ vssd1 vssd1 vccd1 vccd1 _02449_ sky130_fd_sc_hd__a221o_1
X_08290_ net276 _03345_ vssd1 vssd1 vccd1 vccd1 _03426_ sky130_fd_sc_hd__or2_1
XANTENNA__07310__B1 net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_9_clk_A clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07241_ top.DUT.register\[28\]\[10\] net766 net738 top.DUT.register\[12\]\[10\] vssd1
+ vssd1 vccd1 vccd1 _02380_ sky130_fd_sc_hd__a22o_1
XFILLER_0_73_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_183_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06664__A2 net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10409__S net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07172_ top.DUT.register\[19\]\[10\] net535 net515 top.DUT.register\[7\]\[10\] vssd1
+ vssd1 vccd1 vccd1 _02311_ sky130_fd_sc_hd__a22o_1
XFILLER_0_144_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_171_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_200_Left_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_232 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07785__Y _02924_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_479 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_93_1841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08403__A net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_676 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09366__A1 net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10144__S net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout304 net306 vssd1 vssd1 vccd1 vccd1 net304 sky130_fd_sc_hd__buf_2
Xfanout315 net316 vssd1 vssd1 vccd1 vccd1 net315 sky130_fd_sc_hd__buf_2
XANTENNA__07377__B1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout326 _02829_ vssd1 vssd1 vccd1 vccd1 net326 sky130_fd_sc_hd__buf_2
XANTENNA__11173__B2 net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09933__S net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout337 _04995_ vssd1 vssd1 vccd1 vccd1 net337 sky130_fd_sc_hd__clkbuf_8
X_09813_ net828 _04463_ _04829_ vssd1 vssd1 vccd1 vccd1 _04830_ sky130_fd_sc_hd__o21ba_1
Xfanout348 _04991_ vssd1 vssd1 vccd1 vccd1 net348 sky130_fd_sc_hd__clkbuf_8
Xfanout359 net360 vssd1 vssd1 vccd1 vccd1 net359 sky130_fd_sc_hd__buf_4
XANTENNA_fanout386_A _04978_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09744_ top.pc\[12\] _04172_ _04352_ vssd1 vssd1 vccd1 vccd1 _04768_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_94_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06956_ top.DUT.register\[10\]\[23\] net520 net506 top.DUT.register\[27\]\[23\] vssd1
+ vssd1 vccd1 vccd1 _02095_ sky130_fd_sc_hd__a22o_1
XANTENNA__07129__B1 net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_2048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09675_ top.a1.instruction\[10\] net786 vssd1 vssd1 vccd1 vccd1 _04711_ sky130_fd_sc_hd__nand2_2
XANTENNA_fanout553_A _01535_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06887_ _02016_ _02025_ vssd1 vssd1 vccd1 vccd1 _02026_ sky130_fd_sc_hd__nor2_2
X_08626_ _01964_ _03747_ vssd1 vssd1 vccd1 vccd1 _03748_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_139_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12368__Q top.a1.dataIn\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_652 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08629__B1 net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08557_ net883 top.pc\[13\] net694 _03682_ vssd1 vssd1 vccd1 vccd1 _03683_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_120_2248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout720_A _01635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout341_X net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_7_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_34_clk clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_34_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout818_A net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout439_X net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1083_X net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07508_ top.DUT.register\[30\]\[14\] net760 net704 top.DUT.register\[3\]\[14\] vssd1
+ vssd1 vccd1 vccd1 _02647_ sky130_fd_sc_hd__a22o_1
XANTENNA__07689__A net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_193_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_451 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08488_ net423 _03597_ _03616_ _03334_ _03611_ vssd1 vssd1 vccd1 vccd1 _03617_ sky130_fd_sc_hd__a221o_2
XANTENNA__07301__B1 net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_102_1970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_1981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06655__A2 net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07439_ top.DUT.register\[18\]\[15\] net548 net528 top.DUT.register\[26\]\[15\] vssd1
+ vssd1 vccd1 vccd1 _02578_ sky130_fd_sc_hd__a22o_1
XFILLER_0_9_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10319__S net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12189__B1 _05083_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10450_ net200 net2092 net366 vssd1 vssd1 vccd1 vccd1 _00621_ sky130_fd_sc_hd__mux2_1
XFILLER_0_162_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09109_ top.pc\[1\] _02952_ vssd1 vssd1 vccd1 vccd1 _04184_ sky130_fd_sc_hd__nand2_1
XFILLER_0_134_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10381_ net2122 net186 net375 vssd1 vssd1 vccd1 vccd1 _00556_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12120_ _05988_ _05996_ vssd1 vssd1 vccd1 vccd1 _06003_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07080__A2 _02218_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12051_ _05907_ _05917_ vssd1 vssd1 vccd1 vccd1 _05934_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10054__S net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold380 top.DUT.register\[12\]\[29\] vssd1 vssd1 vccd1 vccd1 net1496 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_2_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold391 top.DUT.register\[31\]\[11\] vssd1 vssd1 vccd1 vccd1 net1507 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07368__B1 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08032__B net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07907__A2 _03040_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11002_ net1225 _05035_ net589 vssd1 vssd1 vccd1 vccd1 _01123_ sky130_fd_sc_hd__mux2_1
XANTENNA__08600__X _03724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout860 _01428_ vssd1 vssd1 vccd1 vccd1 net860 sky130_fd_sc_hd__clkbuf_4
Xfanout871 net872 vssd1 vssd1 vccd1 vccd1 net871 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_205_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout882 top.lcd.nextState\[1\] vssd1 vssd1 vccd1 vccd1 net882 sky130_fd_sc_hd__buf_2
XFILLER_0_189_407 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout893 top.a1.instruction\[14\] vssd1 vssd1 vccd1 vccd1 net893 sky130_fd_sc_hd__buf_2
XFILLER_0_204_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12953_ clknet_leaf_14_clk _00545_ net955 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[14\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1080 top.DUT.register\[22\]\[16\] vssd1 vssd1 vccd1 vccd1 net2196 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1091 top.DUT.register\[7\]\[26\] vssd1 vssd1 vccd1 vccd1 net2207 sky130_fd_sc_hd__dlygate4sd3_1
X_11904_ _05779_ _05781_ _05782_ _05785_ vssd1 vssd1 vccd1 vccd1 _05787_ sky130_fd_sc_hd__a31o_1
X_12884_ clknet_leaf_54_clk _00476_ net1031 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[12\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_200_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11835_ _05685_ _05687_ _05712_ _05717_ vssd1 vssd1 vccd1 vccd1 _05718_ sky130_fd_sc_hd__a31o_2
XFILLER_0_114_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06894__A2 net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_25_clk clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_25_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_68_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_2509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_488 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11766_ _05601_ _05620_ _05592_ vssd1 vssd1 vccd1 vccd1 _05649_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_55_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13505_ clknet_leaf_17_clk _01097_ net1030 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[31\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_10717_ net1592 net193 net336 vssd1 vssd1 vccd1 vccd1 _00878_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_60_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_532 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11697_ _05567_ _05573_ _05575_ _05579_ vssd1 vssd1 vccd1 vccd1 _05580_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_125_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08207__B _03122_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13436_ clknet_leaf_0_clk _01028_ net914 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[29\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_779 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_151_2709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10648_ net186 net2150 net345 vssd1 vssd1 vccd1 vccd1 _00812_ sky130_fd_sc_hd__mux2_1
XFILLER_0_141_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11849__A top.a1.dataIn\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13367_ clknet_leaf_2_clk _00959_ net914 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[27\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_10579_ net1788 net225 net351 vssd1 vssd1 vccd1 vccd1 _00745_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12318_ top.pad.button_control.r_counter\[6\] _06120_ net790 vssd1 vssd1 vccd1 vccd1
+ _06123_ sky130_fd_sc_hd__o21ai_1
XANTENNA__09319__A top.pc\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07071__A2 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_184_3208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13298_ clknet_leaf_23_clk _00890_ net1014 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[25\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09348__A1 net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12249_ top.lcd.cnt_20ms\[14\] _06079_ net978 vssd1 vssd1 vccd1 vccd1 _06081_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_139_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_166_2930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08020__A1 _01589_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_166_2941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10899__S net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08510__X _03638_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06949__Y _02088_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08877__B _03987_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06810_ top.DUT.register\[16\]\[17\] net736 _01948_ vssd1 vssd1 vccd1 vccd1 _01949_
+ sky130_fd_sc_hd__a21o_1
X_07790_ top.DUT.register\[11\]\[2\] net523 net515 top.DUT.register\[7\]\[2\] _02928_
+ vssd1 vssd1 vccd1 vccd1 _02929_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_147_Right_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11288__B1_N _05149_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06741_ top.DUT.register\[12\]\[24\] net533 net513 top.DUT.register\[24\]\[24\] _01879_
+ vssd1 vssd1 vccd1 vccd1 _01880_ sky130_fd_sc_hd__a221o_1
XANTENNA__09520__A1 top.pc\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09460_ _02198_ _04514_ vssd1 vssd1 vccd1 vccd1 _04515_ sky130_fd_sc_hd__xor2_1
X_06672_ top.DUT.register\[2\]\[26\] net745 net638 top.DUT.register\[6\]\[26\] vssd1
+ vssd1 vccd1 vccd1 _01811_ sky130_fd_sc_hd__a22o_1
X_08411_ net282 _03542_ vssd1 vssd1 vccd1 vccd1 _03543_ sky130_fd_sc_hd__or2_1
XFILLER_0_176_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09341__X _04403_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09391_ _04448_ _04449_ vssd1 vssd1 vccd1 vccd1 _04450_ sky130_fd_sc_hd__and2b_1
XANTENNA__06885__A2 net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_16_clk clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_16_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_35_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08342_ _03331_ _03475_ net312 vssd1 vssd1 vccd1 vccd1 _03476_ sky130_fd_sc_hd__mux2_1
XFILLER_0_176_679 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10139__S net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06637__A2 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08273_ net316 _03408_ _03406_ vssd1 vssd1 vccd1 vccd1 _03409_ sky130_fd_sc_hd__a21o_1
XFILLER_0_190_126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_172_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout134_A net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07224_ top.a1.instruction\[20\] _01507_ net793 net895 _02362_ vssd1 vssd1 vccd1
+ vccd1 _02363_ sky130_fd_sc_hd__a221o_1
XFILLER_0_80_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07155_ top.DUT.register\[8\]\[11\] net639 net710 top.DUT.register\[11\]\[11\] _02293_
+ vssd1 vssd1 vccd1 vccd1 _02294_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout301_A _02974_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1043_A net1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07598__B1 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07062__A2 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07086_ top.DUT.register\[21\]\[16\] net448 net444 top.DUT.register\[1\]\[16\] _02224_
+ vssd1 vssd1 vccd1 vccd1 _02225_ sky130_fd_sc_hd__a221o_1
XANTENNA__08133__A _02242_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06205__X top.ru.next_iready vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout134 net135 vssd1 vssd1 vccd1 vccd1 net134 sky130_fd_sc_hd__buf_2
XANTENNA_fanout670_A _01599_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout145 net147 vssd1 vssd1 vccd1 vccd1 net145 sky130_fd_sc_hd__buf_2
Xfanout156 _04916_ vssd1 vssd1 vccd1 vccd1 net156 sky130_fd_sc_hd__buf_2
Xfanout167 _04895_ vssd1 vssd1 vccd1 vccd1 net167 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout768_A net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout389_X net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10602__S net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout178 net179 vssd1 vssd1 vccd1 vccd1 net178 sky130_fd_sc_hd__clkbuf_2
Xfanout189 net191 vssd1 vssd1 vccd1 vccd1 net189 sky130_fd_sc_hd__clkbuf_2
X_07988_ top.DUT.register\[4\]\[31\] net669 net775 top.DUT.register\[13\]\[31\] _03126_
+ vssd1 vssd1 vccd1 vccd1 _03127_ sky130_fd_sc_hd__a221o_1
XANTENNA__07770__B1 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_114_Right_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09727_ net826 _04286_ _04752_ top.a1.dataIn\[8\] vssd1 vssd1 vccd1 vccd1 _04755_
+ sky130_fd_sc_hd__a2bb2o_1
X_06939_ top.DUT.register\[18\]\[21\] net729 _02075_ _02077_ vssd1 vssd1 vccd1 vccd1
+ _02078_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout935_A net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout556_X net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10657__A0 _04916_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09658_ _04674_ _04677_ _04678_ _04675_ vssd1 vssd1 vccd1 vccd1 _04698_ sky130_fd_sc_hd__o22a_1
XANTENNA__07522__B1 net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08609_ _03686_ _03731_ net290 vssd1 vssd1 vccd1 vccd1 _03732_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_106_Left_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_194_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06876__A2 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout723_X net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09589_ _04602_ _04615_ _04617_ _04614_ vssd1 vssd1 vccd1 vccd1 _04636_ sky130_fd_sc_hd__a31o_1
XFILLER_0_139_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_775 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11620_ _05451_ _05502_ vssd1 vssd1 vccd1 vccd1 _05503_ sky130_fd_sc_hd__xor2_1
XANTENNA__12490__RESET_B net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_194_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_13_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06628__A2 net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11551_ _05391_ _05433_ vssd1 vssd1 vccd1 vccd1 _05434_ sky130_fd_sc_hd__and2b_1
XFILLER_0_107_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10049__S net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_163_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10502_ net1947 net242 net357 vssd1 vssd1 vccd1 vccd1 _00671_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_42_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11482_ top.a1.dataIn\[15\] _05361_ _05362_ _05363_ vssd1 vssd1 vccd1 vccd1 _05365_
+ sky130_fd_sc_hd__o22a_1
X_13221_ clknet_leaf_35_clk _00813_ net1040 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[22\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09578__B2 net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10433_ net259 net1961 net367 vssd1 vssd1 vccd1 vccd1 _00604_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_133_2439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07053__A2 net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13152_ clknet_leaf_17_clk _00744_ net992 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[20\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_115_Left_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10364_ net2272 net263 net373 vssd1 vssd1 vccd1 vccd1 _00539_ sky130_fd_sc_hd__mux2_1
X_12103_ _05970_ _05981_ _05982_ vssd1 vssd1 vccd1 vccd1 _05986_ sky130_fd_sc_hd__or3_1
X_13083_ clknet_leaf_120_clk _00675_ net933 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[18\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_10295_ _04967_ net399 vssd1 vssd1 vccd1 vccd1 _04979_ sky130_fd_sc_hd__nand2b_1
XANTENNA__07882__A net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12034_ _05881_ _05916_ vssd1 vssd1 vccd1 vccd1 _05917_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_148_2660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10512__S net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_148_2671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout690 _04710_ vssd1 vssd1 vccd1 vccd1 net690 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_70_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06173__A_N top.a1.halfData\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_248 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_161_2860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12936_ clknet_leaf_27_clk _00528_ net1008 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[13\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_124_Left_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_158_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_4_8__f_clk_A clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12867_ clknet_leaf_61_clk _00459_ net1088 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[11\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12507__RESET_B net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11818_ top.a1.dataIn\[7\] _05664_ _05690_ vssd1 vssd1 vccd1 vccd1 _05701_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_32_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12798_ clknet_leaf_18_clk _00390_ net1028 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[9\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09805__A2 net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_185_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06619__A2 net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11749_ _05618_ _05630_ vssd1 vssd1 vccd1 vccd1 _05632_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_154_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09748__S net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_190_3289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13419_ clknet_leaf_48_clk _01011_ net1059 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[28\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_133_Left_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_714 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07044__A2 net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13567__Q top.ramload\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_90_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08960_ net412 net692 net1205 net874 vssd1 vssd1 vccd1 vccd1 _00066_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_121_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_5_clk clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_5_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__11128__A1 net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07911_ _02880_ _02899_ _03049_ vssd1 vssd1 vccd1 vccd1 _03050_ sky130_fd_sc_hd__a21o_1
X_08891_ _01700_ net433 net501 _01699_ _04000_ vssd1 vssd1 vccd1 vccd1 _04001_ sky130_fd_sc_hd__a221o_1
XFILLER_0_166_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09741__A1 _03638_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_66 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07842_ top.DUT.register\[22\]\[0\] net578 net456 top.DUT.register\[25\]\[0\] _02980_
+ vssd1 vssd1 vccd1 vccd1 _02981_ sky130_fd_sc_hd__a221o_1
X_07773_ top.DUT.register\[17\]\[2\] net746 net718 top.DUT.register\[19\]\[2\] vssd1
+ vssd1 vccd1 vccd1 _02912_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_142_Left_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_88_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_2007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09512_ _04544_ _04548_ _04563_ vssd1 vssd1 vccd1 vccd1 _04564_ sky130_fd_sc_hd__a21o_1
XFILLER_0_196_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06724_ top.DUT.register\[7\]\[25\] net662 net765 top.DUT.register\[9\]\[25\] vssd1
+ vssd1 vccd1 vccd1 _01863_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_88_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07504__B1 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09443_ net821 _02501_ net422 vssd1 vssd1 vccd1 vccd1 _04499_ sky130_fd_sc_hd__a21o_2
X_06655_ top.DUT.register\[12\]\[26\] net534 net461 top.DUT.register\[17\]\[26\] _01793_
+ vssd1 vssd1 vccd1 vccd1 _01794_ sky130_fd_sc_hd__a221o_1
XANTENNA__06858__A2 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_176_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12349__S _00016_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout251_A _04741_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout349_A _04991_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09374_ _04413_ _04415_ _04416_ vssd1 vssd1 vccd1 vccd1 _04434_ sky130_fd_sc_hd__a21oi_1
X_06586_ top.DUT.register\[17\]\[28\] net749 net736 top.DUT.register\[16\]\[28\] vssd1
+ vssd1 vccd1 vccd1 _01725_ sky130_fd_sc_hd__a22o_1
XFILLER_0_19_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11064__B1 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08325_ _03448_ _03455_ _03459_ vssd1 vssd1 vccd1 vccd1 _03460_ sky130_fd_sc_hd__or3_2
XFILLER_0_145_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout516_A _01558_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout137_X net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_144_340 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08256_ net1572 net832 net802 _03392_ vssd1 vssd1 vccd1 vccd1 _00020_ sky130_fd_sc_hd__a22o_1
XANTENNA__07283__A2 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_151_Left_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_201_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07207_ _02343_ _02345_ vssd1 vssd1 vccd1 vccd1 _02346_ sky130_fd_sc_hd__nand2_1
XFILLER_0_131_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_535 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08187_ _03324_ vssd1 vssd1 vccd1 vccd1 _03325_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_81_clk_A clknet_4_6__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_2169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07138_ top.DUT.register\[15\]\[11\] net679 net675 top.DUT.register\[31\]\[11\] vssd1
+ vssd1 vccd1 vccd1 _02277_ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout885_A top.ru.state\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07069_ _02202_ _02205_ _02207_ vssd1 vssd1 vccd1 vccd1 _02208_ sky130_fd_sc_hd__or3_1
XANTENNA__07991__B1 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_96_clk_A clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10080_ net2157 net147 net611 vssd1 vssd1 vccd1 vccd1 _00281_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout673_X net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11415__A1_N top.a1.dataIn\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_160_Left_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10332__S net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09406__B _04453_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07743__B1 net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout840_X net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13770_ clknet_leaf_100_clk _01341_ vssd1 vssd1 vccd1 vccd1 top.lcd.cnt_500hz\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_97_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10982_ net1145 _05020_ net590 vssd1 vssd1 vccd1 vccd1 _01118_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_143_2590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12721_ clknet_leaf_113_clk _00313_ net991 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[7\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06849__A2 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_195_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12652_ clknet_leaf_48_clk _00244_ net1060 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[4\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_155_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_238 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_34_clk_A clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08038__A net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_194_284 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11055__B1 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11603_ _05483_ _05484_ _05464_ vssd1 vssd1 vccd1 vccd1 _05486_ sky130_fd_sc_hd__o21ai_1
X_12583_ clknet_leaf_7_clk _00175_ net944 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[2\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_93_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11534_ top.a1.dataIn\[15\] _05396_ _05398_ vssd1 vssd1 vccd1 vccd1 _05417_ sky130_fd_sc_hd__and3_1
XFILLER_0_108_565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13806__RESET_B net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07274__A2 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_49_clk_A clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10507__S net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11465_ _05342_ _05343_ vssd1 vssd1 vccd1 vccd1 _05348_ sky130_fd_sc_hd__and2_1
XFILLER_0_21_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_319 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_59_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13204_ clknet_leaf_56_clk _00796_ net1073 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[22\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_10416_ net1402 net186 net371 vssd1 vssd1 vccd1 vccd1 _00588_ sky130_fd_sc_hd__mux2_1
XANTENNA__07026__A2 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11396_ _05247_ _05278_ vssd1 vssd1 vccd1 vccd1 _05279_ sky130_fd_sc_hd__xor2_1
XFILLER_0_60_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13135_ clknet_leaf_22_clk _00727_ net1024 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[19\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10347_ net1325 net203 net380 vssd1 vssd1 vccd1 vccd1 _00523_ sky130_fd_sc_hd__mux2_1
XFILLER_0_209_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_72_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13066_ clknet_leaf_120_clk _00658_ net933 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[17\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_10278_ net1987 net189 net386 vssd1 vssd1 vccd1 vccd1 _00456_ sky130_fd_sc_hd__mux2_1
X_12017_ _05871_ _05889_ _05896_ vssd1 vssd1 vccd1 vccd1 _05900_ sky130_fd_sc_hd__or3_1
XANTENNA_clkbuf_leaf_107_clk_A clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10242__S net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07734__B1 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08931__C1 _03185_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_179_3129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_177_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11294__B1 _05183_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12919_ clknet_leaf_129_clk _00511_ net911 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[13\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_201_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06440_ _01388_ net896 _01390_ _01502_ vssd1 vssd1 vccd1 vccd1 _01579_ sky130_fd_sc_hd__nand4_2
XTAP_TAPCELL_ROW_192_3329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06371_ top.a1.instruction\[19\] net782 vssd1 vssd1 vccd1 vccd1 _01510_ sky130_fd_sc_hd__and2_1
XFILLER_0_44_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08890__B net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_699 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08110_ _02286_ net328 vssd1 vssd1 vccd1 vccd1 _03249_ sky130_fd_sc_hd__nand2_1
XFILLER_0_43_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13547__RESET_B net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09090_ net895 _01589_ _02332_ net799 _04164_ vssd1 vssd1 vccd1 vccd1 _04165_ sky130_fd_sc_hd__a311o_1
XANTENNA__07265__A2 net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_211_3613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08041_ _02996_ _03172_ vssd1 vssd1 vccd1 vccd1 _03180_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_211_3624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10417__S net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold902 top.ramaddr\[1\] vssd1 vssd1 vccd1 vccd1 net2018 sky130_fd_sc_hd__dlygate4sd3_1
Xhold913 top.DUT.register\[13\]\[23\] vssd1 vssd1 vccd1 vccd1 net2029 sky130_fd_sc_hd__dlygate4sd3_1
Xhold924 top.DUT.register\[22\]\[21\] vssd1 vssd1 vccd1 vccd1 net2040 sky130_fd_sc_hd__dlygate4sd3_1
Xhold935 top.ramload\[25\] vssd1 vssd1 vccd1 vccd1 net2051 sky130_fd_sc_hd__dlygate4sd3_1
Xhold946 top.DUT.register\[21\]\[8\] vssd1 vssd1 vccd1 vccd1 net2062 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold957 top.DUT.register\[29\]\[14\] vssd1 vssd1 vccd1 vccd1 net2073 sky130_fd_sc_hd__dlygate4sd3_1
Xhold968 top.DUT.register\[3\]\[28\] vssd1 vssd1 vccd1 vccd1 net2084 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09992_ net213 net1725 net623 vssd1 vssd1 vccd1 vccd1 _00197_ sky130_fd_sc_hd__mux2_1
Xhold979 top.DUT.register\[4\]\[22\] vssd1 vssd1 vccd1 vccd1 net2095 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_177_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07973__B1 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_177_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08943_ net873 _03267_ vssd1 vssd1 vccd1 vccd1 _04050_ sky130_fd_sc_hd__or2_4
XANTENNA__09507__A net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_2099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_209_3575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10152__S net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_209_3586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08874_ net435 _03979_ _03980_ _03259_ _03984_ vssd1 vssd1 vccd1 vccd1 _03985_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout1006_A net1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07725__B1 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07825_ _02957_ _02959_ _02963_ vssd1 vssd1 vccd1 vccd1 _02964_ sky130_fd_sc_hd__or3_1
X_07756_ top.DUT.register\[11\]\[3\] net526 net506 top.DUT.register\[27\]\[3\] _02894_
+ vssd1 vssd1 vccd1 vccd1 _02895_ sky130_fd_sc_hd__a221o_1
XANTENNA__06866__A _01983_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_196_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06707_ top.DUT.register\[30\]\[25\] net579 net456 top.DUT.register\[25\]\[25\] _01845_
+ vssd1 vssd1 vccd1 vccd1 _01846_ sky130_fd_sc_hd__a221o_1
X_07687_ _02821_ _02823_ _02825_ vssd1 vssd1 vccd1 vccd1 _02826_ sky130_fd_sc_hd__or3_1
XFILLER_0_149_432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout633_A _04714_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09426_ top.pc\[20\] _04471_ vssd1 vssd1 vccd1 vccd1 _04483_ sky130_fd_sc_hd__and2_1
X_06638_ top.DUT.register\[21\]\[27\] net658 net705 top.DUT.register\[3\]\[27\] vssd1
+ vssd1 vccd1 vccd1 _01777_ sky130_fd_sc_hd__a22o_1
XFILLER_0_177_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09357_ _04413_ _04417_ vssd1 vssd1 vccd1 vccd1 _04418_ sky130_fd_sc_hd__xnor2_1
X_06569_ top.DUT.register\[9\]\[28\] net469 net461 top.DUT.register\[17\]\[28\] _01707_
+ vssd1 vssd1 vccd1 vccd1 _01708_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout421_X net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout519_X net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08308_ net321 _03441_ _03437_ vssd1 vssd1 vccd1 vccd1 _03443_ sky130_fd_sc_hd__o21a_1
XFILLER_0_34_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08008__D top.a1.instruction\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07256__A2 net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_660 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09288_ _02443_ _02452_ _04352_ vssd1 vssd1 vccd1 vccd1 _04353_ sky130_fd_sc_hd__o21a_1
XFILLER_0_117_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08239_ _03047_ _03375_ vssd1 vssd1 vccd1 vccd1 _03376_ sky130_fd_sc_hd__or2_1
XFILLER_0_144_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10327__S net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_179 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07008__A2 net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08205__A1 _03334_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11250_ net878 _05118_ _05130_ vssd1 vssd1 vccd1 vccd1 _05143_ sky130_fd_sc_hd__and3_1
XFILLER_0_132_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout888_X net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10201_ net258 net1937 net394 vssd1 vssd1 vccd1 vccd1 _00381_ sky130_fd_sc_hd__mux2_1
X_11181_ _05022_ _05034_ net473 net587 net1168 vssd1 vssd1 vccd1 vccd1 _01239_ sky130_fd_sc_hd__a32o_1
XANTENNA__07964__B1 net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10132_ net185 net1866 net609 vssd1 vssd1 vccd1 vccd1 _00332_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_54_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10062__S net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10063_ net1499 net225 net616 vssd1 vssd1 vccd1 vccd1 _00265_ sky130_fd_sc_hd__mux2_1
XANTENNA_input27_A DAT_I[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_187_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13822_ net1106 vssd1 vssd1 vccd1 vccd1 gpio_out[17] sky130_fd_sc_hd__buf_2
XFILLER_0_15_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13753_ clknet_leaf_99_clk _01324_ vssd1 vssd1 vccd1 vccd1 top.lcd.cnt_20ms\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__11276__B1 _05150_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10965_ top.a1.dataInTemp\[1\] net785 vssd1 vssd1 vccd1 vccd1 _05007_ sky130_fd_sc_hd__or2_1
XANTENNA__12536__CLK clknet_leaf_128_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12704_ clknet_leaf_113_clk _00296_ net991 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[6\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_183_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13684_ clknet_leaf_92_clk _01260_ net999 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07495__A2 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08991__A _03653_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10896_ net1422 net238 net479 vssd1 vssd1 vccd1 vccd1 _01057_ sky130_fd_sc_hd__mux2_1
XANTENNA__11291__A3 _05128_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_182_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_174_3059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12635_ clknet_leaf_120_clk _00227_ net930 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[4\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_799 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12566_ clknet_leaf_12_clk _00158_ net942 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[2\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_124_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_156_2781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_156_2792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11517_ _05380_ _05396_ vssd1 vssd1 vccd1 vccd1 _05400_ sky130_fd_sc_hd__nor2_1
XFILLER_0_163_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10237__S net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12497_ clknet_leaf_93_clk _00089_ net994 vssd1 vssd1 vccd1 vccd1 top.pc\[9\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_151_652 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold209 top.DUT.register\[13\]\[18\] vssd1 vssd1 vccd1 vccd1 net1325 sky130_fd_sc_hd__dlygate4sd3_1
X_11448_ _05329_ _05330_ vssd1 vssd1 vccd1 vccd1 _05331_ sky130_fd_sc_hd__nand2_1
XFILLER_0_151_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_189_3280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11379_ _05228_ _05229_ _05249_ _05250_ _05227_ vssd1 vssd1 vccd1 vccd1 _05262_ sky130_fd_sc_hd__a221o_1
X_13118_ clknet_leaf_18_clk _00710_ net1031 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[19\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_186_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13049_ clknet_leaf_13_clk _00641_ net943 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[17\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12593__RESET_B net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07707__B1 net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08380__B1 net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07610_ _02729_ _02748_ net825 vssd1 vssd1 vccd1 vccd1 _02749_ sky130_fd_sc_hd__mux2_2
X_08590_ _03270_ _03274_ vssd1 vssd1 vccd1 vccd1 _03714_ sky130_fd_sc_hd__nand2_1
XANTENNA__10700__S net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_205_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_3_4_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_3_4_0_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_85_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09062__A _03561_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11267__B1 _05150_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07541_ _02359_ _02679_ vssd1 vssd1 vccd1 vccd1 _02680_ sky130_fd_sc_hd__or2_1
XFILLER_0_48_216 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07486__A2 net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07472_ _02590_ _02610_ vssd1 vssd1 vccd1 vccd1 _02611_ sky130_fd_sc_hd__nand2_1
XFILLER_0_159_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_201_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09211_ _01505_ _04280_ vssd1 vssd1 vccd1 vccd1 _04281_ sky130_fd_sc_hd__nand2_1
X_06423_ net684 _01516_ _01523_ vssd1 vssd1 vccd1 vccd1 _01562_ sky130_fd_sc_hd__and3_4
XANTENNA__11019__B1 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09142_ _02858_ _02899_ vssd1 vssd1 vccd1 vccd1 _04216_ sky130_fd_sc_hd__or2_2
X_06354_ _01490_ _01493_ vssd1 vssd1 vccd1 vccd1 _01494_ sky130_fd_sc_hd__nor2_1
XANTENNA__07238__A2 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_20_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09073_ _01479_ _02334_ _02344_ _04145_ _04147_ vssd1 vssd1 vccd1 vccd1 _04148_ sky130_fd_sc_hd__o311a_1
XFILLER_0_72_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10147__S net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06285_ top.lcd.nextState\[4\] net815 net813 top.lcd.currentState\[4\] net1084 vssd1
+ vssd1 vccd1 vccd1 _01333_ sky130_fd_sc_hd__o221a_2
XANTENNA_fanout214_A _04771_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08024_ _03162_ vssd1 vssd1 vccd1 vccd1 _03163_ sky130_fd_sc_hd__inv_2
XFILLER_0_141_151 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold710 top.DUT.register\[10\]\[5\] vssd1 vssd1 vccd1 vccd1 net1826 sky130_fd_sc_hd__dlygate4sd3_1
Xhold721 top.DUT.register\[28\]\[28\] vssd1 vssd1 vccd1 vccd1 net1837 sky130_fd_sc_hd__dlygate4sd3_1
Xhold732 top.DUT.register\[18\]\[26\] vssd1 vssd1 vccd1 vccd1 net1848 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08199__B1 net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_1883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold743 top.DUT.register\[17\]\[13\] vssd1 vssd1 vccd1 vccd1 net1859 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold754 top.DUT.register\[23\]\[3\] vssd1 vssd1 vccd1 vccd1 net1870 sky130_fd_sc_hd__dlygate4sd3_1
Xhold765 top.DUT.register\[20\]\[6\] vssd1 vssd1 vccd1 vccd1 net1881 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold776 top.DUT.register\[31\]\[31\] vssd1 vssd1 vccd1 vccd1 net1892 sky130_fd_sc_hd__dlygate4sd3_1
Xhold787 top.DUT.register\[5\]\[18\] vssd1 vssd1 vccd1 vccd1 net1903 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09237__A _02544_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07410__A2 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09975_ net1536 net148 net629 vssd1 vssd1 vccd1 vccd1 _00183_ sky130_fd_sc_hd__mux2_1
Xhold798 top.DUT.register\[24\]\[30\] vssd1 vssd1 vccd1 vccd1 net1914 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout583_A _01513_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08926_ _03323_ _03345_ net277 vssd1 vssd1 vccd1 vccd1 _04034_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_99_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_207_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08857_ _03951_ _03968_ vssd1 vssd1 vccd1 vccd1 _03969_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout371_X net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout750_A _01621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout469_X net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07808_ _02945_ _02946_ vssd1 vssd1 vccd1 vccd1 _02947_ sky130_fd_sc_hd__nor2_2
XANTENNA__10610__S net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08788_ _01919_ net433 net501 _01918_ vssd1 vssd1 vccd1 vccd1 _03903_ sky130_fd_sc_hd__a22o_1
XFILLER_0_196_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11258__B1 _05150_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07739_ _02877_ vssd1 vssd1 vccd1 vccd1 _02878_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_0_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout636_X net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10750_ net1484 net181 net418 vssd1 vssd1 vccd1 vccd1 _00911_ sky130_fd_sc_hd__mux2_1
XANTENNA__07477__A2 net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06384__A_N top.a1.instruction\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09409_ _04447_ _04448_ _04449_ vssd1 vssd1 vccd1 vccd1 _04467_ sky130_fd_sc_hd__o21ai_1
XANTENNA__06685__B1 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10681_ net1758 net186 net341 vssd1 vssd1 vccd1 vccd1 _00844_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12420_ clknet_leaf_94_clk top.ru.next_read_i net994 vssd1 vssd1 vccd1 vccd1 top.Ren
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07229__A2 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_7__f_clk clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_7__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_90_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12351_ net2267 net120 _00016_ vssd1 vssd1 vccd1 vccd1 _01376_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10057__S net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11302_ top.a1.row1\[101\] _05189_ net815 vssd1 vssd1 vccd1 vccd1 _05190_ sky130_fd_sc_hd__a21o_1
X_12282_ top.lcd.cnt_500hz\[9\] top.lcd.cnt_500hz\[10\] _06097_ vssd1 vssd1 vccd1
+ vccd1 _06100_ sky130_fd_sc_hd__and3_1
XFILLER_0_133_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11233_ net880 top.lcd.nextState\[0\] _05123_ vssd1 vssd1 vccd1 vccd1 _05126_ sky130_fd_sc_hd__and3_1
XANTENNA__07401__A2 net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11164_ top.a1.row1\[58\] _05091_ _05085_ vssd1 vssd1 vccd1 vccd1 _01229_ sky130_fd_sc_hd__mux2_1
XANTENNA__08051__A _01678_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10115_ net263 net2160 net607 vssd1 vssd1 vccd1 vccd1 _00315_ sky130_fd_sc_hd__mux2_1
X_11095_ net69 net865 vssd1 vssd1 vccd1 vccd1 _05053_ sky130_fd_sc_hd__and2_1
X_10046_ net689 _04713_ _04952_ vssd1 vssd1 vccd1 vccd1 _04954_ sky130_fd_sc_hd__and3_4
XFILLER_0_117_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06777__Y _01916_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold70 top.a1.data\[11\] vssd1 vssd1 vccd1 vccd1 net1186 sky130_fd_sc_hd__dlygate4sd3_1
Xhold81 top.ramstore\[27\] vssd1 vssd1 vccd1 vccd1 net1197 sky130_fd_sc_hd__dlygate4sd3_1
Xhold92 _01167_ vssd1 vssd1 vccd1 vccd1 net1208 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10520__S net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_187_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13805_ clknet_leaf_69_clk _01374_ net1097 vssd1 vssd1 vccd1 vccd1 top.pad.keyCode\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_11997_ _01402_ net126 _05852_ vssd1 vssd1 vccd1 vccd1 _05880_ sky130_fd_sc_hd__a21boi_1
XTAP_TAPCELL_ROW_67_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08973__A1_N _01697_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09311__C1 net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10948_ net1755 net157 net592 vssd1 vssd1 vccd1 vccd1 _01109_ sky130_fd_sc_hd__mux2_1
X_13736_ clknet_leaf_93_clk _01307_ vssd1 vssd1 vccd1 vccd1 top.a1.dataInTemp\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__07468__A2 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08665__B2 _03342_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_158_2810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_158_2821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09032__D _04064_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06676__B1 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13667_ clknet_leaf_90_clk _01243_ net999 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[120\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_80_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10879_ net178 net1676 net596 vssd1 vssd1 vccd1 vccd1 _01040_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_80_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12618_ clknet_leaf_121_clk _00210_ net933 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[3\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08417__A1 net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13598_ clknet_leaf_64_clk net1163 net1091 vssd1 vssd1 vccd1 vccd1 net90 sky130_fd_sc_hd__dfrtp_1
XANTENNA__08417__B2 _03548_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12549_ clknet_leaf_35_clk _00141_ net1041 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[1\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_170_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_436 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_1 _01501_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07640__A2 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07784__B _02922_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09057__A _03121_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout508 _01565_ vssd1 vssd1 vccd1 vccd1 net508 sky130_fd_sc_hd__clkbuf_4
Xfanout519 net522 vssd1 vssd1 vccd1 vccd1 net519 sky130_fd_sc_hd__buf_4
XFILLER_0_67_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06600__B1 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_169_2983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09760_ _04386_ _04776_ _04781_ _04754_ vssd1 vssd1 vccd1 vccd1 _04782_ sky130_fd_sc_hd__a211o_1
X_06972_ _02101_ _02110_ vssd1 vssd1 vccd1 vccd1 _02111_ sky130_fd_sc_hd__nor2_4
XTAP_TAPCELL_ROW_206_3534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08711_ net883 top.pc\[20\] net694 _03829_ vssd1 vssd1 vccd1 vccd1 _03830_ sky130_fd_sc_hd__a22o_1
X_09691_ _03353_ net404 net489 _04725_ vssd1 vssd1 vccd1 vccd1 _04726_ sky130_fd_sc_hd__o211a_4
Xfanout1090 net1091 vssd1 vssd1 vccd1 vccd1 net1090 sky130_fd_sc_hd__clkbuf_4
X_08642_ net496 _03748_ _03763_ net423 vssd1 vssd1 vccd1 vccd1 _03764_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__10430__S net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09504__B top.pc\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08573_ net430 _03696_ _03697_ net426 vssd1 vssd1 vccd1 vccd1 _03698_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_25_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07524_ top.DUT.register\[13\]\[7\] net463 net535 top.DUT.register\[19\]\[7\] _02662_
+ vssd1 vssd1 vccd1 vccd1 _02663_ sky130_fd_sc_hd__a221o_1
XANTENNA__08656__A1 net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07459__A2 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09853__B1 _04151_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06667__B1 net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07455_ top.DUT.register\[24\]\[15\] net643 net743 top.DUT.register\[2\]\[15\] _02593_
+ vssd1 vssd1 vccd1 vccd1 _02594_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout331_A net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout429_A net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1073_A net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06406_ _01520_ _01530_ _01538_ _01544_ vssd1 vssd1 vccd1 vccd1 _01545_ sky130_fd_sc_hd__or4_1
XANTENNA__08408__A1 _02678_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07386_ _02523_ _02524_ vssd1 vssd1 vccd1 vccd1 _02525_ sky130_fd_sc_hd__nand2b_2
XANTENNA__08136__A _02633_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_1912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_1923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_hold1181_A top.ramload\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09125_ _04174_ _04175_ _04142_ vssd1 vssd1 vccd1 vccd1 _04200_ sky130_fd_sc_hd__mux2_1
XFILLER_0_162_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06337_ top.ru.state\[4\] net1733 net887 vssd1 vssd1 vccd1 vccd1 top.ru.next_dready
+ sky130_fd_sc_hd__o21ba_1
XANTENNA__08959__A2 net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_161_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09056_ _03846_ _03945_ _04003_ _03963_ vssd1 vssd1 vccd1 vccd1 _04131_ sky130_fd_sc_hd__or4b_1
XANTENNA__07092__B1 net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_170_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06268_ top.ramload\[29\] net854 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedData\[29\]
+ sky130_fd_sc_hd__and2_1
XANTENNA__07631__A2 net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08007_ top.a1.instruction\[28\] top.a1.instruction\[29\] top.a1.instruction\[30\]
+ top.a1.instruction\[31\] vssd1 vssd1 vccd1 vccd1 _03146_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout798_A _04150_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09908__A1 _03987_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold540 top.DUT.register\[25\]\[18\] vssd1 vssd1 vccd1 vccd1 net1656 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10605__S net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06199_ top.Wen top.Ren vssd1 vssd1 vccd1 vccd1 _01430_ sky130_fd_sc_hd__xnor2_1
Xhold551 top.DUT.register\[30\]\[5\] vssd1 vssd1 vccd1 vccd1 net1667 sky130_fd_sc_hd__dlygate4sd3_1
Xhold562 top.DUT.register\[17\]\[20\] vssd1 vssd1 vccd1 vccd1 net1678 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_491 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_3_3_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold573 top.DUT.register\[1\]\[13\] vssd1 vssd1 vccd1 vccd1 net1689 sky130_fd_sc_hd__dlygate4sd3_1
Xhold584 top.DUT.register\[11\]\[28\] vssd1 vssd1 vccd1 vccd1 net1700 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold595 top.DUT.register\[30\]\[25\] vssd1 vssd1 vccd1 vccd1 net1711 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12444__RESET_B net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout586_X net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout965_A net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_15__f_clk clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_15__leaf_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__11191__A2 net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09958_ net1619 net207 net629 vssd1 vssd1 vccd1 vccd1 _00166_ sky130_fd_sc_hd__mux2_1
X_08909_ net277 _03189_ _03197_ _04017_ net306 vssd1 vssd1 vccd1 vccd1 _04018_ sky130_fd_sc_hd__a311o_1
XANTENNA_fanout753_X net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09889_ top.pc\[27\] _04590_ vssd1 vssd1 vccd1 vccd1 _04898_ sky130_fd_sc_hd__and2_1
XFILLER_0_99_436 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11920_ _05791_ _05802_ vssd1 vssd1 vccd1 vccd1 _05803_ sky130_fd_sc_hd__and2_1
XANTENNA__10340__S net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09414__B _04471_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07698__A2 net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11851_ _05730_ _05731_ _05733_ vssd1 vssd1 vccd1 vccd1 _05734_ sky130_fd_sc_hd__a21o_1
X_10802_ net227 net2310 net598 vssd1 vssd1 vccd1 vccd1 _00963_ sky130_fd_sc_hd__mux2_1
XFILLER_0_184_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11782_ top.a1.dataIn\[7\] _05662_ _05663_ vssd1 vssd1 vccd1 vccd1 _05665_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_49_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09844__B1 net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06658__B1 net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10733_ net1564 net251 net418 vssd1 vssd1 vccd1 vccd1 _00894_ sky130_fd_sc_hd__mux2_1
X_13521_ clknet_leaf_72_clk _01113_ net1080 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[101\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_171_3007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_171_3018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13452_ clknet_leaf_65_clk _01044_ net1095 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[29\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10664_ net2145 net263 net338 vssd1 vssd1 vccd1 vccd1 _00827_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_62_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07870__A2 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_180_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12403_ clknet_leaf_105_clk top.ru.next_FetchedInstr\[15\] net973 vssd1 vssd1 vccd1
+ vccd1 top.a1.instruction\[15\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_63_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_153_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13383_ clknet_leaf_7_clk _00975_ net944 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[27\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_153_2740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10595_ _04713_ _04952_ net400 vssd1 vssd1 vccd1 vccd1 _04991_ sky130_fd_sc_hd__nand3_4
X_12334_ net1231 _06131_ _06132_ vssd1 vssd1 vccd1 vccd1 _01364_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07622__A2 net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06830__B1 net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12265_ _01437_ net686 _06089_ vssd1 vssd1 vccd1 vccd1 _01338_ sky130_fd_sc_hd__and3_1
XFILLER_0_121_655 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10515__S net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_128_Right_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11216_ net845 _05101_ vssd1 vssd1 vccd1 vccd1 _05114_ sky130_fd_sc_hd__and2_1
X_12196_ net1370 _06042_ net688 vssd1 vssd1 vccd1 vccd1 _01303_ sky130_fd_sc_hd__mux2_1
Xoutput60 net60 vssd1 vssd1 vccd1 vccd1 ADR_O[28] sky130_fd_sc_hd__buf_2
Xoutput71 net71 vssd1 vssd1 vccd1 vccd1 ADR_O[9] sky130_fd_sc_hd__buf_2
Xoutput82 net82 vssd1 vssd1 vccd1 vccd1 DAT_O[18] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_128_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput93 net93 vssd1 vssd1 vccd1 vccd1 DAT_O[28] sky130_fd_sc_hd__clkbuf_4
X_11147_ _02952_ _02984_ _02993_ _04191_ vssd1 vssd1 vccd1 vccd1 _05079_ sky130_fd_sc_hd__o31a_1
XFILLER_0_207_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_182_3169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11078_ net94 net872 net836 net1147 vssd1 vssd1 vccd1 vccd1 _01189_ sky130_fd_sc_hd__a22o_1
XFILLER_0_37_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09532__C1 _01393_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10250__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10029_ net2111 net190 net620 vssd1 vssd1 vccd1 vccd1 _00232_ sky130_fd_sc_hd__mux2_1
XANTENNA__07125__A _02242_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06897__B1 net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_201_3464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11870__A top.a1.dataIn\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09835__B1 net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13719_ clknet_leaf_98_clk _01290_ net986 vssd1 vssd1 vccd1 vccd1 top.a1.row2\[33\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_388 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07240_ top.DUT.register\[16\]\[10\] net734 _02366_ _02378_ vssd1 vssd1 vccd1 vccd1
+ _02379_ sky130_fd_sc_hd__a211o_1
XFILLER_0_5_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07171_ _02308_ _02309_ vssd1 vssd1 vccd1 vccd1 _02310_ sky130_fd_sc_hd__nor2_2
XFILLER_0_27_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07074__B1 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_169_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10425__S net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_1842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08403__B net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout305 net306 vssd1 vssd1 vccd1 vccd1 net305 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_1_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout316 _02880_ vssd1 vssd1 vccd1 vccd1 net316 sky130_fd_sc_hd__clkbuf_4
Xfanout327 net328 vssd1 vssd1 vccd1 vccd1 net327 sky130_fd_sc_hd__buf_2
X_09812_ _02679_ net486 net401 top.a1.dataIn\[19\] net397 vssd1 vssd1 vccd1 vccd1
+ _04829_ sky130_fd_sc_hd__a221o_1
Xfanout338 _04993_ vssd1 vssd1 vccd1 vccd1 net338 sky130_fd_sc_hd__buf_6
Xfanout349 _04991_ vssd1 vssd1 vccd1 vccd1 net349 sky130_fd_sc_hd__clkbuf_4
X_09743_ top.pc\[12\] _04172_ _04352_ vssd1 vssd1 vccd1 vccd1 _04767_ sky130_fd_sc_hd__and3_1
X_06955_ top.DUT.register\[26\]\[23\] net528 net453 top.DUT.register\[29\]\[23\] _02093_
+ vssd1 vssd1 vccd1 vccd1 _02094_ sky130_fd_sc_hd__a221o_1
XFILLER_0_94_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_207_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout379_A net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_19_Left_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09674_ top.a1.instruction\[11\] net786 vssd1 vssd1 vccd1 vccd1 _04710_ sky130_fd_sc_hd__nand2_1
XANTENNA__10160__S net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_2049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06886_ _02020_ _02022_ _02024_ vssd1 vssd1 vccd1 vccd1 _02025_ sky130_fd_sc_hd__or3_2
X_08625_ _02266_ _03727_ _02263_ vssd1 vssd1 vccd1 vccd1 _03747_ sky130_fd_sc_hd__o21ba_1
XANTENNA__06888__B1 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_806 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11780__A top.a1.dataIn\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08556_ net423 _03666_ _03669_ _03681_ vssd1 vssd1 vccd1 vccd1 _03682_ sky130_fd_sc_hd__a211o_1
XANTENNA__08565__S net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11228__A3 _05120_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_2249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07507_ top.DUT.register\[7\]\[14\] net660 _02635_ _02645_ vssd1 vssd1 vccd1 vccd1
+ _02646_ sky130_fd_sc_hd__a211o_1
XFILLER_0_182_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08487_ _03614_ _03615_ vssd1 vssd1 vccd1 vccd1 _03616_ sky130_fd_sc_hd__nor2_1
XANTENNA__07689__B _02827_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout334_X net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout713_A _01638_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_463 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_174_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07438_ top.DUT.register\[17\]\[15\] net460 net448 top.DUT.register\[21\]\[15\] _02576_
+ vssd1 vssd1 vccd1 vccd1 _02577_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_102_1971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_1982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07852__A2 net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout501_X net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_28_Left_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07369_ top.DUT.register\[10\]\[8\] net770 net707 top.DUT.register\[15\]\[8\] vssd1
+ vssd1 vccd1 vccd1 _02508_ sky130_fd_sc_hd__a22o_1
XFILLER_0_33_734 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09108_ _04176_ _04182_ vssd1 vssd1 vccd1 vccd1 _04183_ sky130_fd_sc_hd__and2_1
XFILLER_0_60_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07065__B1 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07604__A2 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_2470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10380_ net1486 net203 net375 vssd1 vssd1 vccd1 vccd1 _00555_ sky130_fd_sc_hd__mux2_1
XANTENNA__12625__RESET_B net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06812__B1 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09039_ _02947_ _04113_ _03413_ _01659_ vssd1 vssd1 vccd1 vccd1 _04114_ sky130_fd_sc_hd__or4b_1
XANTENNA__10335__S net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11149__C1 net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12050_ _05909_ _05918_ vssd1 vssd1 vccd1 vccd1 _05933_ sky130_fd_sc_hd__nand2_1
Xhold370 top.DUT.register\[14\]\[18\] vssd1 vssd1 vccd1 vccd1 net1486 sky130_fd_sc_hd__dlygate4sd3_1
Xhold381 top.DUT.register\[17\]\[19\] vssd1 vssd1 vccd1 vccd1 net1497 sky130_fd_sc_hd__dlygate4sd3_1
Xhold392 top.DUT.register\[17\]\[7\] vssd1 vssd1 vccd1 vccd1 net1508 sky130_fd_sc_hd__dlygate4sd3_1
X_11001_ net843 _05033_ _05034_ net849 top.a1.dataIn\[9\] vssd1 vssd1 vccd1 vccd1
+ _05035_ sky130_fd_sc_hd__a32o_1
Xfanout850 net851 vssd1 vssd1 vccd1 vccd1 net850 sky130_fd_sc_hd__clkbuf_2
Xfanout861 net863 vssd1 vssd1 vccd1 vccd1 net861 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_205_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout872 _01427_ vssd1 vssd1 vccd1 vccd1 net872 sky130_fd_sc_hd__buf_2
XANTENNA__06401__X _01540_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout883 net885 vssd1 vssd1 vccd1 vccd1 net883 sky130_fd_sc_hd__buf_2
XANTENNA__06591__A2 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout894 net895 vssd1 vssd1 vccd1 vccd1 net894 sky130_fd_sc_hd__buf_2
XFILLER_0_189_419 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10070__S net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_204_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08868__A1 net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12952_ clknet_leaf_127_clk _00544_ net918 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[14\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08868__B2 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1070 top.DUT.register\[5\]\[10\] vssd1 vssd1 vccd1 vccd1 net2186 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1081 top.DUT.register\[9\]\[15\] vssd1 vssd1 vccd1 vccd1 net2197 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1092 top.DUT.register\[4\]\[29\] vssd1 vssd1 vccd1 vccd1 net2208 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06879__B1 net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11903_ _05779_ _05781_ _05782_ _05785_ vssd1 vssd1 vccd1 vccd1 _05786_ sky130_fd_sc_hd__a31oi_4
X_12883_ clknet_leaf_122_clk _00475_ net932 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[12\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07540__A1 top.a1.instruction\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11834_ _05687_ _05712_ _05684_ vssd1 vssd1 vccd1 vccd1 _05717_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_184_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09160__A net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11765_ _05600_ _05639_ _05647_ vssd1 vssd1 vccd1 vccd1 _05648_ sky130_fd_sc_hd__o21ai_2
XANTENNA__09293__A1 net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09293__B2 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10716_ net1367 net201 net336 vssd1 vssd1 vccd1 vccd1 _00877_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13504_ clknet_leaf_80_clk _01096_ net992 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[31\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_11696_ _05577_ _05578_ vssd1 vssd1 vccd1 vccd1 _05579_ sky130_fd_sc_hd__xor2_4
XANTENNA__07843__A2 net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_544 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13435_ clknet_leaf_125_clk _01027_ net924 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[29\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_130_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10647_ net203 top.DUT.register\[22\]\[18\] net344 vssd1 vssd1 vccd1 vccd1 _00811_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07056__B1 net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13366_ clknet_leaf_11_clk _00958_ net948 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[27\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12366__RESET_B net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10578_ net1439 net190 net351 vssd1 vssd1 vccd1 vccd1 _00744_ sky130_fd_sc_hd__mux2_1
XANTENNA__08504__A net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06803__B1 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12317_ top.pad.button_control.r_counter\[6\] _06120_ vssd1 vssd1 vccd1 vccd1 _06122_
+ sky130_fd_sc_hd__and2_1
XANTENNA__10245__S net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13297_ clknet_leaf_113_clk _00889_ net990 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[25\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09319__B _04370_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_197_Left_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_184_3209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12026__A top.a1.dataIn\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12248_ top.lcd.cnt_20ms\[14\] _06079_ vssd1 vssd1 vccd1 vccd1 _06080_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_75_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_166_2931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12179_ net1555 net847 net797 _05916_ vssd1 vssd1 vccd1 vccd1 _01287_ sky130_fd_sc_hd__a22o_1
XANTENNA__08020__A2 _03157_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_166_2942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08308__B1 _03437_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06740_ top.DUT.register\[19\]\[24\] net538 net520 top.DUT.register\[10\]\[24\] vssd1
+ vssd1 vccd1 vccd1 _01879_ sky130_fd_sc_hd__a22o_1
XFILLER_0_3_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_199_3430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09520__A2 _04543_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06671_ _01809_ vssd1 vssd1 vccd1 vccd1 _01810_ sky130_fd_sc_hd__inv_2
X_08410_ _03419_ _03541_ net313 vssd1 vssd1 vccd1 vccd1 _03542_ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09390_ top.pc\[18\] _04438_ vssd1 vssd1 vccd1 vccd1 _04449_ sky130_fd_sc_hd__or2_1
X_08341_ _03417_ _03474_ net288 vssd1 vssd1 vccd1 vccd1 _03475_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_35_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_87 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08272_ net303 _03407_ _03371_ vssd1 vssd1 vccd1 vccd1 _03408_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_15_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_72 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07223_ top.a1.instruction\[7\] _01474_ vssd1 vssd1 vccd1 vccd1 _02362_ sky130_fd_sc_hd__and2_1
XFILLER_0_116_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07047__B1 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07154_ top.DUT.register\[13\]\[11\] net774 _02291_ _02292_ vssd1 vssd1 vccd1 vccd1
+ _02293_ sky130_fd_sc_hd__a211o_1
XFILLER_0_125_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10155__S net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07085_ top.DUT.register\[16\]\[16\] net546 net504 top.DUT.register\[27\]\[16\] vssd1
+ vssd1 vccd1 vccd1 _02224_ sky130_fd_sc_hd__a22o_1
XFILLER_0_14_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1036_A net1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout496_A net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout135 _04210_ vssd1 vssd1 vccd1 vccd1 net135 sky130_fd_sc_hd__clkbuf_2
Xfanout146 net147 vssd1 vssd1 vccd1 vccd1 net146 sky130_fd_sc_hd__clkbuf_2
Xfanout157 net158 vssd1 vssd1 vccd1 vccd1 net157 sky130_fd_sc_hd__clkbuf_2
XANTENNA_input1_A ACK_I vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout168 net169 vssd1 vssd1 vccd1 vccd1 net168 sky130_fd_sc_hd__buf_2
XFILLER_0_199_706 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout179 _04868_ vssd1 vssd1 vccd1 vccd1 net179 sky130_fd_sc_hd__clkbuf_2
X_07987_ top.DUT.register\[7\]\[31\] net660 net732 top.DUT.register\[14\]\[31\] vssd1
+ vssd1 vccd1 vccd1 _03126_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout284_X net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout663_A _01605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06573__A2 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06938_ top.DUT.register\[4\]\[21\] net670 net761 top.DUT.register\[30\]\[21\] _02076_
+ vssd1 vssd1 vccd1 vccd1 _02077_ sky130_fd_sc_hd__a221o_1
XANTENNA__07036__Y _02175_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09726_ _04172_ net403 _04753_ vssd1 vssd1 vccd1 vccd1 _04754_ sky130_fd_sc_hd__a21boi_4
XFILLER_0_179_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06869_ top.DUT.register\[18\]\[18\] net549 net541 top.DUT.register\[8\]\[18\] vssd1
+ vssd1 vccd1 vccd1 _02008_ sky130_fd_sc_hd__a22o_1
X_09657_ _04679_ _04685_ _04690_ vssd1 vssd1 vccd1 vccd1 _04697_ sky130_fd_sc_hd__or3_1
XANTENNA_fanout451_X net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09899__B _04605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout830_A net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout549_X net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout928_A net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08608_ _03218_ _03241_ vssd1 vssd1 vccd1 vccd1 _03731_ sky130_fd_sc_hd__and2_1
X_09588_ _04633_ _04634_ vssd1 vssd1 vccd1 vccd1 _04635_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_38_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_139_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08539_ _02477_ _03641_ _03064_ vssd1 vssd1 vccd1 vccd1 _03665_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_210_787 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout716_X net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_182_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11550_ _05380_ _05392_ _05399_ vssd1 vssd1 vccd1 vccd1 _05433_ sky130_fd_sc_hd__o21a_1
XANTENNA__11082__A1 net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07286__B1 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10501_ net1951 net251 net357 vssd1 vssd1 vccd1 vccd1 _00670_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11481_ _05362_ _05363_ vssd1 vssd1 vccd1 vccd1 _05364_ sky130_fd_sc_hd__nor2_1
XFILLER_0_190_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13220_ clknet_leaf_37_clk _00812_ net1052 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[22\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10432_ net263 top.DUT.register\[16\]\[2\] net365 vssd1 vssd1 vccd1 vccd1 _00603_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07589__A1 top.a1.instruction\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13151_ clknet_leaf_19_clk _00743_ net1028 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[20\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10065__S net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10363_ net2086 net268 net375 vssd1 vssd1 vccd1 vccd1 _00538_ sky130_fd_sc_hd__mux2_1
X_12102_ _05973_ _05977_ _05984_ _05976_ vssd1 vssd1 vccd1 vccd1 _05985_ sky130_fd_sc_hd__o2bb2a_1
X_13082_ clknet_leaf_5_clk _00674_ net936 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[18\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_10294_ net1405 net140 net388 vssd1 vssd1 vccd1 vccd1 _00472_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13075__CLK clknet_leaf_120_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12033_ _05906_ _05908_ _05914_ _05915_ vssd1 vssd1 vccd1 vccd1 _05916_ sky130_fd_sc_hd__a31o_1
XANTENNA__06779__A _01897_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_148_2661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_8_clk_A clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_148_2672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06564__A2 net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout680 _01547_ vssd1 vssd1 vccd1 vccd1 net680 sky130_fd_sc_hd__buf_2
Xfanout691 net692 vssd1 vssd1 vccd1 vccd1 net691 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_70_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08994__A _03691_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11224__A_N top.lcd.nextState\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_161_2861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12935_ clknet_leaf_7_clk _00527_ net946 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[13\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_158_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12866_ clknet_leaf_9_clk _00458_ net947 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[11\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_815 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11817_ _01401_ net131 _05664_ vssd1 vssd1 vccd1 vccd1 _05700_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_200_264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_194_3360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12797_ clknet_leaf_13_clk _00389_ net919 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[9\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_32_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_141_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07277__B1 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11748_ _05618_ _05630_ vssd1 vssd1 vccd1 vccd1 _05631_ sky130_fd_sc_hd__nand2b_2
XANTENNA__07816__A2 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12547__RESET_B net1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11679_ _05522_ _05558_ vssd1 vssd1 vccd1 vccd1 _05562_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_71_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07029__B1 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13418_ clknet_leaf_118_clk _01010_ net957 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[28\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_180_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_180_Right_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_726 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13349_ clknet_leaf_35_clk _00941_ net1042 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[26\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_44 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08529__B1 _03655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07910_ _02880_ _02899_ _03048_ vssd1 vssd1 vccd1 vccd1 _03049_ sky130_fd_sc_hd__o21ba_1
X_08890_ _01701_ net493 vssd1 vssd1 vccd1 vccd1 _04000_ sky130_fd_sc_hd__nor2_1
XANTENNA__10703__S net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07841_ top.DUT.register\[23\]\[0\] net572 net555 top.DUT.register\[28\]\[0\] vssd1
+ vssd1 vccd1 vccd1 _02980_ sky130_fd_sc_hd__a22o_1
XANTENNA__09741__A2 net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06555__A2 net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07772_ top.DUT.register\[14\]\[2\] net730 net726 top.DUT.register\[18\]\[2\] vssd1
+ vssd1 vccd1 vccd1 _02911_ sky130_fd_sc_hd__a22o_1
X_06723_ top.DUT.register\[21\]\[25\] net655 _01858_ _01861_ vssd1 vssd1 vccd1 vccd1
+ _01862_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_104_2008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09511_ _04561_ _04562_ vssd1 vssd1 vccd1 vccd1 _04563_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_88_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_211_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09442_ _02156_ _04487_ _04490_ vssd1 vssd1 vccd1 vccd1 _04498_ sky130_fd_sc_hd__a21o_1
X_06654_ top.DUT.register\[8\]\[26\] net541 net525 top.DUT.register\[11\]\[26\] vssd1
+ vssd1 vccd1 vccd1 _01793_ sky130_fd_sc_hd__a22o_1
X_09373_ _04431_ _04432_ vssd1 vssd1 vccd1 vccd1 _04433_ sky130_fd_sc_hd__nand2_1
X_06585_ top.DUT.register\[6\]\[28\] net638 net712 top.DUT.register\[11\]\[28\] _01723_
+ vssd1 vssd1 vccd1 vccd1 _01724_ sky130_fd_sc_hd__a221o_1
XFILLER_0_46_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09257__A1 net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout244_A _04745_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09257__B2 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08324_ net428 _03443_ _03444_ _03263_ _03458_ vssd1 vssd1 vccd1 vccd1 _03459_ sky130_fd_sc_hd__a221o_1
XANTENNA__07268__B1 net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11064__B2 top.ramstore\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_522 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_191_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08255_ net885 top.pc\[2\] net696 _03391_ vssd1 vssd1 vccd1 vccd1 _03392_ sky130_fd_sc_hd__a22o_1
XFILLER_0_144_352 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08480__A2 net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout509_A net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07206_ net894 _01477_ vssd1 vssd1 vccd1 vccd1 _02345_ sky130_fd_sc_hd__nand2_1
XFILLER_0_131_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08186_ _03322_ _03323_ vssd1 vssd1 vccd1 vccd1 _03324_ sky130_fd_sc_hd__nand2_1
XANTENNA__08768__B1 net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_558 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07137_ _02269_ _02271_ _02273_ _02275_ vssd1 vssd1 vccd1 vccd1 _02276_ sky130_fd_sc_hd__or4_4
XANTENNA_fanout1039_X net1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07983__A net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07068_ top.DUT.register\[22\]\[22\] net648 net636 top.DUT.register\[6\]\[22\] _02206_
+ vssd1 vssd1 vccd1 vccd1 _02207_ sky130_fd_sc_hd__a221o_1
XANTENNA__07440__B1 net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout780_A _01603_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout878_A top.lcd.nextState\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06794__A2 net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout499_X net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10613__S net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09732__A2 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout666_X net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06546__A2 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06886__X _02025_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09709_ net407 _04739_ vssd1 vssd1 vccd1 vccd1 _04740_ sky130_fd_sc_hd__or2_1
X_10981_ net844 _05018_ _05019_ net849 top.a1.dataIn\[4\] vssd1 vssd1 vccd1 vccd1
+ _05020_ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout833_X net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_260 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12720_ clknet_leaf_28_clk _00312_ net1011 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[6\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_143_2591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07223__A top.a1.instruction\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12651_ clknet_leaf_50_clk _00243_ net1059 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[4\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_4_0__f_clk_X clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_308 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08038__B _02994_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11602_ _05464_ _05483_ _05484_ vssd1 vssd1 vccd1 vccd1 _05485_ sky130_fd_sc_hd__or3_1
XANTENNA__07259__B1 net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_176_3090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12582_ clknet_leaf_32_clk _00174_ net1044 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[2\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_194_296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_154_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11533_ _05396_ _05398_ top.a1.dataIn\[15\] vssd1 vssd1 vccd1 vccd1 _05416_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_108_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11464_ _05316_ _05343_ _05346_ vssd1 vssd1 vccd1 vccd1 _05347_ sky130_fd_sc_hd__nand3b_1
XANTENNA__08054__A _01572_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_536 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13203_ clknet_leaf_122_clk _00795_ net928 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[22\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_59_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10415_ net1310 net203 net370 vssd1 vssd1 vccd1 vccd1 _00587_ sky130_fd_sc_hd__mux2_1
X_11395_ _05246_ _05251_ vssd1 vssd1 vccd1 vccd1 _05278_ sky130_fd_sc_hd__nand2_1
XFILLER_0_150_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13134_ clknet_leaf_42_clk _00726_ net1064 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[19\]\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_10346_ net1552 net218 net379 vssd1 vssd1 vccd1 vccd1 _00522_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_72_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06785__A2 net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13065_ clknet_leaf_50_clk _00657_ net1061 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[17\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10523__S net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10277_ net1414 net196 net386 vssd1 vssd1 vccd1 vccd1 _00455_ sky130_fd_sc_hd__mux2_1
X_12016_ _05870_ _05889_ vssd1 vssd1 vccd1 vccd1 _05899_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_206_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06537__A2 net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09613__A top.a1.halfData\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12918_ clknet_leaf_12_clk _00510_ net942 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[13\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07498__B1 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_192_3319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12849_ clknet_leaf_116_clk _00441_ net957 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[11\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_186_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_291 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06370_ _01500_ net789 vssd1 vssd1 vccd1 vccd1 _01509_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_83_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08516__X _03643_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13240__CLK clknet_leaf_128_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08040_ _03178_ vssd1 vssd1 vccd1 vccd1 _03179_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_211_3614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_211_3625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07670__B1 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold903 top.DUT.register\[25\]\[29\] vssd1 vssd1 vccd1 vccd1 net2019 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold914 top.DUT.register\[2\]\[18\] vssd1 vssd1 vccd1 vccd1 net2030 sky130_fd_sc_hd__dlygate4sd3_1
Xhold925 top.DUT.register\[21\]\[12\] vssd1 vssd1 vccd1 vccd1 net2041 sky130_fd_sc_hd__dlygate4sd3_1
Xhold936 top.DUT.register\[16\]\[18\] vssd1 vssd1 vccd1 vccd1 net2052 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07422__B1 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold947 top.DUT.register\[3\]\[13\] vssd1 vssd1 vccd1 vccd1 net2063 sky130_fd_sc_hd__dlygate4sd3_1
Xhold958 top.DUT.register\[19\]\[10\] vssd1 vssd1 vccd1 vccd1 net2074 sky130_fd_sc_hd__dlygate4sd3_1
Xhold969 top.DUT.register\[21\]\[7\] vssd1 vssd1 vccd1 vccd1 net2085 sky130_fd_sc_hd__dlygate4sd3_1
X_09991_ net222 net1990 net623 vssd1 vssd1 vccd1 vccd1 _00196_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_11__f_clk_X clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08942_ net873 _03267_ vssd1 vssd1 vccd1 vccd1 _04049_ sky130_fd_sc_hd__nor2_4
XANTENNA__10433__S net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_2089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_209_3576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_209_3587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08873_ net284 net429 _03440_ _03983_ vssd1 vssd1 vccd1 vccd1 _03984_ sky130_fd_sc_hd__a31o_1
XANTENNA__06528__A2 net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout194_A _04850_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07824_ top.DUT.register\[29\]\[0\] net722 _02961_ _02962_ vssd1 vssd1 vccd1 vccd1
+ _02963_ sky130_fd_sc_hd__a211o_1
X_07755_ top.DUT.register\[18\]\[3\] net548 net520 top.DUT.register\[10\]\[3\] vssd1
+ vssd1 vccd1 vccd1 _02894_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout361_A net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout459_A net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11285__A1 top.a1.row1\[59\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06706_ top.DUT.register\[18\]\[25\] net550 net503 top.DUT.register\[27\]\[25\] vssd1
+ vssd1 vccd1 vccd1 _01845_ sky130_fd_sc_hd__a22o_1
XANTENNA__07314__Y _02453_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07489__B1 net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07686_ top.DUT.register\[8\]\[4\] net641 net705 top.DUT.register\[3\]\[4\] _02824_
+ vssd1 vssd1 vccd1 vccd1 _02825_ sky130_fd_sc_hd__a221o_1
XANTENNA__08139__A _02286_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_591 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06637_ top.DUT.register\[26\]\[27\] net753 net712 top.DUT.register\[11\]\[27\] vssd1
+ vssd1 vccd1 vccd1 _01776_ sky130_fd_sc_hd__a22o_1
X_09425_ _04465_ _04467_ _04464_ vssd1 vssd1 vccd1 vccd1 _04482_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_19_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_548 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06700__A2 net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06568_ top.DUT.register\[28\]\[28\] net557 net542 top.DUT.register\[8\]\[28\] vssd1
+ vssd1 vccd1 vccd1 _01707_ sky130_fd_sc_hd__a22o_1
XFILLER_0_164_436 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11037__B2 top.ramload\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09356_ _04414_ _04416_ vssd1 vssd1 vccd1 vccd1 _04417_ sky130_fd_sc_hd__nor2_1
XFILLER_0_81_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08307_ net303 net333 _03439_ vssd1 vssd1 vccd1 vccd1 _03442_ sky130_fd_sc_hd__and3_1
XFILLER_0_129_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09287_ net804 _02949_ _04335_ _04351_ vssd1 vssd1 vccd1 vccd1 _04352_ sky130_fd_sc_hd__o22a_2
X_06499_ net787 _01596_ _01600_ vssd1 vssd1 vccd1 vccd1 _01638_ sky130_fd_sc_hd__and3_4
XANTENNA__10608__S net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09650__A1 top.a1.halfData\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08238_ _02947_ _03046_ vssd1 vssd1 vccd1 vccd1 _03375_ sky130_fd_sc_hd__and2_1
XFILLER_0_160_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_160_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08169_ _01983_ net327 vssd1 vssd1 vccd1 vccd1 _03307_ sky130_fd_sc_hd__or2_1
XANTENNA__09402__A1 net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10200_ net259 net2137 net394 vssd1 vssd1 vccd1 vccd1 _00380_ sky130_fd_sc_hd__mux2_1
XANTENNA__07413__B1 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11180_ _05019_ _05030_ net473 net588 net1175 vssd1 vssd1 vccd1 vccd1 _01238_ sky130_fd_sc_hd__a32o_1
XFILLER_0_101_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10131_ net205 net1927 net610 vssd1 vssd1 vccd1 vccd1 _00331_ sky130_fd_sc_hd__mux2_1
XANTENNA__10343__S net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10062_ net1549 net189 net616 vssd1 vssd1 vccd1 vccd1 _00264_ sky130_fd_sc_hd__mux2_1
XANTENNA__09705__A2 net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_145_2620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13113__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13821_ net1105 vssd1 vssd1 vccd1 vccd1 gpio_out[16] sky130_fd_sc_hd__buf_2
XFILLER_0_199_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13752_ clknet_leaf_99_clk net1228 vssd1 vssd1 vccd1 vccd1 top.lcd.cnt_20ms\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_10964_ net1142 _05006_ net589 vssd1 vssd1 vccd1 vccd1 _01114_ sky130_fd_sc_hd__mux2_1
XANTENNA__09720__X _04749_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12703_ clknet_leaf_10_clk _00295_ net949 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[6\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_195_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13683_ clknet_leaf_92_clk _01259_ net997 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_183_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10895_ top.DUT.register\[30\]\[7\] net245 net478 vssd1 vssd1 vccd1 vccd1 _01056_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__13263__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_195_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_174_3049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12634_ clknet_leaf_5_clk _00226_ net936 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[4\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_170_406 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10518__S net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12565_ clknet_leaf_29_clk _00157_ net1019 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[2\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_170_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_156_2782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_156_2793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11516_ _05396_ _05398_ vssd1 vssd1 vccd1 vccd1 _05399_ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_478 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12496_ clknet_leaf_84_clk _00088_ net1000 vssd1 vssd1 vccd1 vccd1 top.pc\[8\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_151_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11447_ _05293_ _05326_ vssd1 vssd1 vccd1 vccd1 _05330_ sky130_fd_sc_hd__xor2_1
XFILLER_0_1_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_189_3281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11378_ _05249_ _05250_ _05227_ vssd1 vssd1 vccd1 vccd1 _05261_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07955__A1 _01810_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10329_ net2117 net147 net377 vssd1 vssd1 vccd1 vccd1 _00505_ sky130_fd_sc_hd__mux2_1
X_13117_ clknet_leaf_3_clk _00709_ net941 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[19\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10253__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13048_ clknet_leaf_128_clk _00640_ net921 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[17\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_179_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07183__A2 net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09343__A _02580_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06391__B1 net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07540_ top.a1.instruction\[27\] net789 net794 top.a1.instruction\[19\] vssd1 vssd1
+ vccd1 vccd1 _02679_ sky130_fd_sc_hd__a22o_2
XFILLER_0_72_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_80_clk_A clknet_4_6__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_504 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07471_ net823 _02609_ _01586_ vssd1 vssd1 vccd1 vccd1 _02610_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_174_712 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06422_ top.a1.instruction\[17\] top.a1.instruction\[18\] net685 _01523_ vssd1 vssd1
+ vccd1 vccd1 _01561_ sky130_fd_sc_hd__and4_4
X_09210_ _04261_ _04266_ _04278_ vssd1 vssd1 vccd1 vccd1 _04280_ sky130_fd_sc_hd__a21o_1
XANTENNA__12216__B1 net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_95_clk_A clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09141_ net132 _04213_ _04214_ vssd1 vssd1 vccd1 vccd1 _04215_ sky130_fd_sc_hd__nor3_1
X_06353_ top.pad.button_control.r_counter\[8\] _01492_ top.pad.button_control.r_counter\[10\]
+ top.pad.button_control.r_counter\[9\] vssd1 vssd1 vccd1 vccd1 _01493_ sky130_fd_sc_hd__o211a_1
XFILLER_0_72_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10428__S net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09072_ _03156_ _01488_ _02343_ vssd1 vssd1 vccd1 vccd1 _04147_ sky130_fd_sc_hd__or3b_1
XFILLER_0_32_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_20_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07643__B1 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06284_ top.lcd.nextState\[3\] net815 net813 top.lcd.currentState\[3\] net1084 vssd1
+ vssd1 vccd1 vccd1 _01332_ sky130_fd_sc_hd__o221a_2
XFILLER_0_4_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08023_ _02343_ _03155_ _01501_ vssd1 vssd1 vccd1 vccd1 _03162_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_141_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold700 top.DUT.register\[28\]\[4\] vssd1 vssd1 vccd1 vccd1 net1816 sky130_fd_sc_hd__dlygate4sd3_1
Xhold711 top.DUT.register\[21\]\[28\] vssd1 vssd1 vccd1 vccd1 net1827 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_112_2129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold722 top.DUT.register\[22\]\[30\] vssd1 vssd1 vccd1 vccd1 net1838 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_96_1884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold733 top.DUT.register\[3\]\[16\] vssd1 vssd1 vccd1 vccd1 net1849 sky130_fd_sc_hd__dlygate4sd3_1
Xhold744 top.DUT.register\[17\]\[12\] vssd1 vssd1 vccd1 vccd1 net1860 sky130_fd_sc_hd__dlygate4sd3_1
Xhold755 top.DUT.register\[1\]\[30\] vssd1 vssd1 vccd1 vccd1 net1871 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06749__A2 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold766 top.DUT.register\[13\]\[16\] vssd1 vssd1 vccd1 vccd1 net1882 sky130_fd_sc_hd__dlygate4sd3_1
Xhold777 top.DUT.register\[14\]\[26\] vssd1 vssd1 vccd1 vccd1 net1893 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10163__S net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold788 top.DUT.register\[2\]\[14\] vssd1 vssd1 vccd1 vccd1 net1904 sky130_fd_sc_hd__dlygate4sd3_1
X_09974_ net2077 net154 net630 vssd1 vssd1 vccd1 vccd1 _00182_ sky130_fd_sc_hd__mux2_1
Xhold799 top.ramaddr\[4\] vssd1 vssd1 vccd1 vccd1 net1915 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07038__A _02155_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_33_clk_A clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09952__S net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08925_ net497 _04032_ vssd1 vssd1 vccd1 vccd1 _04033_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout576_A net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08856_ _03962_ _03964_ _03967_ vssd1 vssd1 vccd1 vccd1 _03968_ sky130_fd_sc_hd__and3_2
XFILLER_0_207_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07174__A2 net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_2350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09253__A _02329_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07807_ _02925_ _02944_ vssd1 vssd1 vccd1 vccd1 _02946_ sky130_fd_sc_hd__nor2_2
X_08787_ net283 _03900_ _03901_ vssd1 vssd1 vccd1 vccd1 _03902_ sky130_fd_sc_hd__o21ba_1
XANTENNA_fanout364_X net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout743_A _01623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06921__A2 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13286__CLK clknet_leaf_40_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_48_clk_A clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07738_ _02868_ _02876_ vssd1 vssd1 vccd1 vccd1 _02877_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_0_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08123__A1 net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_140_2550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09540__X _04590_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout531_X net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout910_A net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11007__B net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07669_ top.a1.instruction\[25\] net806 _02807_ vssd1 vssd1 vccd1 vccd1 _02808_ sky130_fd_sc_hd__a21oi_4
XANTENNA_fanout629_X net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_177_594 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09408_ _04464_ _04465_ vssd1 vssd1 vccd1 vccd1 _04466_ sky130_fd_sc_hd__or2_1
XFILLER_0_137_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10680_ net1479 net206 net340 vssd1 vssd1 vccd1 vccd1 _00843_ sky130_fd_sc_hd__mux2_1
XFILLER_0_192_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09339_ _04389_ _04391_ _04387_ vssd1 vssd1 vccd1 vccd1 _04401_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_35_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10338__S net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_109_Right_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_106_clk_A clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12350_ net2259 net119 _00016_ vssd1 vssd1 vccd1 vccd1 _01375_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06988__A2 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11301_ top.lcd.nextState\[3\] net882 _05128_ _05179_ _05188_ vssd1 vssd1 vccd1 vccd1
+ _05189_ sky130_fd_sc_hd__a311o_1
X_12281_ top.lcd.cnt_500hz\[9\] _06097_ top.lcd.cnt_500hz\[10\] vssd1 vssd1 vccd1
+ vccd1 _06099_ sky130_fd_sc_hd__a21o_1
XFILLER_0_120_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11232_ net880 _01382_ _05123_ vssd1 vssd1 vccd1 vccd1 _05125_ sky130_fd_sc_hd__and3_1
XANTENNA__13091__RESET_B net1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11194__B1 _04668_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10073__S net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11163_ _01378_ _01418_ _05090_ vssd1 vssd1 vccd1 vccd1 _05091_ sky130_fd_sc_hd__o21a_1
XFILLER_0_101_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10114_ net269 net1810 net609 vssd1 vssd1 vccd1 vccd1 _00314_ sky130_fd_sc_hd__mux2_1
XANTENNA__09715__X _04745_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11094_ _01405_ net1537 net860 _05052_ vssd1 vssd1 vccd1 vccd1 _01198_ sky130_fd_sc_hd__a31o_1
XANTENNA__12503__CLK clknet_4_6__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10045_ net2246 net140 net620 vssd1 vssd1 vccd1 vccd1 _00248_ sky130_fd_sc_hd__mux2_1
XANTENNA__10801__S net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold60 top.ramstore\[1\] vssd1 vssd1 vccd1 vccd1 net1176 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08362__A1 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold71 net104 vssd1 vssd1 vccd1 vccd1 net1187 sky130_fd_sc_hd__dlygate4sd3_1
Xhold82 _01187_ vssd1 vssd1 vccd1 vccd1 net1198 sky130_fd_sc_hd__dlygate4sd3_1
Xhold93 net115 vssd1 vssd1 vccd1 vccd1 net1209 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06912__A2 net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13804_ clknet_leaf_69_clk _01373_ net1097 vssd1 vssd1 vccd1 vccd1 top.pad.keyCode\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_11996_ _05857_ _05878_ _05854_ vssd1 vssd1 vccd1 vccd1 _05879_ sky130_fd_sc_hd__a21o_1
XFILLER_0_187_358 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13735_ clknet_leaf_94_clk _01306_ vssd1 vssd1 vccd1 vccd1 top.a1.dataInTemp\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_10947_ net1781 net162 net592 vssd1 vssd1 vccd1 vccd1 _01108_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_158_2811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09862__A1 top.a1.instruction\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_158_2822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13666_ clknet_leaf_72_clk _01242_ net1081 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[111\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__07873__B1 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10878_ net180 net2127 net594 vssd1 vssd1 vccd1 vccd1 _01039_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_80_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12617_ clknet_leaf_50_clk _00209_ net1056 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[3\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10248__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08417__A2 top.pc\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13597_ clknet_leaf_65_clk net1131 net1094 vssd1 vssd1 vccd1 vccd1 net89 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_143_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07625__B1 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12548_ clknet_leaf_37_clk _00140_ net1051 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[1\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09090__A2 _01589_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06979__A2 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12479_ clknet_leaf_64_clk _00074_ net1092 vssd1 vssd1 vccd1 vccd1 top.ramstore\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_2 _01532_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11185__B1 _04668_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07928__A1 _02286_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09057__B _03264_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout509 net510 vssd1 vssd1 vccd1 vccd1 net509 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_158_68 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_169_2984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06971_ _02105_ _02107_ _02109_ vssd1 vssd1 vccd1 vccd1 _02110_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_206_3535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08710_ _02177_ net501 _03828_ vssd1 vssd1 vccd1 vccd1 _03829_ sky130_fd_sc_hd__a21bo_1
XANTENNA__10711__S net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09690_ top.a1.dataIn\[1\] _01489_ _04722_ top.pc\[1\] net407 vssd1 vssd1 vccd1 vccd1
+ _04725_ sky130_fd_sc_hd__a221o_1
XANTENNA__07156__A2 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1080 net1082 vssd1 vssd1 vccd1 vccd1 net1080 sky130_fd_sc_hd__clkbuf_4
Xfanout1091 net1093 vssd1 vssd1 vccd1 vccd1 net1091 sky130_fd_sc_hd__clkbuf_2
X_08641_ _01964_ _03761_ vssd1 vssd1 vccd1 vccd1 _03763_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_109_2080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06903__A2 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08572_ _03499_ _03533_ _03588_ _03695_ vssd1 vssd1 vccd1 vccd1 _03697_ sky130_fd_sc_hd__a211o_1
XFILLER_0_107_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_178_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_25_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07523_ top.DUT.register\[23\]\[7\] net571 net455 top.DUT.register\[25\]\[7\] vssd1
+ vssd1 vccd1 vccd1 _02662_ sky130_fd_sc_hd__a22o_1
XFILLER_0_190_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_122_2280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07454_ top.DUT.register\[21\]\[15\] net656 net652 top.DUT.register\[5\]\[15\] vssd1
+ vssd1 vccd1 vccd1 _02593_ sky130_fd_sc_hd__a22o_1
XFILLER_0_186_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07864__B1 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_190_99 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_174_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06405_ top.DUT.register\[16\]\[30\] net544 net542 top.DUT.register\[8\]\[30\] _01543_
+ vssd1 vssd1 vccd1 vccd1 _01544_ sky130_fd_sc_hd__a221o_1
XFILLER_0_91_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10158__S net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_82 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07385_ _02497_ _02522_ vssd1 vssd1 vccd1 vccd1 _02524_ sky130_fd_sc_hd__nand2_1
XFILLER_0_17_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout324_A net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_1913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09947__S net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06336_ _01481_ top.ru.state\[0\] vssd1 vssd1 vccd1 vccd1 top.ru.next_read_i sky130_fd_sc_hd__and2b_1
X_09124_ _04180_ _04181_ _04045_ vssd1 vssd1 vccd1 vccd1 _04199_ sky130_fd_sc_hd__mux2_1
XANTENNA__07616__B1 net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09055_ _03980_ _04021_ _03905_ _03921_ vssd1 vssd1 vccd1 vccd1 _04130_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_114_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06267_ top.ramload\[28\] net854 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedData\[28\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_32_459 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_483 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08006_ _03143_ _03144_ vssd1 vssd1 vccd1 vccd1 _03145_ sky130_fd_sc_hd__and2b_2
Xhold530 top.ramaddr\[7\] vssd1 vssd1 vccd1 vccd1 net1646 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09908__A2 net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06198_ net1 net860 vssd1 vssd1 vccd1 vccd1 _01429_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_38_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11176__B1 net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout693_A _04049_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold541 top.DUT.register\[5\]\[23\] vssd1 vssd1 vccd1 vccd1 net1657 sky130_fd_sc_hd__dlygate4sd3_1
Xhold552 top.DUT.register\[5\]\[5\] vssd1 vssd1 vccd1 vccd1 net1668 sky130_fd_sc_hd__dlygate4sd3_1
Xhold563 top.DUT.register\[5\]\[1\] vssd1 vssd1 vccd1 vccd1 net1679 sky130_fd_sc_hd__dlygate4sd3_1
Xhold574 top.DUT.register\[31\]\[12\] vssd1 vssd1 vccd1 vccd1 net1690 sky130_fd_sc_hd__dlygate4sd3_1
Xhold585 top.DUT.register\[26\]\[28\] vssd1 vssd1 vccd1 vccd1 net1701 sky130_fd_sc_hd__dlygate4sd3_1
Xhold596 top.DUT.register\[7\]\[25\] vssd1 vssd1 vccd1 vccd1 net1712 sky130_fd_sc_hd__dlygate4sd3_1
X_09957_ net2065 net212 net627 vssd1 vssd1 vccd1 vccd1 _00165_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout481_X net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout860_A _01428_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout958_A net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout579_X net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08908_ _03193_ net289 _03190_ vssd1 vssd1 vccd1 vccd1 _04017_ sky130_fd_sc_hd__and3b_1
XANTENNA__10621__S net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09888_ _04889_ _04890_ _04887_ vssd1 vssd1 vccd1 vccd1 _04897_ sky130_fd_sc_hd__a21o_1
XANTENNA__09541__B1 _04590_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08839_ _03930_ _03950_ vssd1 vssd1 vccd1 vccd1 _03952_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout746_X net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11850_ _05702_ _05719_ _05724_ _05732_ vssd1 vssd1 vccd1 vccd1 _05733_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_169_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10801_ net231 net1992 net598 vssd1 vssd1 vccd1 vccd1 _00962_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11781_ _05662_ _05663_ vssd1 vssd1 vccd1 vccd1 _05664_ sky130_fd_sc_hd__or2_1
XANTENNA__09844__A1 _03869_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13520_ clknet_leaf_31_clk _01112_ net1018 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[31\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_10732_ net1916 net258 net419 vssd1 vssd1 vccd1 vccd1 _00893_ sky130_fd_sc_hd__mux2_1
XFILLER_0_177_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_171_3008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_326 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13451_ clknet_leaf_50_clk _01043_ net1059 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[29\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_94_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10068__S net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_180_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_62_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10663_ net1730 net269 net340 vssd1 vssd1 vccd1 vccd1 _00826_ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_62_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_540 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12402_ clknet_leaf_103_clk top.ru.next_FetchedInstr\[14\] net976 vssd1 vssd1 vccd1
+ vccd1 top.a1.instruction\[14\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__07607__B1 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13382_ clknet_leaf_33_clk _00974_ net1044 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[27\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_10594_ net1750 net141 net351 vssd1 vssd1 vccd1 vccd1 _00760_ sky130_fd_sc_hd__mux2_1
XANTENNA__08614__X _03737_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_153_2741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12333_ top.pad.button_control.r_counter\[12\] _06131_ net791 vssd1 vssd1 vccd1 vccd1
+ _06132_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_180_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_3_3_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_3_3_0_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__09158__A _04216_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12264_ top.lcd.cnt_500hz\[1\] top.lcd.cnt_500hz\[0\] top.lcd.cnt_500hz\[2\] top.lcd.cnt_500hz\[3\]
+ vssd1 vssd1 vccd1 vccd1 _06089_ sky130_fd_sc_hd__a31o_1
XFILLER_0_10_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08062__A _01853_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_186_3240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11215_ _05113_ net1252 net472 vssd1 vssd1 vccd1 vccd1 _01258_ sky130_fd_sc_hd__mux2_1
XANTENNA__13451__CLK clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12195_ net1124 _06048_ net688 vssd1 vssd1 vccd1 vccd1 _01302_ sky130_fd_sc_hd__mux2_1
Xoutput50 net50 vssd1 vssd1 vccd1 vccd1 ADR_O[19] sky130_fd_sc_hd__buf_2
XFILLER_0_120_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08997__A _03556_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput61 net61 vssd1 vssd1 vccd1 vccd1 ADR_O[29] sky130_fd_sc_hd__buf_2
Xoutput72 net72 vssd1 vssd1 vccd1 vccd1 CYC_O sky130_fd_sc_hd__buf_2
Xoutput83 net83 vssd1 vssd1 vccd1 vccd1 DAT_O[19] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_101_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11146_ _01332_ _01469_ _05078_ _01448_ vssd1 vssd1 vccd1 vccd1 _01224_ sky130_fd_sc_hd__o211a_1
Xoutput94 net94 vssd1 vssd1 vccd1 vccd1 DAT_O[29] sky130_fd_sc_hd__clkbuf_4
XANTENNA__10390__A1 _04916_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_207_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11077_ net93 net872 net836 net1235 vssd1 vssd1 vccd1 vccd1 _01188_ sky130_fd_sc_hd__a22o_1
XANTENNA__10531__S net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07138__A2 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10028_ net1395 net197 net620 vssd1 vssd1 vccd1 vccd1 _00231_ sky130_fd_sc_hd__mux2_1
XFILLER_0_144_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_201_3454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_201_3465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_829 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11979_ top.a1.dataIn\[4\] _05852_ vssd1 vssd1 vccd1 vccd1 _05862_ sky130_fd_sc_hd__nor2_1
XANTENNA__09835__A1 _03848_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13718_ clknet_leaf_97_clk _01289_ net984 vssd1 vssd1 vccd1 vccd1 top.a1.row2\[32\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07846__B1 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_570 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07310__A2 net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_186 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13649_ clknet_leaf_89_clk _01228_ net1003 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[57\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_211_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09767__S net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07170_ _02286_ _02306_ vssd1 vssd1 vccd1 vccd1 _02309_ sky130_fd_sc_hd__nor2_1
XFILLER_0_81_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_30_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10706__S net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_120_clk clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_120_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_152_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08810__A2 net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_10_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_93_1843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12490__Q top.pc\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08023__B1 _01501_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout306 net307 vssd1 vssd1 vccd1 vccd1 net306 sky130_fd_sc_hd__buf_2
XANTENNA__07377__A2 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout317 net318 vssd1 vssd1 vccd1 vccd1 net317 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09771__B1 _04752_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09811_ _04824_ _04827_ vssd1 vssd1 vccd1 vccd1 _04828_ sky130_fd_sc_hd__xnor2_1
Xfanout328 net329 vssd1 vssd1 vccd1 vccd1 net328 sky130_fd_sc_hd__clkbuf_2
Xfanout339 _04993_ vssd1 vssd1 vccd1 vccd1 net339 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06585__B1 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload11_A clknet_leaf_128_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_185_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09742_ net1574 net222 net631 vssd1 vssd1 vccd1 vccd1 _00132_ sky130_fd_sc_hd__mux2_1
XANTENNA__10441__S net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06954_ top.DUT.register\[23\]\[23\] net572 net568 top.DUT.register\[6\]\[23\] vssd1
+ vssd1 vccd1 vccd1 _02093_ sky130_fd_sc_hd__a22o_1
XANTENNA__07129__A2 net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09673_ top.a1.instruction\[11\] net786 vssd1 vssd1 vccd1 vccd1 _04709_ sky130_fd_sc_hd__and2_1
X_06885_ top.DUT.register\[10\]\[18\] net520 net453 top.DUT.register\[29\]\[18\] _02023_
+ vssd1 vssd1 vccd1 vccd1 _02024_ sky130_fd_sc_hd__a221o_1
X_08624_ net1611 net833 net803 _03746_ vssd1 vssd1 vccd1 vccd1 _00034_ sky130_fd_sc_hd__a22o_1
XFILLER_0_96_407 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08555_ _02433_ net499 net494 _02434_ _03680_ vssd1 vssd1 vccd1 vccd1 _03681_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_120_2239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout441_A _01566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_204_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout539_A _01540_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_367 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07506_ top.DUT.register\[9\]\[14\] net763 net732 top.DUT.register\[14\]\[14\] _02634_
+ vssd1 vssd1 vccd1 vccd1 _02645_ sky130_fd_sc_hd__a221o_1
XFILLER_0_147_520 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07837__B1 net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08147__A _02899_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_194_Right_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08486_ _02389_ _03613_ vssd1 vssd1 vccd1 vccd1 _03615_ sky130_fd_sc_hd__nor2_1
XANTENNA__10396__B _04155_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07301__A2 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07437_ top.DUT.register\[8\]\[15\] net540 net531 top.DUT.register\[12\]\[15\] vssd1
+ vssd1 vccd1 vccd1 _02576_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_102_1972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_475 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout706_A _01640_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_1983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12189__A2 net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07368_ top.DUT.register\[26\]\[8\] net751 net711 top.DUT.register\[11\]\[8\] vssd1
+ vssd1 vccd1 vccd1 _02507_ sky130_fd_sc_hd__a22o_1
XFILLER_0_18_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_746 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09107_ _04181_ _04180_ _04045_ vssd1 vssd1 vccd1 vccd1 _04182_ sky130_fd_sc_hd__mux2_1
X_06319_ top.pad.count\[0\] top.pad.count\[1\] vssd1 vssd1 vccd1 vccd1 net117 sky130_fd_sc_hd__nor2_1
XFILLER_0_162_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10616__S net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07299_ top.DUT.register\[22\]\[12\] net575 net507 top.DUT.register\[4\]\[12\] _02437_
+ vssd1 vssd1 vccd1 vccd1 _02438_ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_111_clk clknet_4_6__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_111_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_103_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_135_2471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09038_ _01877_ _02803_ _02852_ vssd1 vssd1 vccd1 vccd1 _04113_ sky130_fd_sc_hd__nand3_1
XFILLER_0_60_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout696_X net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08972__A1_N _01741_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold360 top.ramaddr\[0\] vssd1 vssd1 vccd1 vccd1 net1476 sky130_fd_sc_hd__dlygate4sd3_1
Xhold371 top.DUT.register\[13\]\[15\] vssd1 vssd1 vccd1 vccd1 net1487 sky130_fd_sc_hd__dlygate4sd3_1
Xhold382 top.DUT.register\[6\]\[11\] vssd1 vssd1 vccd1 vccd1 net1498 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07368__A2 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11000_ top.a1.data\[5\] net783 vssd1 vssd1 vccd1 vccd1 _05034_ sky130_fd_sc_hd__or2_1
Xhold393 top.DUT.register\[23\]\[15\] vssd1 vssd1 vccd1 vccd1 net1509 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06576__B1 net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10372__A1 net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout863_X net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout840 _05042_ vssd1 vssd1 vccd1 vccd1 net840 sky130_fd_sc_hd__clkbuf_2
Xfanout851 _04662_ vssd1 vssd1 vccd1 vccd1 net851 sky130_fd_sc_hd__clkbuf_2
XANTENNA__10351__S net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout862 net863 vssd1 vssd1 vccd1 vccd1 net862 sky130_fd_sc_hd__clkbuf_2
Xfanout873 net877 vssd1 vssd1 vccd1 vccd1 net873 sky130_fd_sc_hd__buf_4
Xfanout884 net885 vssd1 vssd1 vccd1 vccd1 net884 sky130_fd_sc_hd__clkbuf_2
Xfanout895 top.a1.instruction\[12\] vssd1 vssd1 vccd1 vccd1 net895 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_99_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12951_ clknet_leaf_129_clk _00543_ net911 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[14\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09144__C _04217_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1060 top.DUT.register\[21\]\[22\] vssd1 vssd1 vccd1 vccd1 net2176 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1071 top.DUT.register\[29\]\[7\] vssd1 vssd1 vccd1 vccd1 net2187 sky130_fd_sc_hd__dlygate4sd3_1
X_11902_ _05760_ _05766_ vssd1 vssd1 vccd1 vccd1 _05785_ sky130_fd_sc_hd__nand2b_1
Xhold1082 top.DUT.register\[22\]\[26\] vssd1 vssd1 vccd1 vccd1 net2198 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1093 top.DUT.register\[10\]\[16\] vssd1 vssd1 vccd1 vccd1 net2209 sky130_fd_sc_hd__dlygate4sd3_1
X_12882_ clknet_leaf_23_clk _00474_ net1021 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[12\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07540__A2 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_464 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11833_ _05705_ _05710_ _05711_ _05713_ _05715_ vssd1 vssd1 vccd1 vccd1 _05716_ sky130_fd_sc_hd__o311ai_4
XTAP_TAPCELL_ROW_64_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11764_ _05597_ _05599_ _05620_ _05598_ vssd1 vssd1 vccd1 vccd1 _05647_ sky130_fd_sc_hd__a31o_1
XFILLER_0_95_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_161_Right_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13503_ clknet_leaf_19_clk _01095_ net1026 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[31\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_10715_ net1565 net184 net335 vssd1 vssd1 vccd1 vccd1 _00876_ sky130_fd_sc_hd__mux2_1
XANTENNA__06500__B1 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11695_ _05537_ _05541_ _05570_ vssd1 vssd1 vccd1 vccd1 _05578_ sky130_fd_sc_hd__and3_1
XFILLER_0_193_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13434_ clknet_leaf_1_clk _01026_ net916 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[29\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_10646_ net218 net1918 net342 vssd1 vssd1 vccd1 vccd1 _00810_ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08253__B1 _03363_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13365_ clknet_leaf_30_clk _00957_ net1019 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[27\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_102_clk clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_102_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__10526__S net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10577_ net1856 net198 net351 vssd1 vssd1 vccd1 vccd1 _00743_ sky130_fd_sc_hd__mux2_1
X_12316_ _06120_ _06121_ vssd1 vssd1 vccd1 vccd1 _01357_ sky130_fd_sc_hd__nor2_1
XFILLER_0_2_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13296_ clknet_leaf_28_clk _00888_ net1018 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[24\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12026__B _05879_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12247_ _06079_ net978 _06078_ vssd1 vssd1 vccd1 vccd1 _01324_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_75_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08556__A1 net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07835__S net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_166_2932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12178_ net1258 net848 net796 _05937_ vssd1 vssd1 vccd1 vccd1 _01286_ sky130_fd_sc_hd__a22o_1
XANTENNA__06567__B1 net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_166_2943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09335__B _04386_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10261__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11129_ net56 net869 vssd1 vssd1 vccd1 vccd1 _05070_ sky130_fd_sc_hd__and2_1
XFILLER_0_3_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09505__B1 top.pc\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_199_3431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06670_ _01799_ _01808_ vssd1 vssd1 vccd1 vccd1 _01809_ sky130_fd_sc_hd__nor2_2
XANTENNA__07531__A2 net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08340_ _03286_ _03293_ vssd1 vssd1 vccd1 vccd1 _03474_ sky130_fd_sc_hd__nand2_1
XANTENNA__07819__B1 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_35_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08271_ _03316_ _03325_ net276 vssd1 vssd1 vccd1 vccd1 _03407_ sky130_fd_sc_hd__mux2_1
XANTENNA__13123__RESET_B net1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11105__B net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_99 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07222_ _02359_ _02360_ vssd1 vssd1 vccd1 vccd1 _02361_ sky130_fd_sc_hd__nor2_1
XANTENNA__08254__X _03391_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07153_ top.DUT.register\[23\]\[11\] net671 net647 top.DUT.register\[22\]\[11\] vssd1
+ vssd1 vccd1 vccd1 _02292_ sky130_fd_sc_hd__a22o_1
XANTENNA__10436__S net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07598__A2 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07084_ _02092_ _02136_ _02179_ _02222_ vssd1 vssd1 vccd1 vccd1 _02223_ sky130_fd_sc_hd__and4b_1
XFILLER_0_66_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1029_A net1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_2390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout391_A net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout136 net139 vssd1 vssd1 vccd1 vccd1 net136 sky130_fd_sc_hd__clkbuf_4
Xfanout147 _04724_ vssd1 vssd1 vccd1 vccd1 net147 sky130_fd_sc_hd__buf_2
XANTENNA_fanout489_A net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout158 _04916_ vssd1 vssd1 vccd1 vccd1 net158 sky130_fd_sc_hd__buf_2
XANTENNA__10171__S net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout169 net171 vssd1 vssd1 vccd1 vccd1 net169 sky130_fd_sc_hd__clkbuf_2
X_07986_ top.DUT.register\[29\]\[31\] net724 net717 top.DUT.register\[27\]\[31\] _03124_
+ vssd1 vssd1 vccd1 vccd1 _03125_ sky130_fd_sc_hd__a221o_1
XFILLER_0_199_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07770__A2 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09960__S net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09725_ top.a1.dataIn\[7\] _04750_ net407 vssd1 vssd1 vccd1 vccd1 _04753_ sky130_fd_sc_hd__a21o_1
X_06937_ top.DUT.register\[23\]\[21\] net673 net637 top.DUT.register\[6\]\[21\] vssd1
+ vssd1 vccd1 vccd1 _02076_ sky130_fd_sc_hd__a22o_1
XANTENNA__11303__B1 _05136_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout277_X net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout656_A _01609_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09656_ top.a1.halfData\[1\] _01471_ _04696_ net1086 vssd1 vssd1 vccd1 vccd1 _00116_
+ sky130_fd_sc_hd__o211a_1
XANTENNA__08429__X _03560_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06868_ _02005_ _02006_ vssd1 vssd1 vccd1 vccd1 _02007_ sky130_fd_sc_hd__nand2b_4
XANTENNA__07522__A2 net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07333__X _02472_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08607_ _02266_ _03073_ vssd1 vssd1 vccd1 vccd1 _03730_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_194_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09587_ top.pc\[29\] _04597_ top.pc\[30\] vssd1 vssd1 vccd1 vccd1 _04634_ sky130_fd_sc_hd__a21o_1
XFILLER_0_139_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06730__B1 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout444_X net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06799_ top.DUT.register\[28\]\[17\] net558 net452 top.DUT.register\[29\]\[17\] _01937_
+ vssd1 vssd1 vccd1 vccd1 _01938_ sky130_fd_sc_hd__a221o_1
XFILLER_0_210_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_648 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08538_ top.ramaddr\[12\] net832 net802 _03664_ vssd1 vssd1 vccd1 vccd1 _00030_ sky130_fd_sc_hd__a22o_1
XFILLER_0_210_799 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12395__Q top.a1.instruction\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_137_2500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08469_ _03171_ _03358_ _03366_ net279 vssd1 vssd1 vccd1 vccd1 _03598_ sky130_fd_sc_hd__o22a_2
XANTENNA_fanout611_X net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout709_X net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10500_ net1742 net255 net358 vssd1 vssd1 vccd1 vccd1 _00669_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11480_ _05328_ net273 _01396_ vssd1 vssd1 vccd1 vccd1 _05363_ sky130_fd_sc_hd__and3b_1
XFILLER_0_107_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08235__B1 _03370_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10431_ net267 net1823 net367 vssd1 vssd1 vccd1 vccd1 _00602_ sky130_fd_sc_hd__mux2_1
XANTENNA__10346__S net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_150_2700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08786__A1 net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08786__B2 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13150_ clknet_leaf_20_clk _00742_ net1033 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[20\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout980_X net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10362_ net2281 net144 net373 vssd1 vssd1 vccd1 vccd1 _00537_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_226 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06797__B1 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12101_ _05973_ _05975_ _05978_ vssd1 vssd1 vccd1 vccd1 _05984_ sky130_fd_sc_hd__and3_1
XFILLER_0_14_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10293_ net1406 net151 net387 vssd1 vssd1 vccd1 vccd1 _00471_ sky130_fd_sc_hd__mux2_1
X_13081_ clknet_leaf_13_clk _00673_ net955 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[18\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08538__A1 top.ramaddr\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12032_ _05895_ net125 vssd1 vssd1 vccd1 vccd1 _05915_ sky130_fd_sc_hd__nor2_1
XANTENNA__09735__B1 _04752_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold190 top.DUT.register\[15\]\[2\] vssd1 vssd1 vccd1 vccd1 net1306 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10081__S net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_148_2662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_148_2673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout670 _01599_ vssd1 vssd1 vccd1 vccd1 net670 sky130_fd_sc_hd__clkbuf_4
Xfanout681 _01547_ vssd1 vssd1 vccd1 vccd1 net681 sky130_fd_sc_hd__clkbuf_8
Xfanout692 _04050_ vssd1 vssd1 vccd1 vccd1 net692 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_70_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12934_ clknet_leaf_32_clk _00526_ net1045 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[13\]\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_161_2862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_16_Right_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_198_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_200_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12865_ clknet_leaf_16_clk _00457_ net964 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[11\]\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_158_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06721__B1 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_1_Left_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_185_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11816_ _01401_ _05690_ vssd1 vssd1 vccd1 vccd1 _05699_ sky130_fd_sc_hd__xnor2_2
XTAP_TAPCELL_ROW_194_3350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12796_ clknet_leaf_0_clk _00388_ net915 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[9\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_201_799 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_194_3361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_276 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11747_ _05603_ _05611_ _05620_ vssd1 vssd1 vccd1 vccd1 _05630_ sky130_fd_sc_hd__o21a_1
XFILLER_0_55_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09671__C1 net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11678_ _05557_ _05560_ vssd1 vssd1 vccd1 vccd1 _05561_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_510 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13417_ clknet_leaf_52_clk _01009_ net1034 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[28\]\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10256__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10629_ net146 net2220 net342 vssd1 vssd1 vccd1 vccd1 _00793_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_25_Right_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08234__B net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_180_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13348_ clknet_leaf_36_clk _00940_ net1049 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[26\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_738 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06788__B1 net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_47_Left_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_90_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13279_ clknet_leaf_24_clk _00871_ net1013 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[24\]\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08529__B2 net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11128__A3 net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08250__A net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_208_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11533__B1 top.a1.dataIn\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07840_ top.DUT.register\[21\]\[0\] net447 net507 top.DUT.register\[4\]\[0\] _02978_
+ vssd1 vssd1 vccd1 vccd1 _02979_ sky130_fd_sc_hd__a221o_1
XFILLER_0_208_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07752__A2 net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07771_ top.DUT.register\[7\]\[2\] net659 _02905_ _02907_ _02909_ vssd1 vssd1 vccd1
+ vccd1 _02910_ sky130_fd_sc_hd__a2111o_1
XPHY_EDGE_ROW_34_Right_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06960__B1 net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09510_ _01854_ _04560_ vssd1 vssd1 vccd1 vccd1 _04562_ sky130_fd_sc_hd__or2_1
X_06722_ top.DUT.register\[17\]\[25\] net746 _01860_ vssd1 vssd1 vccd1 vccd1 _01861_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_79_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_104_2009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09081__A top.a1.instruction\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07504__A2 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire412_X net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_604 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09441_ _04494_ _04495_ vssd1 vssd1 vccd1 vccd1 _04497_ sky130_fd_sc_hd__nor2_1
X_06653_ top.DUT.register\[9\]\[26\] net469 net529 top.DUT.register\[26\]\[26\] _01791_
+ vssd1 vssd1 vccd1 vccd1 _01792_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_56_Left_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06712__B1 net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_602 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09372_ top.pc\[17\] _04420_ vssd1 vssd1 vccd1 vccd1 _04432_ sky130_fd_sc_hd__or2_1
X_06584_ top.DUT.register\[28\]\[28\] net768 net741 top.DUT.register\[12\]\[28\] vssd1
+ vssd1 vccd1 vccd1 _01723_ sky130_fd_sc_hd__a22o_1
XFILLER_0_24_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08323_ _03342_ _03457_ vssd1 vssd1 vccd1 vccd1 _03458_ sky130_fd_sc_hd__nor2_1
XANTENNA__08465__B1 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10955__A _00016_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout237_A _04757_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_534 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_180 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_2230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08254_ _03263_ _03374_ _03390_ net430 _03388_ vssd1 vssd1 vccd1 vccd1 _03391_ sky130_fd_sc_hd__a221o_4
XANTENNA__08425__A net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_43_Right_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07205_ _01391_ net893 vssd1 vssd1 vccd1 vccd1 _02344_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_41_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10166__S net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08185_ _01572_ net330 vssd1 vssd1 vccd1 vccd1 _03323_ sky130_fd_sc_hd__nand2_1
XFILLER_0_172_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout404_A net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09955__S net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07136_ top.DUT.register\[11\]\[11\] net523 net519 top.DUT.register\[10\]\[11\] _02274_
+ vssd1 vssd1 vccd1 vccd1 _02275_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_132_2430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_598 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_65_Left_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07067_ top.DUT.register\[25\]\[22\] net778 net710 top.DUT.register\[11\]\[22\] vssd1
+ vssd1 vccd1 vccd1 _02206_ sky130_fd_sc_hd__a22o_1
XFILLER_0_140_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07991__A2 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout773_A _01614_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout394_X net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09193__A1 _02773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_52_Right_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07743__A2 net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07969_ top.DUT.register\[20\]\[31\] net566 net533 top.DUT.register\[12\]\[31\] _03107_
+ vssd1 vssd1 vccd1 vccd1 _03108_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout561_X net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout659_X net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09708_ top.a1.dataIn\[5\] net795 net798 top.pc\[5\] _04738_ vssd1 vssd1 vccd1 vccd1
+ _04739_ sky130_fd_sc_hd__a221o_1
X_10980_ top.a1.dataInTemp\[4\] _04999_ vssd1 vssd1 vccd1 vccd1 _05019_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_74_Left_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09639_ top.pad.keyCode\[5\] top.pad.keyCode\[6\] top.pad.keyCode\[7\] top.pad.keyCode\[4\]
+ vssd1 vssd1 vccd1 vccd1 _04681_ sky130_fd_sc_hd__or4b_2
XFILLER_0_179_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_143_2592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout826_X net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06703__B1 net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12650_ clknet_leaf_115_clk _00242_ net957 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[4\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_194_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11601_ _05409_ _05441_ vssd1 vssd1 vccd1 vccd1 _05484_ sky130_fd_sc_hd__xnor2_2
XANTENNA__11055__A2 net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_176_3080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12581_ clknet_leaf_33_clk _00173_ net1040 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[2\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_176_3091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_240 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_61_Right_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11532_ _05369_ _05413_ _05414_ vssd1 vssd1 vccd1 vccd1 _05415_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_80_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08335__A net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06407__X _01546_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10076__S net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11463_ _05317_ _05344_ vssd1 vssd1 vccd1 vccd1 _05346_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_151_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_83_Left_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09865__S net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13202_ clknet_leaf_25_clk _00794_ net1014 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[22\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_123_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_59_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10414_ net1319 net215 net369 vssd1 vssd1 vccd1 vccd1 _00586_ sky130_fd_sc_hd__mux2_1
X_11394_ _05260_ _05265_ _05276_ vssd1 vssd1 vccd1 vccd1 _05277_ sky130_fd_sc_hd__a21bo_1
X_13133_ clknet_leaf_42_clk _00725_ net1064 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[19\]\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_150_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10804__S net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10345_ net1882 net225 net379 vssd1 vssd1 vccd1 vccd1 _00521_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09708__B1 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13064_ clknet_leaf_27_clk _00656_ net1008 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[17\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08070__A _02156_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10276_ net1501 net208 net388 vssd1 vssd1 vccd1 vccd1 _00454_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_70_Right_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12015_ _05897_ vssd1 vssd1 vccd1 vccd1 _05898_ sky130_fd_sc_hd__inv_2
XFILLER_0_206_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08931__A1 _03122_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07734__A2 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_205_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_205_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06942__B1 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_502 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_17_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12917_ clknet_leaf_32_clk _00509_ net1023 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[13\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11294__A2 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12848_ clknet_leaf_28_clk _00440_ net1010 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[10\]\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_201_574 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_158_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_68 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12779_ clknet_leaf_46_clk _00371_ net1065 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[8\]\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_83_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08998__A1 net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_211_3604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_211_3615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_211_3626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold904 top.DUT.register\[21\]\[6\] vssd1 vssd1 vccd1 vccd1 net2020 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08214__A3 net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold915 top.a1.row1\[108\] vssd1 vssd1 vccd1 vccd1 net2031 sky130_fd_sc_hd__dlygate4sd3_1
Xhold926 top.DUT.register\[18\]\[15\] vssd1 vssd1 vccd1 vccd1 net2042 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08899__B _04008_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold937 top.DUT.register\[21\]\[10\] vssd1 vssd1 vccd1 vccd1 net2053 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_114_2160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold948 top.DUT.register\[29\]\[30\] vssd1 vssd1 vccd1 vccd1 net2064 sky130_fd_sc_hd__dlygate4sd3_1
Xhold959 top.DUT.register\[1\]\[26\] vssd1 vssd1 vccd1 vccd1 net2075 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_177_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09990_ net229 net1731 net623 vssd1 vssd1 vccd1 vccd1 _00195_ sky130_fd_sc_hd__mux2_1
XANTENNA__10714__S net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_177_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07973__A2 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08941_ net1295 net831 net801 _04048_ vssd1 vssd1 vccd1 vccd1 _00049_ sky130_fd_sc_hd__a22o_1
XFILLER_0_209_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08872_ _01745_ net493 net433 _01744_ vssd1 vssd1 vccd1 vccd1 _03983_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_209_3577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07186__B1 net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_209_3588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06212__B net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07725__A2 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07823_ top.DUT.register\[5\]\[0\] net651 net742 top.DUT.register\[2\]\[0\] vssd1
+ vssd1 vccd1 vccd1 _02962_ sky130_fd_sc_hd__a22o_1
XFILLER_0_208_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06933__B1 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout187_A _04832_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07754_ top.DUT.register\[14\]\[3\] net585 net462 top.DUT.register\[17\]\[3\] _02892_
+ vssd1 vssd1 vccd1 vccd1 _02893_ sky130_fd_sc_hd__a221o_1
XFILLER_0_211_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_168_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06705_ top.DUT.register\[15\]\[25\] net679 net675 top.DUT.register\[31\]\[25\] vssd1
+ vssd1 vccd1 vccd1 _01844_ sky130_fd_sc_hd__a22o_1
XANTENNA__11285__A2 _05136_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07685_ top.DUT.register\[20\]\[4\] net665 net658 top.DUT.register\[21\]\[4\] vssd1
+ vssd1 vccd1 vccd1 _02824_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout354_A _04989_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1096_A net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_91_clk clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_91_clk
+ sky130_fd_sc_hd__clkbuf_8
X_09424_ net137 _04480_ vssd1 vssd1 vccd1 vccd1 _04481_ sky130_fd_sc_hd__nor2_1
X_06636_ top.DUT.register\[23\]\[27\] net673 net729 top.DUT.register\[18\]\[27\] vssd1
+ vssd1 vccd1 vccd1 _01775_ sky130_fd_sc_hd__a22o_1
XFILLER_0_149_456 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09355_ top.pc\[16\] _04403_ vssd1 vssd1 vccd1 vccd1 _04416_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout521_A net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06567_ top.DUT.register\[13\]\[28\] net464 net525 top.DUT.register\[11\]\[28\] _01705_
+ vssd1 vssd1 vccd1 vccd1 _01706_ sky130_fd_sc_hd__a221o_1
XANTENNA__13065__CLK clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout619_A net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10245__A0 net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08306_ net298 _03440_ _03439_ vssd1 vssd1 vccd1 vccd1 _03441_ sky130_fd_sc_hd__o21a_2
X_09286_ net821 _02363_ vssd1 vssd1 vccd1 vccd1 _04351_ sky130_fd_sc_hd__and2_1
XFILLER_0_145_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08155__A _02773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06498_ net788 _01596_ _01600_ vssd1 vssd1 vccd1 vccd1 _01637_ sky130_fd_sc_hd__and3_4
XANTENNA__07110__B1 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_830 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_7_clk_A clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08237_ net317 _03373_ _03363_ vssd1 vssd1 vccd1 vccd1 _03374_ sky130_fd_sc_hd__a21o_1
XFILLER_0_7_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout407_X net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_479 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08168_ _03302_ _03305_ net287 vssd1 vssd1 vccd1 vccd1 _03306_ sky130_fd_sc_hd__mux2_1
XANTENNA__11012__C net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout890_A net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout988_A net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07119_ top.DUT.register\[24\]\[16\] net644 net743 top.DUT.register\[2\]\[16\] _02253_
+ vssd1 vssd1 vccd1 vccd1 _02258_ sky130_fd_sc_hd__a221o_1
XFILLER_0_120_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10624__S net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08099_ net319 net298 vssd1 vssd1 vccd1 vccd1 _03238_ sky130_fd_sc_hd__nor2_1
XANTENNA__12902__CLK clknet_leaf_40_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10130_ net217 net1681 net608 vssd1 vssd1 vccd1 vccd1 _00330_ sky130_fd_sc_hd__mux2_1
XANTENNA__07964__A2 net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout776_X net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_54_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_54_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10061_ net1845 net196 net616 vssd1 vssd1 vccd1 vccd1 _00263_ sky130_fd_sc_hd__mux2_1
XANTENNA__13297__RESET_B net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07177__B1 net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09714__A net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_2621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06924__B1 net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13820_ net1104 vssd1 vssd1 vccd1 vccd1 gpio_out[15] sky130_fd_sc_hd__buf_2
XFILLER_0_203_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_178_3120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13751_ clknet_leaf_99_clk _01322_ vssd1 vssd1 vccd1 vccd1 top.lcd.cnt_20ms\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_3_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10963_ top.a1.dataIn\[0\] net850 _04667_ net888 _05005_ vssd1 vssd1 vccd1 vccd1
+ _05006_ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_82_clk clknet_4_6__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_82_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08992__C_N _03777_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_376 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12702_ clknet_leaf_18_clk _00294_ net1028 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[6\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13682_ clknet_leaf_90_clk _01258_ net999 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08617__X _03740_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10894_ top.DUT.register\[30\]\[6\] net242 net478 vssd1 vssd1 vccd1 vccd1 _01055_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12633_ clknet_leaf_14_clk _00225_ net955 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[4\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_183_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11190__S net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_182_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12564_ clknet_leaf_58_clk _00156_ net1075 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[2\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_91_Left_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07101__B1 net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_182_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11515_ _05375_ _05379_ _05395_ _05397_ vssd1 vssd1 vccd1 vccd1 _05398_ sky130_fd_sc_hd__a211o_2
XTAP_TAPCELL_ROW_156_2783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12495_ clknet_leaf_93_clk _00087_ net1000 vssd1 vssd1 vccd1 vccd1 top.pc\[7\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_108_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11446_ top.a1.dataIn\[16\] _05326_ _05327_ vssd1 vssd1 vccd1 vccd1 _05329_ sky130_fd_sc_hd__or3_1
XANTENNA__10539__A1 _04760_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_507 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10534__S net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08601__B1 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_189_3282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11377_ _05255_ _05256_ _05259_ vssd1 vssd1 vccd1 vccd1 _05260_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_0_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13116_ clknet_leaf_130_clk _00708_ net910 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[19\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_10328_ _04153_ _04713_ net400 vssd1 vssd1 vccd1 vccd1 _04980_ sky130_fd_sc_hd__and3_1
XFILLER_0_147_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13047_ clknet_leaf_2_clk _00639_ net918 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[17\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_10259_ net155 net2287 net391 vssd1 vssd1 vccd1 vccd1 _00438_ sky130_fd_sc_hd__mux2_1
XANTENNA__07707__A2 net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06915__B1 net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10711__A1 net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09343__B _02589_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_507 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09062__C _03623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11267__A2 _05149_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_73_clk clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_73_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_76_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07470_ _02601_ _02608_ vssd1 vssd1 vccd1 vccd1 _02609_ sky130_fd_sc_hd__or2_2
XANTENNA__07340__B1 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_724 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06421_ top.DUT.register\[7\]\[30\] net517 net513 top.DUT.register\[24\]\[30\] vssd1
+ vssd1 vccd1 vccd1 _01560_ sky130_fd_sc_hd__a22o_1
XFILLER_0_201_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11019__A2 net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10709__S net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_711 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09140_ _04211_ _04212_ vssd1 vssd1 vccd1 vccd1 _04214_ sky130_fd_sc_hd__and2_1
X_06352_ top.pad.button_control.r_counter\[5\] top.pad.button_control.r_counter\[6\]
+ top.pad.button_control.r_counter\[7\] vssd1 vssd1 vccd1 vccd1 _01492_ sky130_fd_sc_hd__o21a_1
XFILLER_0_16_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09071_ net894 _01485_ vssd1 vssd1 vccd1 vccd1 _04146_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_20_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06283_ _01437_ _01443_ _01445_ vssd1 vssd1 vccd1 vccd1 _01446_ sky130_fd_sc_hd__nor3_2
XANTENNA__08840__B1 top.pc\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_479 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_800 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06207__B net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08022_ net333 _03142_ _03151_ _03159_ vssd1 vssd1 vccd1 vccd1 _03161_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_142_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold701 top.DUT.register\[19\]\[29\] vssd1 vssd1 vccd1 vccd1 net1817 sky130_fd_sc_hd__dlygate4sd3_1
Xhold712 top.DUT.register\[21\]\[18\] vssd1 vssd1 vccd1 vccd1 net1828 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10952__B _04668_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold723 top.DUT.register\[16\]\[5\] vssd1 vssd1 vccd1 vccd1 net1839 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_112_2119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold734 top.DUT.register\[5\]\[2\] vssd1 vssd1 vccd1 vccd1 net1850 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_96_1885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10444__S net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold745 top.DUT.register\[16\]\[28\] vssd1 vssd1 vccd1 vccd1 net1861 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold756 top.DUT.register\[12\]\[31\] vssd1 vssd1 vccd1 vccd1 net1872 sky130_fd_sc_hd__dlygate4sd3_1
Xhold767 top.DUT.register\[27\]\[5\] vssd1 vssd1 vccd1 vccd1 net1883 sky130_fd_sc_hd__dlygate4sd3_1
Xhold778 top.DUT.register\[3\]\[23\] vssd1 vssd1 vccd1 vccd1 net1894 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09973_ net1873 net157 net630 vssd1 vssd1 vccd1 vccd1 _00181_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_139_Left_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold789 top.DUT.register\[11\]\[20\] vssd1 vssd1 vccd1 vccd1 net1905 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08924_ _03145_ _04031_ vssd1 vssd1 vccd1 vccd1 _04032_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07159__B1 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1011_A net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08855_ net424 _03966_ _03955_ net497 vssd1 vssd1 vccd1 vccd1 _03967_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA_fanout471_A net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout569_A _01525_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_2351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_2_Right_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07806_ _02925_ _02944_ vssd1 vssd1 vccd1 vccd1 _02945_ sky130_fd_sc_hd__and2_1
X_08786_ net319 _03555_ _03734_ net274 vssd1 vssd1 vccd1 vccd1 _03901_ sky130_fd_sc_hd__a22o_1
XFILLER_0_211_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11258__A2 _05149_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07737_ _02870_ _02872_ _02874_ _02875_ vssd1 vssd1 vccd1 vccd1 _02876_ sky130_fd_sc_hd__or4_1
XANTENNA__08659__B1 _03264_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout736_A net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_64_clk clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_64_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08123__A2 _03176_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout357_X net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_2540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_2551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07668_ _02359_ _02805_ _02806_ _01580_ vssd1 vssd1 vccd1 vccd1 _02807_ sky130_fd_sc_hd__o211a_1
XPHY_EDGE_ROW_148_Left_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07331__B1 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09407_ top.pc\[19\] _04453_ vssd1 vssd1 vccd1 vccd1 _04465_ sky130_fd_sc_hd__nor2_1
X_06619_ top.DUT.register\[1\]\[27\] net445 _01755_ _01757_ vssd1 vssd1 vccd1 vccd1
+ _01758_ sky130_fd_sc_hd__a211o_1
XANTENNA__06685__A2 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10619__S net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_746 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07599_ top.DUT.register\[5\]\[6\] net651 net635 top.DUT.register\[6\]\[6\] _02736_
+ vssd1 vssd1 vccd1 vccd1 _02738_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout524_X net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09338_ _04398_ _04399_ vssd1 vssd1 vccd1 vccd1 _04400_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_192_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09269_ _01579_ _01583_ vssd1 vssd1 vccd1 vccd1 _04335_ sky130_fd_sc_hd__and2_2
XFILLER_0_105_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11300_ net879 _05122_ top.lcd.nextState\[3\] vssd1 vssd1 vccd1 vccd1 _05188_ sky130_fd_sc_hd__and3b_1
XFILLER_0_16_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12280_ net1966 _06097_ _06098_ vssd1 vssd1 vccd1 vccd1 _01344_ sky130_fd_sc_hd__o21a_1
XANTENNA__09709__A net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_490 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11231_ _05120_ _05123_ vssd1 vssd1 vccd1 vccd1 _05124_ sky130_fd_sc_hd__and2_1
XANTENNA__10354__S net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07398__B1 net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11162_ _01385_ _01418_ _01409_ vssd1 vssd1 vccd1 vccd1 _05090_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_101_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10113_ net146 net1996 net607 vssd1 vssd1 vccd1 vccd1 _00313_ sky130_fd_sc_hd__mux2_1
X_11093_ net68 net864 vssd1 vssd1 vccd1 vccd1 _05052_ sky130_fd_sc_hd__and2_1
XANTENNA_input32_A DAT_I[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09444__A _02070_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10044_ net2189 net149 net620 vssd1 vssd1 vccd1 vccd1 _00247_ sky130_fd_sc_hd__mux2_1
XANTENNA__06420__X _01559_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold50 top.ramstore\[20\] vssd1 vssd1 vccd1 vccd1 net1166 sky130_fd_sc_hd__dlygate4sd3_1
Xhold61 _01161_ vssd1 vssd1 vccd1 vccd1 net1177 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold72 net79 vssd1 vssd1 vccd1 vccd1 net1188 sky130_fd_sc_hd__dlygate4sd3_1
Xhold83 top.ramstore\[13\] vssd1 vssd1 vccd1 vccd1 net1199 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold94 net95 vssd1 vssd1 vccd1 vccd1 net1210 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07570__B1 net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13803_ clknet_leaf_71_clk _01372_ net1087 vssd1 vssd1 vccd1 vccd1 top.pad.keyCode\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_11995_ _05865_ _05872_ _05874_ _05876_ vssd1 vssd1 vccd1 vccd1 _05878_ sky130_fd_sc_hd__a211o_1
XFILLER_0_58_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_55_clk clknet_4_12__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_55_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__09311__A1 net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13734_ clknet_leaf_94_clk _01305_ vssd1 vssd1 vccd1 vccd1 top.a1.dataInTemp\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__09311__B2 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10946_ net1392 net166 net592 vssd1 vssd1 vccd1 vccd1 _01107_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_27_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07322__B1 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_158_2812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_404 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_158_2823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06676__A2 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13665_ clknet_leaf_91_clk _01241_ net996 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[115\]
+ sky130_fd_sc_hd__dfrtp_1
X_10877_ net193 net1875 net597 vssd1 vssd1 vccd1 vccd1 _01038_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_763 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12616_ clknet_leaf_7_clk _00208_ net946 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[3\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_651 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13596_ clknet_leaf_46_clk net1183 net1067 vssd1 vssd1 vccd1 vccd1 net88 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_171_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_143_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12547_ clknet_leaf_61_clk _00139_ net1088 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[1\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_170_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12478_ clknet_leaf_47_clk _00073_ net1067 vssd1 vssd1 vccd1 vccd1 top.ramstore\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_3 _02748_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11429_ _05269_ _05311_ vssd1 vssd1 vccd1 vccd1 _05312_ sky130_fd_sc_hd__nand2_1
XANTENNA__10264__S net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07389__B1 net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09057__C _03737_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_191_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06600__A2 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_169_2974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_169_2985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06970_ top.DUT.register\[30\]\[23\] net581 net468 top.DUT.register\[9\]\[23\] _02108_
+ vssd1 vssd1 vccd1 vccd1 _02109_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_206_3536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1070 net1071 vssd1 vssd1 vccd1 vccd1 net1070 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_174_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08640_ _03761_ vssd1 vssd1 vccd1 vccd1 _03762_ sky130_fd_sc_hd__inv_2
Xfanout1081 net1082 vssd1 vssd1 vccd1 vccd1 net1081 sky130_fd_sc_hd__clkbuf_4
Xfanout1092 net1093 vssd1 vssd1 vccd1 vccd1 net1092 sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_175_Right_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_109_2081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_178_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08571_ _03498_ _03533_ _03695_ vssd1 vssd1 vccd1 vccd1 _03696_ sky130_fd_sc_hd__a21o_1
XFILLER_0_83_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_46_clk clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_46_clk
+ sky130_fd_sc_hd__clkbuf_8
X_07522_ top.DUT.register\[9\]\[7\] net467 net439 top.DUT.register\[5\]\[7\] _02660_
+ vssd1 vssd1 vccd1 vccd1 _02661_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_122_2270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_122_2281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06667__A2 net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07453_ top.DUT.register\[30\]\[15\] net759 net715 top.DUT.register\[27\]\[15\] vssd1
+ vssd1 vccd1 vccd1 _02592_ sky130_fd_sc_hd__a22o_1
XFILLER_0_147_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10439__S net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06404_ top.DUT.register\[19\]\[30\] net537 net534 top.DUT.register\[12\]\[30\] vssd1
+ vssd1 vccd1 vccd1 _01543_ sky130_fd_sc_hd__a22o_1
XANTENNA__09066__B1 _04140_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07384_ _02497_ _02522_ vssd1 vssd1 vccd1 vccd1 _02523_ sky130_fd_sc_hd__nor2_1
XFILLER_0_123_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_174_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09123_ _04190_ _04194_ _04196_ _04197_ _01505_ vssd1 vssd1 vccd1 vccd1 _04198_ sky130_fd_sc_hd__o311a_1
XTAP_TAPCELL_ROW_98_1914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06335_ top.d_ready _01475_ _01480_ vssd1 vssd1 vccd1 vccd1 _01481_ sky130_fd_sc_hd__nor3_1
XFILLER_0_96_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout317_A net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1059_A net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09054_ _04125_ _04126_ _04127_ _04128_ vssd1 vssd1 vccd1 vccd1 _04129_ sky130_fd_sc_hd__or4_1
X_06266_ top.ramload\[27\] net854 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedData\[27\]
+ sky130_fd_sc_hd__and2_1
XANTENNA__07092__A2 net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08005_ _03122_ _03142_ vssd1 vssd1 vccd1 vccd1 _03144_ sky130_fd_sc_hd__nand2_1
Xhold520 top.DUT.register\[5\]\[27\] vssd1 vssd1 vccd1 vccd1 net1636 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10174__S net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_38_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06197_ wb.curr_state\[2\] wb.curr_state\[1\] vssd1 vssd1 vccd1 vccd1 _01428_ sky130_fd_sc_hd__or2_2
Xhold531 top.DUT.register\[19\]\[12\] vssd1 vssd1 vccd1 vccd1 net1647 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_38_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold542 top.DUT.register\[31\]\[16\] vssd1 vssd1 vccd1 vccd1 net1658 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09963__S net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold553 top.DUT.register\[18\]\[8\] vssd1 vssd1 vccd1 vccd1 net1669 sky130_fd_sc_hd__dlygate4sd3_1
Xhold564 top.DUT.register\[28\]\[20\] vssd1 vssd1 vccd1 vccd1 net1680 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold575 top.DUT.register\[4\]\[0\] vssd1 vssd1 vccd1 vccd1 net1691 sky130_fd_sc_hd__dlygate4sd3_1
Xhold586 top.DUT.register\[28\]\[9\] vssd1 vssd1 vccd1 vccd1 net1702 sky130_fd_sc_hd__dlygate4sd3_1
Xhold597 top.DUT.register\[11\]\[24\] vssd1 vssd1 vccd1 vccd1 net1713 sky130_fd_sc_hd__dlygate4sd3_1
X_09956_ net1989 net220 net627 vssd1 vssd1 vccd1 vccd1 _00164_ sky130_fd_sc_hd__mux2_1
XANTENNA__10902__S net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_5_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08907_ net325 _03690_ vssd1 vssd1 vccd1 vccd1 _04016_ sky130_fd_sc_hd__nor2_1
X_09887_ _03968_ net407 vssd1 vssd1 vccd1 vccd1 _04896_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout474_X net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout853_A net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09541__A1 _01754_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08838_ _03930_ _03950_ vssd1 vssd1 vccd1 vccd1 _03951_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_142_Right_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07552__B1 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12398__Q top.a1.instruction\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08769_ net426 _03881_ _03882_ _03884_ _03880_ vssd1 vssd1 vccd1 vccd1 _03885_ sky130_fd_sc_hd__a2111o_1
XANTENNA_fanout641_X net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_37_clk clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_37_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout739_X net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06646__A_N _01764_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10800_ net235 net1901 net599 vssd1 vssd1 vccd1 vccd1 _00961_ sky130_fd_sc_hd__mux2_1
X_11780_ top.a1.dataIn\[8\] _05655_ _05656_ vssd1 vssd1 vccd1 vccd1 _05663_ sky130_fd_sc_hd__and3_1
XANTENNA__11100__A1 net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09844__A2 net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12453__RESET_B net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10731_ net1581 net259 net419 vssd1 vssd1 vccd1 vccd1 _00892_ sky130_fd_sc_hd__mux2_1
XANTENNA__10349__S net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06658__A2 net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout906_X net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_171_3009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13450_ clknet_leaf_115_clk _01042_ net963 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[29\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10662_ net1687 net145 net338 vssd1 vssd1 vccd1 vccd1 _00825_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_338 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12401_ clknet_leaf_103_clk top.ru.next_FetchedInstr\[13\] net976 vssd1 vssd1 vccd1
+ vccd1 top.a1.instruction\[13\] sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_62_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13381_ clknet_leaf_33_clk _00973_ net1042 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[27\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_10593_ net1356 net150 net351 vssd1 vssd1 vccd1 vccd1 _00759_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_153_2742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12332_ _06131_ net790 _06130_ vssd1 vssd1 vccd1 vccd1 _01363_ sky130_fd_sc_hd__and3b_1
XANTENNA__08280__A1 net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06415__X _01554_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08280__B2 net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06830__A2 net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12263_ _01435_ net686 _06088_ vssd1 vssd1 vccd1 vccd1 _01337_ sky130_fd_sc_hd__and3_1
XANTENNA__10084__S net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_186_3230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_186_3241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11214_ _04664_ _05100_ vssd1 vssd1 vccd1 vccd1 _05113_ sky130_fd_sc_hd__and2_1
X_12194_ net1126 _06046_ net688 vssd1 vssd1 vccd1 vccd1 _01301_ sky130_fd_sc_hd__mux2_1
Xoutput40 net40 vssd1 vssd1 vccd1 vccd1 ADR_O[0] sky130_fd_sc_hd__buf_2
XANTENNA__08997__B _03580_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput51 net51 vssd1 vssd1 vccd1 vccd1 ADR_O[1] sky130_fd_sc_hd__buf_2
Xoutput62 net62 vssd1 vssd1 vccd1 vccd1 ADR_O[2] sky130_fd_sc_hd__buf_2
Xoutput73 net73 vssd1 vssd1 vccd1 vccd1 DAT_O[0] sky130_fd_sc_hd__clkbuf_4
X_11145_ _01333_ _01469_ vssd1 vssd1 vccd1 vccd1 _05078_ sky130_fd_sc_hd__nand2_1
XFILLER_0_208_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_207_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput84 net84 vssd1 vssd1 vccd1 vccd1 DAT_O[1] sky130_fd_sc_hd__clkbuf_4
XANTENNA__10812__S net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07791__B1 net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput95 net95 vssd1 vssd1 vccd1 vccd1 DAT_O[2] sky130_fd_sc_hd__buf_2
XANTENNA__07246__X _02385_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09174__A _02773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11076_ net92 net872 net836 net1197 vssd1 vssd1 vccd1 vccd1 _01187_ sky130_fd_sc_hd__a22o_1
XFILLER_0_207_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_94_clk_A clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13692__Q top.lcd.nextState\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09532__A1 _01505_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10027_ net1620 net210 net620 vssd1 vssd1 vccd1 vccd1 _00230_ sky130_fd_sc_hd__mux2_1
XFILLER_0_208_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06897__A2 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_203_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_28_clk clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_28_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_201_3455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_201_3466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11978_ _05859_ _05860_ _05858_ vssd1 vssd1 vccd1 vccd1 _05861_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_53_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_175_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09835__A2 net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13717_ clknet_leaf_96_clk _01288_ net984 vssd1 vssd1 vccd1 vccd1 top.a1.row2\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_10929_ net1985 net232 net593 vssd1 vssd1 vccd1 vccd1 _01090_ sky130_fd_sc_hd__mux2_1
XANTENNA__10259__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_184_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_582 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13126__CLK clknet_leaf_40_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_32_clk_A clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13648_ clknet_leaf_89_clk _01227_ net1003 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[56\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_171_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13579_ clknet_leaf_106_clk net1218 net970 vssd1 vssd1 vccd1 vccd1 net101 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07074__A2 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13329__RESET_B net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_47_clk_A clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_460 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_1844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_99_Right_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout307 _02925_ vssd1 vssd1 vccd1 vccd1 net307 sky130_fd_sc_hd__dlymetal6s2s_1
X_09810_ _04825_ _04826_ vssd1 vssd1 vccd1 vccd1 _04827_ sky130_fd_sc_hd__nor2_1
XANTENNA__10722__S net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09771__B2 top.a1.dataIn\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout318 _02830_ vssd1 vssd1 vccd1 vccd1 net318 sky130_fd_sc_hd__clkbuf_2
Xfanout329 net332 vssd1 vssd1 vccd1 vccd1 net329 sky130_fd_sc_hd__clkbuf_2
XANTENNA__06585__A1 top.DUT.register\[6\]\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07782__B1 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09084__A top.a1.instruction\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09741_ _03638_ net403 net488 _04765_ vssd1 vssd1 vccd1 vccd1 _04766_ sky130_fd_sc_hd__o211a_4
X_06953_ _02090_ _02091_ vssd1 vssd1 vccd1 vccd1 _02092_ sky130_fd_sc_hd__nor2_1
XANTENNA_clkbuf_leaf_105_clk_A clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09672_ _01500_ _01507_ net793 vssd1 vssd1 vccd1 vccd1 _04708_ sky130_fd_sc_hd__or3_4
X_06884_ top.DUT.register\[22\]\[18\] net576 net533 top.DUT.register\[12\]\[18\] vssd1
+ vssd1 vccd1 vccd1 _02023_ sky130_fd_sc_hd__a22o_1
XANTENNA__07534__B1 net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06220__B net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_124_2310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08623_ net886 top.pc\[16\] net697 _03745_ vssd1 vssd1 vccd1 vccd1 _03746_ sky130_fd_sc_hd__a22o_1
XANTENNA__06888__A2 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13107__Q top.DUT.register\[19\]\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10958__A net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_19_clk clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_19_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_11_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout267_A _04726_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08554_ _02431_ net431 net428 _03673_ _03679_ vssd1 vssd1 vccd1 vccd1 _03680_ sky130_fd_sc_hd__a221o_1
XANTENNA__08428__A net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07505_ _02638_ _02640_ _02641_ _02643_ vssd1 vssd1 vccd1 vccd1 _02644_ sky130_fd_sc_hd__or4_2
XFILLER_0_187_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10169__S net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08485_ _02389_ _03613_ vssd1 vssd1 vccd1 vccd1 _03614_ sky130_fd_sc_hd__and2_1
XFILLER_0_175_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout434_A _03169_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_532 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10396__C _04708_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09958__S net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07436_ top.DUT.register\[25\]\[15\] net455 net516 top.DUT.register\[7\]\[15\] _02574_
+ vssd1 vssd1 vccd1 vccd1 _02575_ sky130_fd_sc_hd__a221o_1
XFILLER_0_91_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_102_1973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_190_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_749 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07367_ top.DUT.register\[23\]\[8\] net672 net715 top.DUT.register\[27\]\[8\] _02505_
+ vssd1 vssd1 vccd1 vccd1 _02506_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout601_A _04965_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_162_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09106_ _04172_ _04179_ vssd1 vssd1 vccd1 vccd1 _04181_ sky130_fd_sc_hd__nand2_1
XFILLER_0_45_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06318_ _01334_ _01460_ _01470_ vssd1 vssd1 vccd1 vccd1 _00004_ sky130_fd_sc_hd__o21a_1
XFILLER_0_60_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07065__A2 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_758 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07298_ top.DUT.register\[18\]\[12\] net547 net523 top.DUT.register\[11\]\[12\] vssd1
+ vssd1 vccd1 vccd1 _02437_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_135_2472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09037_ _04105_ _04106_ _04111_ _04104_ vssd1 vssd1 vccd1 vccd1 _04112_ sky130_fd_sc_hd__o31a_1
X_06249_ net2313 net855 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedData\[10\] sky130_fd_sc_hd__and2_1
XFILLER_0_102_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06812__A2 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11149__A1 _01393_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_211_Right_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold350 top.DUT.register\[18\]\[18\] vssd1 vssd1 vccd1 vccd1 net1466 sky130_fd_sc_hd__dlygate4sd3_1
Xhold361 top.DUT.register\[15\]\[15\] vssd1 vssd1 vccd1 vccd1 net1477 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout591_X net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold372 top.DUT.register\[12\]\[13\] vssd1 vssd1 vccd1 vccd1 net1488 sky130_fd_sc_hd__dlygate4sd3_1
Xhold383 top.DUT.register\[5\]\[16\] vssd1 vssd1 vccd1 vccd1 net1499 sky130_fd_sc_hd__dlygate4sd3_1
Xhold394 top.DUT.register\[15\]\[5\] vssd1 vssd1 vccd1 vccd1 net1510 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10632__S net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07773__B1 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout830 net832 vssd1 vssd1 vccd1 vccd1 net830 sky130_fd_sc_hd__buf_2
Xfanout841 net842 vssd1 vssd1 vccd1 vccd1 net841 sky130_fd_sc_hd__buf_2
Xfanout852 net855 vssd1 vssd1 vccd1 vccd1 net852 sky130_fd_sc_hd__buf_2
X_09939_ top.a1.instruction\[31\] net486 net401 top.a1.dataIn\[31\] net397 vssd1 vssd1
+ vccd1 vccd1 _04944_ sky130_fd_sc_hd__a221o_2
XANTENNA_fanout856_X net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout863 _01428_ vssd1 vssd1 vccd1 vccd1 net863 sky130_fd_sc_hd__buf_2
Xfanout874 net875 vssd1 vssd1 vccd1 vccd1 net874 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_181_3160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout885 top.ru.state\[5\] vssd1 vssd1 vccd1 vccd1 net885 sky130_fd_sc_hd__clkbuf_4
Xfanout896 top.a1.instruction\[4\] vssd1 vssd1 vccd1 vccd1 net896 sky130_fd_sc_hd__buf_2
X_12950_ clknet_leaf_4_clk _00542_ net940 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[14\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07525__B1 net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1050 top.DUT.register\[16\]\[7\] vssd1 vssd1 vccd1 vccd1 net2166 sky130_fd_sc_hd__dlygate4sd3_1
X_11901_ _05779_ _05781_ _05782_ vssd1 vssd1 vccd1 vccd1 _05784_ sky130_fd_sc_hd__nand3_1
Xhold1061 top.DUT.register\[13\]\[3\] vssd1 vssd1 vccd1 vccd1 net2177 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1072 top.DUT.register\[7\]\[28\] vssd1 vssd1 vccd1 vccd1 net2188 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06879__A2 net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1083 top.DUT.register\[30\]\[10\] vssd1 vssd1 vccd1 vccd1 net2199 sky130_fd_sc_hd__dlygate4sd3_1
X_12881_ clknet_leaf_116_clk _00473_ net957 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[12\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1094 top.DUT.register\[17\]\[25\] vssd1 vssd1 vccd1 vccd1 net2210 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11832_ _05681_ _05714_ vssd1 vssd1 vccd1 vccd1 _05715_ sky130_fd_sc_hd__xnor2_2
XANTENNA__07513__Y _02652_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_169_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11763_ _05635_ _05645_ vssd1 vssd1 vccd1 vccd1 _05646_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_68_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13502_ clknet_leaf_21_clk _01094_ net1034 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[31\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_10714_ net2298 net206 net336 vssd1 vssd1 vccd1 vccd1 _00875_ sky130_fd_sc_hd__mux2_1
X_11694_ _05544_ _05576_ vssd1 vssd1 vccd1 vccd1 _05577_ sky130_fd_sc_hd__nor2_2
XFILLER_0_71_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13433_ clknet_leaf_118_clk _01025_ net956 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[29\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_180_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10645_ net225 net2196 net343 vssd1 vssd1 vccd1 vccd1 _00809_ sky130_fd_sc_hd__mux2_1
XANTENNA__10807__S net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09045__A3 _03370_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07056__A2 net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13364_ clknet_leaf_56_clk _00956_ net1075 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[27\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_63_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10576_ net1420 net208 net351 vssd1 vssd1 vccd1 vccd1 _00742_ sky130_fd_sc_hd__mux2_1
X_12315_ net2132 _06118_ net790 vssd1 vssd1 vccd1 vccd1 _06121_ sky130_fd_sc_hd__o21ai_1
XANTENNA__06803__A2 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11311__C_N top.lcd.nextState\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13295_ clknet_leaf_22_clk _00887_ net1022 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[24\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_12246_ top.lcd.cnt_20ms\[13\] top.lcd.cnt_20ms\[12\] _06075_ vssd1 vssd1 vccd1 vccd1
+ _06079_ sky130_fd_sc_hd__and3_1
XFILLER_0_139_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_75_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12177_ _05948_ _05083_ net846 net1288 vssd1 vssd1 vccd1 vccd1 _01285_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__10542__S _04989_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07937__A_N _02026_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_166_2933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11128_ net906 net1298 net861 _05069_ vssd1 vssd1 vccd1 vccd1 _01215_ sky130_fd_sc_hd__a31o_1
XANTENNA__08308__A2 _03441_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09505__A1 top.pc\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11059_ net1193 net866 net837 top.ramstore\[10\] vssd1 vssd1 vccd1 vccd1 _01170_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_199_3432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_106_2040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_148_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_157_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_156_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08270_ net296 _03405_ vssd1 vssd1 vccd1 vccd1 _03406_ sky130_fd_sc_hd__and2_1
XFILLER_0_73_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_671 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07221_ top.a1.instruction\[30\] net789 net793 top.a1.instruction\[22\] vssd1 vssd1
+ vccd1 vccd1 _02360_ sky130_fd_sc_hd__a22o_1
XFILLER_0_104_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10717__S net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07152_ top.DUT.register\[15\]\[11\] net706 net698 top.DUT.register\[31\]\[11\] vssd1
+ vssd1 vccd1 vccd1 _02291_ sky130_fd_sc_hd__a22o_1
XANTENNA__09079__A top.a1.instruction\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07047__A2 net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11121__B net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07083_ _02220_ _02221_ vssd1 vssd1 vccd1 vccd1 _02222_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_112_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_8_clk clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_8_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_140_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06215__B net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_196_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09744__A1 top.pc\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10452__S net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_2391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout126 _05879_ vssd1 vssd1 vccd1 vccd1 net126 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_10_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07755__B1 net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout137 net139 vssd1 vssd1 vccd1 vccd1 net137 sky130_fd_sc_hd__clkbuf_4
Xfanout148 _04938_ vssd1 vssd1 vccd1 vccd1 net148 sky130_fd_sc_hd__clkbuf_2
Xfanout159 net160 vssd1 vssd1 vccd1 vccd1 net159 sky130_fd_sc_hd__buf_2
XANTENNA__06231__A top.ramload\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07985_ top.DUT.register\[2\]\[31\] net744 net720 top.DUT.register\[19\]\[31\] vssd1
+ vssd1 vccd1 vccd1 _03124_ sky130_fd_sc_hd__a22o_1
X_09724_ _04172_ _04750_ _04751_ vssd1 vssd1 vccd1 vccd1 _04752_ sky130_fd_sc_hd__a21bo_2
X_06936_ top.DUT.register\[22\]\[21\] net650 _02074_ vssd1 vssd1 vccd1 vccd1 _02075_
+ sky130_fd_sc_hd__a21o_1
XANTENNA__09542__A _01764_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09655_ _04683_ _04693_ _04694_ _04695_ vssd1 vssd1 vccd1 vccd1 _04696_ sky130_fd_sc_hd__or4_1
X_06867_ _01983_ _02004_ vssd1 vssd1 vccd1 vccd1 _02006_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout551_A _01535_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08606_ net496 _03728_ vssd1 vssd1 vccd1 vccd1 _03729_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout649_A _01612_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_3_2_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_3_2_0_clk sky130_fd_sc_hd__clkbuf_8
X_09586_ top.pc\[29\] top.pc\[30\] _04597_ vssd1 vssd1 vccd1 vccd1 _04633_ sky130_fd_sc_hd__and3_1
X_06798_ top.DUT.register\[25\]\[17\] net456 net516 top.DUT.register\[7\]\[17\] vssd1
+ vssd1 vccd1 vccd1 _01937_ sky130_fd_sc_hd__a22o_1
XFILLER_0_194_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_167_627 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_139_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08537_ net885 top.pc\[12\] net696 _03663_ vssd1 vssd1 vccd1 vccd1 _03664_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_46_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout437_X net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_182_608 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13441__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07286__A2 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08468_ _02389_ _03596_ vssd1 vssd1 vccd1 vccd1 _03597_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_175_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11082__A3 net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_2501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06494__B1 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07419_ _02551_ _02553_ _02556_ _02557_ vssd1 vssd1 vccd1 vccd1 _02558_ sky130_fd_sc_hd__or4_1
XFILLER_0_162_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08399_ _03530_ vssd1 vssd1 vccd1 vccd1 _03531_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout604_X net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10627__S net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_708 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10430_ net146 net1779 net368 vssd1 vssd1 vccd1 vccd1 _00601_ sky130_fd_sc_hd__mux2_1
XANTENNA__08235__A1 net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_150_2701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_150_549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10361_ _04153_ _04947_ net399 vssd1 vssd1 vccd1 vccd1 _04981_ sky130_fd_sc_hd__and3_4
XFILLER_0_33_588 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12100_ _05981_ _05982_ vssd1 vssd1 vccd1 vccd1 _05983_ sky130_fd_sc_hd__nor2_1
X_13080_ clknet_leaf_126_clk _00672_ net929 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[18\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_238 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09717__A net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10292_ net1729 net154 net387 vssd1 vssd1 vccd1 vccd1 _00470_ sky130_fd_sc_hd__mux2_1
X_12031_ _05893_ _05899_ _05910_ _05911_ vssd1 vssd1 vccd1 vccd1 _05914_ sky130_fd_sc_hd__and4bb_1
XANTENNA__09196__C1 _01393_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08538__A2 net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10362__S net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09735__B2 top.a1.dataIn\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold180 top.ramaddr\[22\] vssd1 vssd1 vccd1 vccd1 net1296 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold191 top.DUT.register\[30\]\[17\] vssd1 vssd1 vccd1 vccd1 net1307 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07746__B1 net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_148_2663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout660 net662 vssd1 vssd1 vccd1 vccd1 net660 sky130_fd_sc_hd__clkbuf_8
XANTENNA__11982__A top.a1.dataIn\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout671 _01597_ vssd1 vssd1 vccd1 vccd1 net671 sky130_fd_sc_hd__buf_4
Xfanout682 _01547_ vssd1 vssd1 vccd1 vccd1 net682 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_70_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout693 _04049_ vssd1 vssd1 vccd1 vccd1 net693 sky130_fd_sc_hd__buf_6
X_12933_ clknet_leaf_33_clk _00525_ net1042 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[13\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_161_2863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11046__X _05045_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_201_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08710__A2 net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08068__A _02111_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12864_ clknet_leaf_80_clk _00456_ net991 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[11\]\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_200_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_205_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11058__B1 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11815_ _05667_ net131 _05696_ _05697_ vssd1 vssd1 vccd1 vccd1 _05698_ sky130_fd_sc_hd__a31oi_4
XFILLER_0_96_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12795_ clknet_leaf_124_clk _00387_ net923 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[9\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_139_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_194_3351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_194_3362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_200_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_32_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11746_ _01400_ _05624_ _05626_ _05627_ vssd1 vssd1 vccd1 vccd1 _05629_ sky130_fd_sc_hd__a211o_1
XANTENNA__07277__A2 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11677_ _05505_ _05526_ _05559_ vssd1 vssd1 vccd1 vccd1 _05560_ sky130_fd_sc_hd__o21ai_2
XANTENNA__10537__S net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_181_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07029__A2 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10628_ _04947_ _04952_ net400 vssd1 vssd1 vccd1 vccd1 _04992_ sky130_fd_sc_hd__nand3_4
X_13416_ clknet_leaf_27_clk _01008_ net1010 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[28\]\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08226__B2 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_181_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_180_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_77_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13347_ clknet_leaf_54_clk _00939_ net1037 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[26\]\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_10559_ net1817 net153 net356 vssd1 vssd1 vccd1 vccd1 _00726_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07985__B1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13278_ clknet_leaf_21_clk _00870_ net1034 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[24\]\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_90_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09726__A1 _04172_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12229_ top.lcd.cnt_20ms\[6\] _06053_ top.lcd.cnt_20ms\[7\] vssd1 vssd1 vccd1 vccd1
+ _06068_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_102_Left_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10272__S net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_208_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07770_ top.DUT.register\[9\]\[2\] net762 net635 top.DUT.register\[6\]\[2\] _02908_
+ vssd1 vssd1 vccd1 vccd1 _02909_ sky130_fd_sc_hd__a221o_1
X_06721_ top.DUT.register\[24\]\[25\] net643 net710 top.DUT.register\[11\]\[25\] _01859_
+ vssd1 vssd1 vccd1 vccd1 _01860_ sky130_fd_sc_hd__a221o_1
XFILLER_0_79_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_189_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13464__CLK clknet_leaf_128_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09440_ _04494_ _04495_ vssd1 vssd1 vccd1 vccd1 _04496_ sky130_fd_sc_hd__and2_1
X_06652_ top.DUT.register\[30\]\[26\] net582 net574 top.DUT.register\[23\]\[26\] vssd1
+ vssd1 vccd1 vccd1 _01791_ sky130_fd_sc_hd__a22o_1
XFILLER_0_189_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09081__B top.a1.instruction\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_68 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09371_ top.pc\[17\] _04420_ vssd1 vssd1 vccd1 vccd1 _04431_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_111_Left_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06583_ _01721_ vssd1 vssd1 vccd1 vccd1 _01722_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06992__Y _02131_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08322_ _03051_ _03456_ vssd1 vssd1 vccd1 vccd1 _03457_ sky130_fd_sc_hd__nand2_1
XFILLER_0_191_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_176_479 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08465__A1 net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07268__A2 net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08465__B2 _03594_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08253_ net317 _03389_ _03363_ vssd1 vssd1 vccd1 vccd1 _03390_ sky130_fd_sc_hd__a21o_1
XFILLER_0_144_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10447__S net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_119_2231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout132_A net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07204_ net895 _02332_ vssd1 vssd1 vccd1 vccd1 _02343_ sky130_fd_sc_hd__or2_2
XFILLER_0_144_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08184_ _01678_ net330 vssd1 vssd1 vccd1 vccd1 _03322_ sky130_fd_sc_hd__or2_1
XFILLER_0_6_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06226__A top.ramload\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_171_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10024__A1 net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08768__A2 net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07135_ top.DUT.register\[23\]\[11\] net571 net535 top.DUT.register\[19\]\[11\] vssd1
+ vssd1 vccd1 vccd1 _02274_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_132_2420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_132_2431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07976__B1 net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07609__X _02748_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_120_Left_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07066_ top.DUT.register\[17\]\[22\] net747 _02201_ _02204_ vssd1 vssd1 vccd1 vccd1
+ _02205_ sky130_fd_sc_hd__a211o_1
XFILLER_0_2_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07440__A2 net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout599_A _04965_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07728__B1 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09971__S net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout387_X net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout766_A net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10910__S net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07968_ top.DUT.register\[22\]\[31\] net576 net569 top.DUT.register\[6\]\[31\] vssd1
+ vssd1 vccd1 vccd1 _03107_ sky130_fd_sc_hd__a22o_1
XANTENNA__09272__A _02286_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06919_ top.DUT.register\[30\]\[21\] net582 net570 top.DUT.register\[6\]\[21\] _02057_
+ vssd1 vssd1 vccd1 vccd1 _02058_ sky130_fd_sc_hd__a221o_1
X_09707_ net827 _04238_ vssd1 vssd1 vccd1 vccd1 _04738_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout554_X net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07899_ top.DUT.register\[30\]\[1\] net581 net468 top.DUT.register\[9\]\[1\] _03037_
+ vssd1 vssd1 vccd1 vccd1 _03038_ sky130_fd_sc_hd__a221o_1
XANTENNA__11307__A _05123_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09638_ top.pad.keyCode\[1\] top.pad.keyCode\[0\] top.pad.keyCode\[3\] top.pad.keyCode\[2\]
+ vssd1 vssd1 vccd1 vccd1 _04680_ sky130_fd_sc_hd__or4b_2
XFILLER_0_69_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_143_2593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09569_ _04600_ _04601_ vssd1 vssd1 vccd1 vccd1 _04617_ sky130_fd_sc_hd__nand2b_1
XANTENNA_fanout721_X net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout819_X net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_468 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11600_ net234 _05476_ _05468_ _05470_ vssd1 vssd1 vccd1 vccd1 _05483_ sky130_fd_sc_hd__a211o_1
XFILLER_0_155_619 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12580_ clknet_leaf_37_clk _00172_ net1051 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[2\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_194_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07259__A2 net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_176_3081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_176_3092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08616__A _03121_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_455 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_182_438 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11531_ _05396_ _05398_ _05366_ _05373_ vssd1 vssd1 vccd1 vccd1 _05414_ sky130_fd_sc_hd__a211o_1
XANTENNA__10357__S net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11462_ _05287_ _05324_ _05317_ _05306_ vssd1 vssd1 vccd1 vccd1 _05345_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_20_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13201_ clknet_leaf_113_clk _00793_ net991 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[22\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_10413_ net1450 net226 net372 vssd1 vssd1 vccd1 vccd1 _00585_ sky130_fd_sc_hd__mux2_1
X_11393_ _05273_ _05274_ _05243_ _05272_ vssd1 vssd1 vccd1 vccd1 _05276_ sky130_fd_sc_hd__and4b_1
XTAP_TAPCELL_ROW_59_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07967__B1 net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13132_ clknet_leaf_48_clk _00724_ net1060 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[19\]\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_103_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10344_ net1487 net191 net379 vssd1 vssd1 vccd1 vccd1 _00520_ sky130_fd_sc_hd__mux2_1
XANTENNA__06423__X _01562_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09708__A1 top.a1.dataIn\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10092__S net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13063_ clknet_leaf_8_clk _00655_ net945 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[17\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_10275_ net1472 net214 net385 vssd1 vssd1 vccd1 vccd1 _00453_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_72_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12014_ _05889_ _05896_ vssd1 vssd1 vccd1 vccd1 _05897_ sky130_fd_sc_hd__nor2_1
XANTENNA__08931__A2 _03142_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13487__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10820__S net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout490 net491 vssd1 vssd1 vccd1 vccd1 net490 sky130_fd_sc_hd__buf_4
XANTENNA__09182__A net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_514 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12916_ clknet_leaf_55_clk _00508_ net1072 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[13\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07498__A2 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_186_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09910__A _04008_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_185_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12847_ clknet_leaf_32_clk _00439_ net1045 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[10\]\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_201_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_201_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_173_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08526__A net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12778_ clknet_leaf_115_clk _00370_ net957 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[8\]\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_83_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07430__A _02544_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10267__S net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11729_ _05567_ net163 _05581_ _05553_ vssd1 vssd1 vccd1 vccd1 _05612_ sky130_fd_sc_hd__a22o_2
XFILLER_0_9_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08245__B _03185_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_211_3605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_211_3616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07670__A2 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_211_3627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold905 top.DUT.register\[12\]\[27\] vssd1 vssd1 vccd1 vccd1 net2021 sky130_fd_sc_hd__dlygate4sd3_1
Xhold916 top.DUT.register\[14\]\[21\] vssd1 vssd1 vccd1 vccd1 net2032 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold927 top.DUT.register\[19\]\[15\] vssd1 vssd1 vccd1 vccd1 net2043 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_114_2150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07422__A2 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_114_2161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold938 top.DUT.register\[16\]\[31\] vssd1 vssd1 vccd1 vccd1 net2054 sky130_fd_sc_hd__dlygate4sd3_1
Xhold949 top.DUT.register\[2\]\[12\] vssd1 vssd1 vccd1 vccd1 net2065 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06630__B1 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08940_ net695 _04046_ _04047_ top.pc\[31\] net884 vssd1 vssd1 vccd1 vccd1 _04048_
+ sky130_fd_sc_hd__a32o_1
XANTENNA__12390__RESET_B net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_177_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08871_ _03096_ _03981_ vssd1 vssd1 vccd1 vccd1 _03982_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_209_3578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_208_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07822_ top.DUT.register\[14\]\[0\] net730 net635 top.DUT.register\[6\]\[0\] _02960_
+ vssd1 vssd1 vccd1 vccd1 _02961_ sky130_fd_sc_hd__a221o_1
XANTENNA__10730__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09092__A _01505_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07753_ top.DUT.register\[20\]\[3\] net566 net541 top.DUT.register\[8\]\[3\] vssd1
+ vssd1 vccd1 vccd1 _02892_ sky130_fd_sc_hd__a22o_1
XFILLER_0_193_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06704_ _01836_ _01838_ _01840_ _01842_ vssd1 vssd1 vccd1 vccd1 _01843_ sky130_fd_sc_hd__or4_1
XANTENNA__09332__C1 net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_177_711 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07684_ top.DUT.register\[4\]\[4\] net669 net732 top.DUT.register\[14\]\[4\] _02822_
+ vssd1 vssd1 vccd1 vccd1 _02823_ sky130_fd_sc_hd__a221o_1
XANTENNA__07489__A2 net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09423_ _04478_ _04479_ vssd1 vssd1 vccd1 vccd1 _04480_ sky130_fd_sc_hd__or2_1
X_06635_ top.DUT.register\[17\]\[27\] net748 net709 top.DUT.register\[15\]\[27\] vssd1
+ vssd1 vccd1 vccd1 _01774_ sky130_fd_sc_hd__a22o_1
XANTENNA__06697__B1 net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout347_A _04991_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_468 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1089_A net1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09354_ _04414_ vssd1 vssd1 vccd1 vccd1 _04415_ sky130_fd_sc_hd__inv_2
X_06566_ top.DUT.register\[12\]\[28\] net534 net529 top.DUT.register\[26\]\[28\] vssd1
+ vssd1 vccd1 vccd1 _01705_ sky130_fd_sc_hd__a22o_1
XFILLER_0_118_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08438__A1 net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08438__B2 _03334_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08305_ net305 _03196_ vssd1 vssd1 vccd1 vccd1 _03440_ sky130_fd_sc_hd__nor2_2
XFILLER_0_90_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09285_ _04346_ _04349_ vssd1 vssd1 vccd1 vccd1 _04350_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10177__S net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06497_ top.DUT.register\[13\]\[30\] net776 net748 top.DUT.register\[17\]\[30\] vssd1
+ vssd1 vccd1 vccd1 _01636_ sky130_fd_sc_hd__a22o_1
XFILLER_0_19_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout514_A _01559_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout135_X net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08236_ net298 _03372_ _03367_ vssd1 vssd1 vccd1 vccd1 _03373_ sky130_fd_sc_hd__o21ai_1
XANTENNA__09966__S net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_145_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08167_ _03303_ _03304_ vssd1 vssd1 vccd1 vccd1 _03305_ sky130_fd_sc_hd__nand2_1
XFILLER_0_30_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10905__S net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07118_ top.DUT.register\[20\]\[16\] net664 net771 top.DUT.register\[10\]\[16\] _02252_
+ vssd1 vssd1 vccd1 vccd1 _02257_ sky130_fd_sc_hd__a221o_1
X_08098_ _03227_ _03229_ _03236_ net311 net285 vssd1 vssd1 vccd1 vccd1 _03237_ sky130_fd_sc_hd__o221a_1
XANTENNA__07413__A2 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout883_A net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_189_Right_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06621__B1 net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07049_ _02181_ _02183_ _02185_ _02187_ vssd1 vssd1 vccd1 vccd1 _02188_ sky130_fd_sc_hd__or4_4
XFILLER_0_140_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_54_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10060_ net1653 net210 net617 vssd1 vssd1 vccd1 vccd1 _00262_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_54_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout671_X net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout769_X net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10640__S net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_2622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07515__A _02633_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_207_Left_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_3_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08677__A1 net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_178_3110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13750_ clknet_leaf_99_clk _01321_ vssd1 vssd1 vccd1 vccd1 top.lcd.cnt_20ms\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_10962_ net888 net784 _05004_ net844 vssd1 vssd1 vccd1 vccd1 _05005_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_178_3121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09874__B1 net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06688__B1 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12701_ clknet_leaf_118_clk _00293_ net955 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[6\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10893_ net1667 net252 net478 vssd1 vssd1 vccd1 vccd1 _01054_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13681_ clknet_leaf_75_clk _01257_ net1079 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[15\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_155_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08429__A1 net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_191_3310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12632_ clknet_leaf_127_clk _00224_ net929 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[4\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_155_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12563_ clknet_leaf_120_clk _00155_ net932 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[2\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10087__S net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_202_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_182_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11514_ _05386_ _05392_ vssd1 vssd1 vccd1 vccd1 _05397_ sky130_fd_sc_hd__or2_1
XFILLER_0_53_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09729__X _04757_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_156_2784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07652__A2 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12494_ clknet_leaf_84_clk _00086_ net994 vssd1 vssd1 vccd1 vccd1 top.pc\[6\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_124_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_22_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06860__B1 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11445_ _05326_ _05327_ vssd1 vssd1 vccd1 vccd1 _05328_ sky130_fd_sc_hd__or2_1
XANTENNA__12727__CLK clknet_leaf_128_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10815__S net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_491 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_519 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11376_ _05257_ _05258_ _05223_ _05251_ vssd1 vssd1 vccd1 vccd1 _05259_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_33_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08601__A1 net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_189_3283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13695__Q net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08601__B2 _03724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06612__B1 net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_156_Right_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13115_ clknet_leaf_127_clk _00707_ net929 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[19\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_10327_ net141 net1872 net382 vssd1 vssd1 vccd1 vccd1 _00504_ sky130_fd_sc_hd__mux2_1
X_13046_ clknet_leaf_3_clk _00638_ net940 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[17\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_10258_ net157 net1324 net391 vssd1 vssd1 vccd1 vccd1 _00437_ sky130_fd_sc_hd__mux2_1
XANTENNA__12877__CLK clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10550__S net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10189_ _04968_ vssd1 vssd1 vccd1 vccd1 _04969_ sky130_fd_sc_hd__inv_2
XFILLER_0_206_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_206_656 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09343__C _04403_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_205_155 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08117__B1 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06391__A2 net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_205_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_178_519 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_85_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09062__D _03655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06679__B1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_186_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06420_ net685 _01521_ _01527_ vssd1 vssd1 vccd1 vccd1 _01559_ sky130_fd_sc_hd__and3_4
XFILLER_0_29_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_146_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_174_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_146_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06351_ top.pad.button_control.r_counter\[10\] top.pad.button_control.r_counter\[9\]
+ top.pad.button_control.r_counter\[7\] top.pad.button_control.r_counter\[5\] vssd1
+ vssd1 vccd1 vccd1 _01491_ sky130_fd_sc_hd__nand4_1
XFILLER_0_8_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09786__S net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09070_ _01475_ _02346_ _04144_ net829 vssd1 vssd1 vccd1 vccd1 _04145_ sky130_fd_sc_hd__o211a_1
X_06282_ _01404_ top.lcd.cnt_500hz\[13\] top.lcd.cnt_500hz\[12\] _01444_ vssd1 vssd1
+ vccd1 vccd1 _01445_ sky130_fd_sc_hd__or4_1
XFILLER_0_126_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07643__A2 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08021_ _01501_ _03151_ vssd1 vssd1 vccd1 vccd1 _03160_ sky130_fd_sc_hd__or2_2
XANTENNA__06851__B1 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_812 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10725__S net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold702 top.DUT.register\[20\]\[22\] vssd1 vssd1 vccd1 vccd1 net1818 sky130_fd_sc_hd__dlygate4sd3_1
Xhold713 top.DUT.register\[30\]\[2\] vssd1 vssd1 vccd1 vccd1 net1829 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_4_1__f_clk_A clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold724 top.DUT.register\[26\]\[16\] vssd1 vssd1 vccd1 vccd1 net1840 sky130_fd_sc_hd__dlygate4sd3_1
Xhold735 top.DUT.register\[22\]\[27\] vssd1 vssd1 vccd1 vccd1 net1851 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_96_1886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold746 top.DUT.register\[30\]\[0\] vssd1 vssd1 vccd1 vccd1 net1862 sky130_fd_sc_hd__dlygate4sd3_1
Xhold757 top.DUT.register\[2\]\[28\] vssd1 vssd1 vccd1 vccd1 net1873 sky130_fd_sc_hd__dlygate4sd3_1
Xhold768 top.DUT.register\[27\]\[13\] vssd1 vssd1 vccd1 vccd1 net1884 sky130_fd_sc_hd__dlygate4sd3_1
X_09972_ net1964 net162 net630 vssd1 vssd1 vccd1 vccd1 _00180_ sky130_fd_sc_hd__mux2_1
Xhold779 top.ramaddr\[10\] vssd1 vssd1 vccd1 vccd1 net1895 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_123_Right_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06223__B net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08923_ _01659_ _04013_ _01657_ vssd1 vssd1 vccd1 vccd1 _04031_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_41_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout297_A net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10460__S net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08854_ _03095_ _03965_ vssd1 vssd1 vccd1 vccd1 _03966_ sky130_fd_sc_hd__nor2_1
XANTENNA__09534__B _04577_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07805_ _02934_ _02943_ vssd1 vssd1 vccd1 vccd1 _02944_ sky130_fd_sc_hd__or2_4
XFILLER_0_98_108 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_2352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08785_ _03822_ _03899_ net308 vssd1 vssd1 vccd1 vccd1 _03900_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout464_A net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07736_ top.DUT.register\[21\]\[3\] net657 net649 top.DUT.register\[22\]\[3\] _02869_
+ vssd1 vssd1 vccd1 vccd1 _02875_ sky130_fd_sc_hd__a221o_1
XFILLER_0_197_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08659__A1 _02048_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_2541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07667_ top.a1.instruction\[25\] _01508_ net411 vssd1 vssd1 vccd1 vccd1 _02806_ sky130_fd_sc_hd__a21o_1
XFILLER_0_94_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_140_2552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_211_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout631_A _04714_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_177_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout729_A _01628_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06618_ top.DUT.register\[16\]\[27\] net544 net529 top.DUT.register\[26\]\[27\] _01756_
+ vssd1 vssd1 vccd1 vccd1 _01757_ sky130_fd_sc_hd__a221o_1
XFILLER_0_165_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09406_ top.pc\[19\] _04453_ vssd1 vssd1 vccd1 vccd1 _04464_ sky130_fd_sc_hd__and2_1
XFILLER_0_137_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08166__A _02198_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07598_ top.DUT.register\[4\]\[6\] net667 net663 top.DUT.register\[20\]\[6\] _02732_
+ vssd1 vssd1 vccd1 vccd1 _02737_ sky130_fd_sc_hd__a221o_1
XFILLER_0_94_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_165_758 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06549_ _01681_ _01685_ _01686_ _01687_ vssd1 vssd1 vccd1 vccd1 _01688_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_173_3040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09337_ _04380_ _04381_ _04382_ vssd1 vssd1 vccd1 vccd1 _04399_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout517_X net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09696__S net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09268_ _04321_ _04322_ _04319_ vssd1 vssd1 vccd1 vccd1 _04334_ sky130_fd_sc_hd__o21ai_1
X_08219_ _03246_ _03250_ net291 vssd1 vssd1 vccd1 vccd1 _03356_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06842__B1 net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10635__S net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09199_ top.pc\[6\] _04236_ top.pc\[7\] vssd1 vssd1 vccd1 vccd1 _04269_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_105_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_688 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11230_ top.lcd.nextState\[3\] net879 _05122_ vssd1 vssd1 vccd1 vccd1 _05123_ sky130_fd_sc_hd__and3_2
XANTENNA_fanout886_X net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11194__A2 net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_686 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11161_ top.a1.row1\[57\] _05089_ _05085_ vssd1 vssd1 vccd1 vccd1 _01228_ sky130_fd_sc_hd__mux2_1
X_10112_ _04156_ _04709_ _04952_ vssd1 vssd1 vccd1 vccd1 _04956_ sky130_fd_sc_hd__or3b_4
XTAP_TAPCELL_ROW_8_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11092_ net908 net1462 net863 _05051_ vssd1 vssd1 vccd1 vccd1 _01197_ sky130_fd_sc_hd__a31o_1
X_10043_ net2208 net152 net621 vssd1 vssd1 vccd1 vccd1 _00246_ sky130_fd_sc_hd__mux2_1
XANTENNA__10370__S net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09444__B _04499_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08898__A1 net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold40 top.a1.dataInTemp\[8\] vssd1 vssd1 vccd1 vccd1 net1156 sky130_fd_sc_hd__dlygate4sd3_1
Xhold51 _01180_ vssd1 vssd1 vccd1 vccd1 net1167 sky130_fd_sc_hd__dlygate4sd3_1
Xhold62 top.ramload\[16\] vssd1 vssd1 vccd1 vccd1 net1178 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07245__A _02383_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input25_A DAT_I[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold73 _01175_ vssd1 vssd1 vccd1 vccd1 net1189 sky130_fd_sc_hd__dlygate4sd3_1
Xhold84 _01173_ vssd1 vssd1 vccd1 vccd1 net1200 sky130_fd_sc_hd__dlygate4sd3_1
Xhold95 _01162_ vssd1 vssd1 vccd1 vccd1 net1211 sky130_fd_sc_hd__dlygate4sd3_1
X_13802_ clknet_leaf_71_clk _01371_ net1086 vssd1 vssd1 vccd1 vccd1 top.pad.keyCode\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_98_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_203_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11994_ _05804_ _05875_ vssd1 vssd1 vccd1 vccd1 _05877_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_58_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09460__A _02198_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_12__f_clk_A clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13733_ clknet_leaf_94_clk _01304_ vssd1 vssd1 vccd1 vccd1 top.a1.dataInTemp\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_67_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10945_ net2124 net169 _04960_ vssd1 vssd1 vccd1 vccd1 _01106_ sky130_fd_sc_hd__mux2_1
XFILLER_0_168_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_158_2813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13664_ clknet_leaf_91_clk _01240_ net996 vssd1 vssd1 vccd1 vccd1 top.a1.row1\[114\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06295__S net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08076__A _01983_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10876_ net201 net2026 net597 vssd1 vssd1 vccd1 vccd1 _01037_ sky130_fd_sc_hd__mux2_1
XANTENNA__07873__A2 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_80_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12615_ clknet_leaf_5_clk _00207_ net937 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[3\]\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13595_ clknet_leaf_65_clk net1174 net1095 vssd1 vssd1 vccd1 vccd1 net87 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_183_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09459__X _04514_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07086__B1 net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07625__A2 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12546_ clknet_leaf_10_clk _00138_ net948 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[1\]\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_164_791 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06833__B1 net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10545__S net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12477_ clknet_leaf_65_clk _00072_ net1094 vssd1 vssd1 vccd1 vccd1 top.ramstore\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_34_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_4 top.a1.dataIn\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11230__A top.lcd.nextState\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11428_ _05241_ _05268_ _05243_ vssd1 vssd1 vccd1 vccd1 _05311_ sky130_fd_sc_hd__a21o_1
XFILLER_0_158_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11185__A2 net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11359_ _05241_ vssd1 vssd1 vccd1 vccd1 _05242_ sky130_fd_sc_hd__inv_2
XANTENNA__09057__D _03881_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_169_2975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_169_2986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13029_ clknet_leaf_35_clk _00621_ net1041 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[16\]\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10280__S net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_206_3537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08889__A1 net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1060 net1061 vssd1 vssd1 vccd1 vccd1 net1060 sky130_fd_sc_hd__buf_2
Xfanout1071 net1098 vssd1 vssd1 vccd1 vccd1 net1071 sky130_fd_sc_hd__buf_4
XANTENNA__09922__X _04929_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_6_clk_A clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1082 net1083 vssd1 vssd1 vccd1 vccd1 net1082 sky130_fd_sc_hd__clkbuf_2
Xfanout1093 net1096 vssd1 vssd1 vccd1 vccd1 net1093 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_179_806 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_109_2082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08570_ _03694_ vssd1 vssd1 vccd1 vccd1 _03695_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10012__C top.a1.instruction\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07521_ top.DUT.register\[6\]\[7\] net567 net531 top.DUT.register\[12\]\[7\] vssd1
+ vssd1 vccd1 vccd1 _02660_ sky130_fd_sc_hd__a22o_1
XFILLER_0_202_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_122_2271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07452_ top.DUT.register\[15\]\[15\] net707 net699 top.DUT.register\[31\]\[15\] vssd1
+ vssd1 vccd1 vccd1 _02591_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_122_2282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07864__A2 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06403_ net683 _01527_ _01533_ vssd1 vssd1 vccd1 vccd1 _01542_ sky130_fd_sc_hd__and3_4
X_07383_ _02502_ _02521_ net825 vssd1 vssd1 vccd1 vccd1 _02522_ sky130_fd_sc_hd__mux2_2
X_09122_ _04190_ _04194_ _04196_ vssd1 vssd1 vccd1 vccd1 _04197_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_8_179 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06334_ top.d_ready _01480_ _01476_ top.ru.state\[0\] vssd1 vssd1 vccd1 vccd1 top.ru.next_write_i
+ sky130_fd_sc_hd__and4bb_1
XANTENNA__07077__B1 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07616__A2 net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_1915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_199_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09053_ _03560_ _03585_ _03610_ _03626_ vssd1 vssd1 vccd1 vccd1 _04128_ sky130_fd_sc_hd__or4_1
XFILLER_0_115_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06265_ top.ramload\[26\] net853 vssd1 vssd1 vccd1 vccd1 top.ru.next_FetchedData\[26\]
+ sky130_fd_sc_hd__and2_1
XANTENNA__10455__S net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08004_ _03122_ _03142_ vssd1 vssd1 vccd1 vccd1 _03143_ sky130_fd_sc_hd__nor2_1
XFILLER_0_130_603 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold510 top.DUT.register\[24\]\[8\] vssd1 vssd1 vccd1 vccd1 net1626 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08026__C1 _03162_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06196_ wb.curr_state\[2\] wb.curr_state\[1\] vssd1 vssd1 vccd1 vccd1 _01427_ sky130_fd_sc_hd__nor2_4
XANTENNA__06234__A top.ramload\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold521 top.DUT.register\[10\]\[13\] vssd1 vssd1 vccd1 vccd1 net1637 sky130_fd_sc_hd__dlygate4sd3_1
Xhold532 top.DUT.register\[20\]\[24\] vssd1 vssd1 vccd1 vccd1 net1648 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold543 top.DUT.register\[20\]\[19\] vssd1 vssd1 vccd1 vccd1 net1659 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold554 top.DUT.register\[28\]\[1\] vssd1 vssd1 vccd1 vccd1 net1670 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold565 top.DUT.register\[7\]\[17\] vssd1 vssd1 vccd1 vccd1 net1681 sky130_fd_sc_hd__dlygate4sd3_1
Xhold576 top.DUT.register\[5\]\[21\] vssd1 vssd1 vccd1 vccd1 net1692 sky130_fd_sc_hd__dlygate4sd3_1
Xhold587 top.ramaddr\[20\] vssd1 vssd1 vccd1 vccd1 net1703 sky130_fd_sc_hd__dlygate4sd3_1
Xhold598 top.DUT.register\[6\]\[18\] vssd1 vssd1 vccd1 vccd1 net1714 sky130_fd_sc_hd__dlygate4sd3_1
X_09955_ net1683 net229 net627 vssd1 vssd1 vccd1 vccd1 _00163_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout581_A _01514_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout679_A _01547_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08906_ net497 _04014_ vssd1 vssd1 vccd1 vccd1 _04015_ sky130_fd_sc_hd__nor2_1
X_09886_ net2075 net165 net634 vssd1 vssd1 vccd1 vccd1 _00147_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout1007_X net1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07001__B1 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09832__X _04847_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09541__A2 _01763_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08837_ net497 _03936_ _03949_ vssd1 vssd1 vccd1 vccd1 _03950_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout467_X net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout846_A net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08768_ _02134_ net433 net501 _02135_ _03883_ vssd1 vssd1 vccd1 vccd1 _03884_ sky130_fd_sc_hd__a221o_1
XANTENNA__09280__A top.pc\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07719_ _02857_ vssd1 vssd1 vccd1 vccd1 _02858_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout634_X net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08699_ net321 _03441_ vssd1 vssd1 vccd1 vccd1 _03818_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_49_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10730_ net1447 net265 net418 vssd1 vssd1 vccd1 vccd1 _00891_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_24_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10661_ _04155_ _04952_ net399 vssd1 vssd1 vccd1 vccd1 _04993_ sky130_fd_sc_hd__and3_4
XFILLER_0_94_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12493__RESET_B net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12400_ clknet_leaf_103_clk top.ru.next_FetchedInstr\[12\] net976 vssd1 vssd1 vccd1
+ vccd1 top.a1.instruction\[12\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_62_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07068__B1 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13380_ clknet_leaf_36_clk _00972_ net1049 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[27\]\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_180_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10592_ top.DUT.register\[20\]\[29\] net154 net352 vssd1 vssd1 vccd1 vccd1 _00758_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__07607__A2 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12331_ top.pad.button_control.r_counter\[11\] top.pad.button_control.r_counter\[10\]
+ _06127_ vssd1 vssd1 vccd1 vccd1 _06131_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_153_2743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10365__S net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12262_ top.lcd.cnt_500hz\[1\] top.lcd.cnt_500hz\[0\] top.lcd.cnt_500hz\[2\] vssd1
+ vssd1 vccd1 vccd1 _06088_ sky130_fd_sc_hd__a21o_1
XANTENNA__08911__X _04020_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11213_ net1979 net472 _04668_ vssd1 vssd1 vccd1 vccd1 _01257_ sky130_fd_sc_hd__a21o_1
XANTENNA__08568__B1 _03691_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_186_3231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_186_3242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12193_ net1127 _06045_ net688 vssd1 vssd1 vccd1 vccd1 _01300_ sky130_fd_sc_hd__mux2_1
Xoutput41 net41 vssd1 vssd1 vccd1 vccd1 ADR_O[10] sky130_fd_sc_hd__buf_2
Xoutput52 net52 vssd1 vssd1 vccd1 vccd1 ADR_O[20] sky130_fd_sc_hd__buf_2
XANTENNA__08997__C _03606_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11144_ net907 net1295 net862 _05077_ vssd1 vssd1 vccd1 vccd1 _01223_ sky130_fd_sc_hd__a31o_1
Xoutput63 net63 vssd1 vssd1 vccd1 vccd1 ADR_O[30] sky130_fd_sc_hd__buf_2
Xoutput74 net74 vssd1 vssd1 vccd1 vccd1 DAT_O[10] sky130_fd_sc_hd__buf_2
Xoutput85 net85 vssd1 vssd1 vccd1 vccd1 DAT_O[20] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_207_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput96 net96 vssd1 vssd1 vccd1 vccd1 DAT_O[30] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_101_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11075_ net91 net872 net836 net1229 vssd1 vssd1 vccd1 vccd1 _01186_ sky130_fd_sc_hd__a22o_1
XANTENNA__06150__Y _01393_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10026_ net2229 net211 net619 vssd1 vssd1 vccd1 vccd1 _00229_ sky130_fd_sc_hd__mux2_1
XANTENNA_input28_X net28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12915__CLK clknet_leaf_120_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09190__A _02723_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_201_3456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_201_3467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11977_ _05795_ _05833_ _05829_ vssd1 vssd1 vccd1 vccd1 _05860_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_58_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11225__A top.lcd.nextState\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13716_ clknet_leaf_97_clk _01287_ net984 vssd1 vssd1 vccd1 vccd1 top.a1.row2\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07846__A2 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10928_ net2036 net237 net593 vssd1 vssd1 vccd1 vccd1 _01089_ sky130_fd_sc_hd__mux2_1
XFILLER_0_168_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09048__A1 net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13647_ clknet_leaf_94_clk net873 net983 vssd1 vssd1 vccd1 vccd1 top.ru.state\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10859_ net260 net1719 net596 vssd1 vssd1 vccd1 vccd1 _01020_ sky130_fd_sc_hd__mux2_1
XFILLER_0_171_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_144_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_167_Left_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13578_ clknet_leaf_89_clk net1215 net1003 vssd1 vssd1 vccd1 vccd1 net100 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10275__S net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12529_ clknet_leaf_112_clk _00121_ net988 vssd1 vssd1 vccd1 vccd1 top.DUT.register\[1\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_112_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_10_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_1834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_1845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07231__B1 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout308 net310 vssd1 vssd1 vccd1 vccd1 net308 sky130_fd_sc_hd__clkbuf_4
Xfanout319 _02830_ vssd1 vssd1 vccd1 vccd1 net319 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_185_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06585__A2 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06952_ _02069_ _02089_ vssd1 vssd1 vccd1 vccd1 _02091_ sky130_fd_sc_hd__nor2_1
XANTENNA__09084__B top.a1.instruction\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09740_ top.pc\[11\] net799 _04754_ _04764_ vssd1 vssd1 vccd1 vccd1 _04765_ sky130_fd_sc_hd__a211o_1
.ends

