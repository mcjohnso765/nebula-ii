* NGSPICE file created from team_10.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_2 abstract view
.subckt sky130_fd_sc_hd__dfstp_2 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinvlp_4 abstract view
.subckt sky130_fd_sc_hd__clkinvlp_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_1 abstract view
.subckt sky130_fd_sc_hd__clkinv_1 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_12 abstract view
.subckt sky130_fd_sc_hd__inv_12 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_8 abstract view
.subckt sky130_fd_sc_hd__clkinv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_8 abstract view
.subckt sky130_fd_sc_hd__inv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__bufinv_16 abstract view
.subckt sky130_fd_sc_hd__bufinv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_16 abstract view
.subckt sky130_fd_sc_hd__inv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_2 abstract view
.subckt sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_4 abstract view
.subckt sky130_fd_sc_hd__and3b_4 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_2 abstract view
.subckt sky130_fd_sc_hd__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_2 abstract view
.subckt sky130_fd_sc_hd__a2111oi_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_2 abstract view
.subckt sky130_fd_sc_hd__o2111ai_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_2 abstract view
.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

.subckt team_10 clk en gpio_in[0] gpio_in[10] gpio_in[11] gpio_in[12] gpio_in[13]
+ gpio_in[14] gpio_in[15] gpio_in[16] gpio_in[17] gpio_in[18] gpio_in[19] gpio_in[1]
+ gpio_in[20] gpio_in[21] gpio_in[22] gpio_in[23] gpio_in[24] gpio_in[25] gpio_in[26]
+ gpio_in[27] gpio_in[28] gpio_in[29] gpio_in[2] gpio_in[30] gpio_in[31] gpio_in[32]
+ gpio_in[33] gpio_in[3] gpio_in[4] gpio_in[5] gpio_in[6] gpio_in[7] gpio_in[8] gpio_in[9]
+ gpio_oeb[0] gpio_oeb[10] gpio_oeb[11] gpio_oeb[12] gpio_oeb[13] gpio_oeb[14] gpio_oeb[15]
+ gpio_oeb[16] gpio_oeb[17] gpio_oeb[18] gpio_oeb[19] gpio_oeb[1] gpio_oeb[20] gpio_oeb[21]
+ gpio_oeb[22] gpio_oeb[23] gpio_oeb[24] gpio_oeb[25] gpio_oeb[26] gpio_oeb[27] gpio_oeb[28]
+ gpio_oeb[29] gpio_oeb[2] gpio_oeb[30] gpio_oeb[31] gpio_oeb[32] gpio_oeb[33] gpio_oeb[3]
+ gpio_oeb[4] gpio_oeb[5] gpio_oeb[6] gpio_oeb[7] gpio_oeb[8] gpio_oeb[9] gpio_out[0]
+ gpio_out[10] gpio_out[11] gpio_out[12] gpio_out[13] gpio_out[14] gpio_out[15] gpio_out[16]
+ gpio_out[17] gpio_out[18] gpio_out[19] gpio_out[1] gpio_out[20] gpio_out[21] gpio_out[22]
+ gpio_out[23] gpio_out[24] gpio_out[25] gpio_out[26] gpio_out[27] gpio_out[28] gpio_out[29]
+ gpio_out[2] gpio_out[30] gpio_out[31] gpio_out[32] gpio_out[33] gpio_out[3] gpio_out[4]
+ gpio_out[5] gpio_out[6] gpio_out[7] gpio_out[8] gpio_out[9] nrst vccd1 vssd1
XFILLER_0_94_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3155_ clknet_leaf_16_clk _0131_ net222 vssd1 vssd1 vccd1 vccd1 keypadplayer.scan_col\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__1911__X _0764_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3086_ clknet_leaf_18_clk _0076_ net219 vssd1 vssd1 vccd1 vccd1 message_reg.msg\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2106_ hostdisp.curr_word\[34\] net99 _0855_ gamelogic.letter\[2\] vssd1 vssd1 vccd1
+ vccd1 hostdisp.next_curr_word\[34\] sky130_fd_sc_hd__o22a_1
X_2037_ net143 net91 net76 net458 vssd1 vssd1 vccd1 vccd1 hostdisp.next_curr_guesses\[43\]
+ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout162_A net165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_94 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2939_ net482 net88 net65 net460 vssd1 vssd1 vccd1 vccd1 _0306_ sky130_fd_sc_hd__a22o_1
XFILLER_0_150_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2954__A1 host_message_reg.setLetter\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2954__B2 gamelogic.setWord\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_157_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2706__A1 gamelogic.letter\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout75_A _0830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_169_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_169_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3282__CLK clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2642__B1 _0360_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1996__A2 net92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_180_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_180 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_171_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2633__B1 _1086_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_155 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2724_ gamelogic.indexCorrect\[0\] _1236_ _1286_ _0921_ vssd1 vssd1 vccd1 vccd1 _0196_
+ sky130_fd_sc_hd__a22o_1
X_2655_ dispFSM.guesses\[63\] net118 net108 dispFSM.msg\[7\] vssd1 vssd1 vccd1 vccd1
+ _1226_ sky130_fd_sc_hd__a22o_1
XFILLER_0_89_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1606_ _0539_ _0540_ vssd1 vssd1 vccd1 vccd1 _0541_ sky130_fd_sc_hd__nor2_1
XFILLER_0_120_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2586_ _0360_ _1147_ _1153_ _1160_ vssd1 vssd1 vccd1 vccd1 _1161_ sky130_fd_sc_hd__a211o_1
X_1537_ _0419_ net128 keypadFSMPlayer.prev_key\[5\] vssd1 vssd1 vccd1 vccd1 _0485_
+ sky130_fd_sc_hd__a21oi_1
Xfanout116 _0732_ vssd1 vssd1 vccd1 vccd1 net116 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_129_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout105 _1081_ vssd1 vssd1 vccd1 vccd1 net105 sky130_fd_sc_hd__buf_4
Xfanout127 _0630_ vssd1 vssd1 vccd1 vccd1 net127 sky130_fd_sc_hd__clkbuf_4
Xfanout138 lcdPlayer.nextState\[1\] vssd1 vssd1 vccd1 vccd1 net138 sky130_fd_sc_hd__buf_2
X_1468_ _0418_ _0419_ vssd1 vssd1 vccd1 vccd1 _0420_ sky130_fd_sc_hd__nor2_1
XFILLER_0_129_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout149 uart_receiver.bit_index\[1\] vssd1 vssd1 vccd1 vccd1 net149 sky130_fd_sc_hd__clkbuf_2
XANTENNA__3342__Q gamelogic.letter\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3207_ clknet_leaf_27_clk _0183_ vssd1 vssd1 vccd1 vccd1 lcdPlayer.currentState\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_3138_ clknet_leaf_26_clk _0114_ vssd1 vssd1 vccd1 vccd1 lcdPlayer.cnt_20ms\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_107_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3069_ clknet_leaf_15_clk _0062_ _0031_ vssd1 vssd1 vccd1 vccd1 dispFSM.msg\[4\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_0_54_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout165_X net165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_159_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_92 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_115_Left_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold170 dispFSM.guesses\[29\] vssd1 vssd1 vccd1 vccd1 net434 sky130_fd_sc_hd__dlygate4sd3_1
Xhold181 _0290_ vssd1 vssd1 vccd1 vccd1 net445 sky130_fd_sc_hd__dlygate4sd3_1
Xhold192 lcdPlayer.cnt_20ms\[7\] vssd1 vssd1 vccd1 vccd1 net456 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_18_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_31_clk_A clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3602__236 vssd1 vssd1 vccd1 vccd1 _3602__236/HI net236 sky130_fd_sc_hd__conb_1
XPHY_EDGE_ROW_124_Left_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1711__B net100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2615__A0 hostdisp.bottom\[101\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_330 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2823__A net100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_177_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_119 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2091__B2 net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_180_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_133_Left_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3178__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2440_ net130 host_message_reg.setLetter\[2\] hostdisp.curr_word\[18\] net73 net71
+ vssd1 vssd1 vccd1 vccd1 _1042_ sky130_fd_sc_hd__a221o_1
XFILLER_0_11_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_166_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2371_ lcdPlayer.cnt_20ms\[10\] _1004_ net167 vssd1 vssd1 vccd1 vccd1 _1006_ sky130_fd_sc_hd__o21ai_1
XANTENNA__3223__RESET_B net223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3162__Q hostdisp.top\[46\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_79 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_142_Left_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2854__A0 gamelogic.letter\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2606__B1 net108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2082__B2 gamelogic.letter\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_151_Left_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout125_A net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2707_ net143 gamelogic.setWord\[19\] vssd1 vssd1 vccd1 vccd1 _1271_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_154_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2638_ hostdisp.bottom\[54\] net114 _1098_ hostdisp.top\[46\] vssd1 vssd1 vccd1 vccd1
+ _1210_ sky130_fd_sc_hd__a22o_1
X_2569_ hostdisp.bottom\[51\] net114 _1095_ hostdisp.top\[75\] vssd1 vssd1 vccd1 vccd1
+ _1144_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_160_Left_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_7_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_165_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_137_Right_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3470__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_172_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2128__A2 net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_142_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1940_ _0765_ _0768_ vssd1 vssd1 vccd1 vccd1 _0786_ sky130_fd_sc_hd__nor2_1
X_1871_ uart_transmitter.clk_count\[0\] net290 _0733_ vssd1 vssd1 vccd1 vccd1 uart_transmitter.next_clk_count\[1\]
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_16_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_104_Right_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3610_ gamelogic.red vssd1 vssd1 vccd1 vccd1 net35 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_141_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3541_ clknet_leaf_14_clk hostdisp.next_curr_guesses\[23\] net206 vssd1 vssd1 vccd1
+ vccd1 hostdisp.curr_guesses\[23\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_12_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3472_ clknet_leaf_1_clk _0350_ net175 vssd1 vssd1 vccd1 vccd1 gamelogic.setWord\[34\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_10_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2423_ hostdisp.curr_word\[8\] _0830_ net70 net368 _1034_ vssd1 vssd1 vccd1 vccd1
+ _0140_ sky130_fd_sc_hd__a221o_1
X_2354_ net167 _0946_ _0995_ _0955_ vssd1 vssd1 vccd1 vccd1 _0110_ sky130_fd_sc_hd__a31o_1
X_2285_ _0953_ vssd1 vssd1 vccd1 vccd1 _0954_ sky130_fd_sc_hd__inv_2
XFILLER_0_193_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3343__CLK clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2055__B2 net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_191_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_144_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3493__CLK clknet_leaf_30_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3067__Q dispFSM.msg\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1807__A _0693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input2_X net2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2597__A2 _1072_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_174_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_94_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2521__A2 _1095_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_59 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3366__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2070_ hostdisp.curr_word\[13\] net96 _0841_ net141 vssd1 vssd1 vccd1 vccd1 hostdisp.next_curr_word\[13\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_163_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_146_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2972_ gamelogic.setWord\[11\] net51 net47 gamelogic.setWord\[19\] vssd1 vssd1 vccd1
+ vccd1 _0335_ sky130_fd_sc_hd__o22a_1
XANTENNA__2037__A1 net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2588__A2 net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1923_ _0773_ vssd1 vssd1 vccd1 vccd1 _0187_ sky130_fd_sc_hd__inv_2
X_3615__246 vssd1 vssd1 vccd1 vccd1 _3615__246/HI net246 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_192_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1854_ clock_div.count\[25\] _0725_ vssd1 vssd1 vccd1 vccd1 _0727_ sky130_fd_sc_hd__and2_1
XFILLER_0_21_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1627__A net3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1785_ clock_div.count\[23\] clock_div.count\[22\] clock_div.count\[25\] clock_div.count\[24\]
+ vssd1 vssd1 vccd1 vccd1 _0683_ sky130_fd_sc_hd__or4_1
XFILLER_0_12_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3524_ clknet_leaf_5_clk hostdisp.next_curr_guesses\[6\] net193 vssd1 vssd1 vccd1
+ vccd1 hostdisp.curr_guesses\[6\] sky130_fd_sc_hd__dfstp_1
XFILLER_0_12_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_151_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3455_ clknet_leaf_7_clk _0333_ net195 vssd1 vssd1 vccd1 vccd1 gamelogic.setWord\[17\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_12_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2406_ _0361_ _0430_ vssd1 vssd1 vccd1 vccd1 _1028_ sky130_fd_sc_hd__nor2_1
X_3386_ clknet_leaf_25_clk _0275_ net183 vssd1 vssd1 vccd1 vccd1 dispFSM.guesses\[40\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_110_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout192_A net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2337_ lcdPlayer.cnt_500hz\[18\] _0984_ lcdPlayer.cnt_500hz\[19\] vssd1 vssd1 vccd1
+ vccd1 _0987_ sky130_fd_sc_hd__a21o_1
XANTENNA__2512__A2 _1084_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2268_ dispFSM.msg\[2\] _0941_ _0942_ net302 vssd1 vssd1 vccd1 vccd1 _0077_ sky130_fd_sc_hd__a22o_1
XFILLER_0_98_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_162_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2199_ net129 gamelogic.setWord\[34\] vssd1 vssd1 vccd1 vccd1 _0902_ sky130_fd_sc_hd__and2_1
XFILLER_0_189_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold30 message_reg.msg\[1\] vssd1 vssd1 vccd1 vccd1 net294 sky130_fd_sc_hd__dlygate4sd3_1
Xhold41 buffer.Rx_byte\[6\] vssd1 vssd1 vccd1 vccd1 net305 sky130_fd_sc_hd__dlygate4sd3_1
Xhold52 _0242_ vssd1 vssd1 vccd1 vccd1 net316 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold74 uart_receiver.clk_count\[4\] vssd1 vssd1 vccd1 vccd1 net338 sky130_fd_sc_hd__dlygate4sd3_1
Xhold63 _0068_ vssd1 vssd1 vccd1 vccd1 net327 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold96 keypadFSMHost.prev_key\[1\] vssd1 vssd1 vccd1 vccd1 net360 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2267__A1 dispFSM.msg\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold85 hostdisp.top\[63\] vssd1 vssd1 vccd1 vccd1 net349 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1570_ _0466_ _0517_ _0450_ vssd1 vssd1 vccd1 vccd1 _0518_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_158_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3240_ clknet_leaf_9_clk keypadFSMHost.next_state\[1\] net215 vssd1 vssd1 vccd1 vccd1
+ _1397_ sky130_fd_sc_hd__dfrtp_1
X_3171_ clknet_leaf_30_clk net348 net185 vssd1 vssd1 vccd1 vccd1 hostdisp.top\[55\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_177_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2122_ hostdisp.curr_guesses\[3\] net119 _0863_ net132 vssd1 vssd1 vccd1 vccd1 hostdisp.nextBottom\[43\]
+ sky130_fd_sc_hd__o211a_1
X_2053_ hostdisp.curr_word\[1\] net98 _0835_ net144 vssd1 vssd1 vccd1 vccd1 hostdisp.next_curr_word\[1\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_76_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_193_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2955_ host_message_reg.setLetter\[2\] net52 net48 gamelogic.setWord\[2\] vssd1 vssd1
+ vccd1 vccd1 _0318_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_20_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1906_ _0752_ _0758_ vssd1 vssd1 vccd1 vccd1 _0759_ sky130_fd_sc_hd__nor2_1
X_2886_ dispFSM.guesses\[26\] net84 net58 net486 vssd1 vssd1 vccd1 vccd1 _0253_ sky130_fd_sc_hd__o22a_1
XFILLER_0_154_291 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1837_ _0716_ _0717_ vssd1 vssd1 vccd1 vccd1 clock_div.next_count\[17\] sky130_fd_sc_hd__nor2_1
XFILLER_0_114_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2981__A2 net52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1768_ _0399_ _0661_ _0667_ _0668_ net328 vssd1 vssd1 vccd1 vccd1 uart_transmitter.next_state\[0\]
+ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout205_A net206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2194__A0 gamelogic.setWord\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3345__Q gamelogic.letter\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3507_ clknet_leaf_29_clk hostdisp.next_curr_word\[29\] net181 vssd1 vssd1 vccd1
+ vccd1 hostdisp.curr_word\[29\] sky130_fd_sc_hd__dfrtp_1
X_1699_ keypadFSMPlayer.state\[4\] keypadFSMPlayer.state\[0\] _0443_ _0449_ _0615_
+ vssd1 vssd1 vccd1 vccd1 _0616_ sky130_fd_sc_hd__o32a_1
XFILLER_0_12_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3438_ clknet_leaf_13_clk _0316_ net199 vssd1 vssd1 vccd1 vccd1 gamelogic.setWord\[0\]
+ sky130_fd_sc_hd__dfstp_1
X_3369_ clknet_leaf_21_clk net407 net202 vssd1 vssd1 vccd1 vccd1 dispFSM.guesses\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_110_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2421__B2 hostdisp.top\[47\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2709__C1 gamelogic.indexCorrect\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_259 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput42 net42 vssd1 vssd1 vccd1 vccd1 gpio_out[32] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_130_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput31 net31 vssd1 vssd1 vccd1 vccd1 gpio_out[12] sky130_fd_sc_hd__buf_2
Xoutput20 net20 vssd1 vssd1 vccd1 vccd1 gpio_oeb[28] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_91_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_187_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1999__B1 net80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3404__CLK clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2740_ keypadFSMHost.state\[1\] keypadFSMHost.state\[4\] vssd1 vssd1 vccd1 vccd1
+ _1294_ sky130_fd_sc_hd__nor2_1
XFILLER_0_26_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2671_ gamelogic.setWord\[33\] net144 vssd1 vssd1 vccd1 vccd1 _1237_ sky130_fd_sc_hd__or2_1
XFILLER_0_26_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1622_ _0542_ _0545_ _0552_ _0540_ vssd1 vssd1 vccd1 vccd1 _0557_ sky130_fd_sc_hd__o211a_2
XFILLER_0_41_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1553_ _0414_ _0416_ vssd1 vssd1 vccd1 vccd1 _0501_ sky130_fd_sc_hd__or2_1
XFILLER_0_111_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1484_ _0417_ _0418_ _0419_ net128 vssd1 vssd1 vccd1 vccd1 _0436_ sky130_fd_sc_hd__or4bb_1
X_3223_ clknet_leaf_16_clk _0197_ net223 vssd1 vssd1 vccd1 vccd1 keypadFSMHost.prev_key\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_185_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3154_ clknet_leaf_16_clk _0130_ net222 vssd1 vssd1 vccd1 vccd1 keypadplayer.scan_col\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_118_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_19_Left_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3085_ clknet_leaf_19_clk _0075_ net211 vssd1 vssd1 vccd1 vccd1 message_reg.msg\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_2105_ hostdisp.curr_word\[33\] net99 _0855_ net144 vssd1 vssd1 vccd1 vccd1 hostdisp.next_curr_word\[33\]
+ sky130_fd_sc_hd__o22a_1
X_2036_ gamelogic.letter\[2\] net91 net76 net527 vssd1 vssd1 vccd1 vccd1 hostdisp.next_curr_guesses\[42\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_166_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3084__CLK clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2938_ dispFSM.guesses\[78\] net87 net60 net543 vssd1 vssd1 vccd1 vccd1 _0305_ sky130_fd_sc_hd__o22a_1
XFILLER_0_17_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_28_Left_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_150_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2954__A2 net53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_157_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2869_ dispFSM.guesses\[9\] net86 net62 net423 vssd1 vssd1 vccd1 vccd1 _0236_ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout110_X net110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3587__259 vssd1 vssd1 vccd1 vccd1 net259 _3587__259/LO sky130_fd_sc_hd__conb_1
XFILLER_0_7_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_168_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_37_Left_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout68_A net69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3427__CLK clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_127_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_184_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_46_Left_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_180_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_180_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_5_clk_A clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_171_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_190_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_30_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_340 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2723_ _1282_ _1283_ _1285_ vssd1 vssd1 vccd1 vccd1 _1286_ sky130_fd_sc_hd__and3b_1
X_2654_ dispFSM.guesses\[15\] _1078_ _1086_ dispFSM.guesses\[79\] _0360_ vssd1 vssd1
+ vccd1 vccd1 _1225_ sky130_fd_sc_hd__a221o_1
X_1605_ net229 net232 vssd1 vssd1 vccd1 vccd1 _0540_ sky130_fd_sc_hd__and2b_1
XANTENNA__1906__Y _0759_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2585_ net139 _1123_ _1154_ net108 _1159_ vssd1 vssd1 vccd1 vccd1 _1160_ sky130_fd_sc_hd__a221o_1
X_1536_ keypadFSMPlayer.prev_key\[5\] _0419_ net128 vssd1 vssd1 vccd1 vccd1 _0484_
+ sky130_fd_sc_hd__and3_1
Xfanout128 _0424_ vssd1 vssd1 vccd1 vccd1 net128 sky130_fd_sc_hd__buf_2
Xfanout106 _0759_ vssd1 vssd1 vccd1 vccd1 net106 sky130_fd_sc_hd__clkbuf_4
Xfanout117 net118 vssd1 vssd1 vccd1 vccd1 net117 sky130_fd_sc_hd__buf_4
X_1467_ net4 net231 vssd1 vssd1 vccd1 vccd1 _0419_ sky130_fd_sc_hd__and2_1
XFILLER_0_38_71 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout139 lcdPlayer.nextState\[0\] vssd1 vssd1 vccd1 vccd1 net139 sky130_fd_sc_hd__buf_2
X_3206_ clknet_leaf_27_clk _0182_ vssd1 vssd1 vccd1 vccd1 lcdPlayer.currentState\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_3137_ clknet_leaf_26_clk _0113_ vssd1 vssd1 vccd1 vccd1 lcdPlayer.cnt_20ms\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_3068_ clknet_leaf_17_clk _0061_ _0030_ vssd1 vssd1 vccd1 vccd1 dispFSM.msg\[3\]
+ sky130_fd_sc_hd__dfstp_2
XPHY_EDGE_ROW_118_Right_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_107_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2019_ hostdisp.curr_guesses\[33\] net93 net78 net463 vssd1 vssd1 vccd1 vccd1 hostdisp.next_curr_guesses\[25\]
+ sky130_fd_sc_hd__o22a_1
XANTENNA__2624__B2 _1078_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_53_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2405__S _0934_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_334 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_162_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold171 _0264_ vssd1 vssd1 vccd1 vccd1 net435 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2140__S net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold160 hostdisp.curr_guesses\[3\] vssd1 vssd1 vccd1 vccd1 net424 sky130_fd_sc_hd__dlygate4sd3_1
Xhold193 hostdisp.curr_guesses\[9\] vssd1 vssd1 vccd1 vccd1 net457 sky130_fd_sc_hd__dlygate4sd3_1
Xhold182 dispFSM.guesses\[13\] vssd1 vssd1 vccd1 vccd1 net446 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2560__B1 net109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2823__B _0827_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_177_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_386 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3000__A net221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_188_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2370_ _1004_ _1005_ vssd1 vssd1 vccd1 vccd1 _0116_ sky130_fd_sc_hd__nor2_1
XANTENNA__2551__B1 _1096_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_147_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2706_ gamelogic.letter\[1\] _0389_ gamelogic.setWord\[18\] _0379_ _1269_ vssd1 vssd1
+ vccd1 vccd1 _1270_ sky130_fd_sc_hd__a221o_1
XFILLER_0_6_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_154_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_12_Right_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2637_ hostdisp.top\[78\] _1095_ _1097_ hostdisp.top\[54\] vssd1 vssd1 vccd1 vccd1
+ _1209_ sky130_fd_sc_hd__a22o_1
XFILLER_0_64_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2542__B1 net108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2568_ hostdisp.top\[67\] _1096_ _1097_ hostdisp.top\[51\] _1141_ vssd1 vssd1 vccd1
+ vccd1 _1143_ sky130_fd_sc_hd__a221o_1
X_1519_ net146 _0462_ vssd1 vssd1 vccd1 vccd1 _0467_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_113_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2499_ dispFSM.guesses\[64\] _1072_ net114 dispFSM.guesses\[24\] vssd1 vssd1 vccd1
+ vccd1 _1077_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_58_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_165_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_21_Right_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_66_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2135__S net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_30_Right_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_231 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2533__B1 _1096_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_185_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_142_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1870_ uart_transmitter.clk_count\[0\] net290 net116 vssd1 vssd1 vccd1 vccd1 _0733_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_126_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3540_ clknet_leaf_6_clk hostdisp.next_curr_guesses\[22\] net191 vssd1 vssd1 vccd1
+ vccd1 hostdisp.curr_guesses\[22\] sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_12_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_66 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3471_ clknet_leaf_7_clk _0349_ net195 vssd1 vssd1 vccd1 vccd1 gamelogic.setWord\[33\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_10_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2422_ net133 _0822_ _0857_ vssd1 vssd1 vccd1 vccd1 _1034_ sky130_fd_sc_hd__and3_4
XANTENNA__2524__B1 net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2353_ lcdPlayer.cnt_20ms\[2\] lcdPlayer.cnt_20ms\[1\] lcdPlayer.cnt_20ms\[0\] net567
+ vssd1 vssd1 vccd1 vccd1 _0995_ sky130_fd_sc_hd__a31o_1
XFILLER_0_19_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2284_ _0949_ _0950_ _0952_ vssd1 vssd1 vccd1 vccd1 _0953_ sky130_fd_sc_hd__or3_1
XFILLER_0_193_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3516__SET_B net165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2463__B _0827_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2460__C1 _1034_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_30_clk_A clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1999_ hostdisp.curr_guesses\[13\] net95 net80 net335 vssd1 vssd1 vccd1 vccd1 hostdisp.next_curr_guesses\[5\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_27_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_115_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_167_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3185__RESET_B net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_170_Right_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3168__CLK clknet_leaf_30_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_324 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_174_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_133_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_163_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2564__A _0764_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_204 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2971_ gamelogic.setWord\[10\] net51 net47 gamelogic.setWord\[18\] vssd1 vssd1 vccd1
+ vccd1 _0334_ sky130_fd_sc_hd__o22a_1
XFILLER_0_8_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1922_ net181 _0772_ vssd1 vssd1 vccd1 vccd1 _0773_ sky130_fd_sc_hd__nand2_1
X_1853_ net503 _0725_ vssd1 vssd1 vccd1 vccd1 _0726_ sky130_fd_sc_hd__nor2_1
XFILLER_0_122_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_276 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1784_ clock_div.count\[27\] clock_div.count\[26\] clock_div.count\[29\] clock_div.count\[28\]
+ vssd1 vssd1 vccd1 vccd1 _0682_ sky130_fd_sc_hd__or4_1
X_3523_ clknet_leaf_15_clk net336 net208 vssd1 vssd1 vccd1 vccd1 hostdisp.curr_guesses\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3454_ clknet_leaf_5_clk _0332_ net196 vssd1 vssd1 vccd1 vccd1 gamelogic.setWord\[16\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_97_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2405_ _0441_ keypadplayer.scan_col\[1\] _0934_ vssd1 vssd1 vccd1 vccd1 _0129_ sky130_fd_sc_hd__mux2_1
X_3385_ clknet_leaf_21_clk net385 net207 vssd1 vssd1 vccd1 vccd1 dispFSM.guesses\[39\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_110_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2336_ net452 _0984_ _0986_ vssd1 vssd1 vccd1 vccd1 _0101_ sky130_fd_sc_hd__o21a_1
XANTENNA__2458__B net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2267_ dispFSM.msg\[1\] _0941_ _0942_ net294 vssd1 vssd1 vccd1 vccd1 _0076_ sky130_fd_sc_hd__a22o_1
XFILLER_0_137_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout185_A net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_162_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2198_ net135 hostdisp.curr_guesses\[41\] net124 _0901_ vssd1 vssd1 vccd1 vccd1 hostdisp.nextBottom\[81\]
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_79_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3460__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout140_X net140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout98_A net100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold20 message_reg.msg\[0\] vssd1 vssd1 vccd1 vccd1 net284 sky130_fd_sc_hd__dlygate4sd3_1
Xhold31 net29 vssd1 vssd1 vccd1 vccd1 net295 sky130_fd_sc_hd__dlygate4sd3_1
Xhold64 uart_transmitter.state\[2\] vssd1 vssd1 vccd1 vccd1 net328 sky130_fd_sc_hd__dlygate4sd3_1
Xhold42 _0073_ vssd1 vssd1 vccd1 vccd1 net306 sky130_fd_sc_hd__dlygate4sd3_1
Xhold53 buffer.Rx_byte\[0\] vssd1 vssd1 vccd1 vccd1 net317 sky130_fd_sc_hd__dlygate4sd3_1
Xhold75 uart_transmitter.bit_index\[2\] vssd1 vssd1 vccd1 vccd1 net339 sky130_fd_sc_hd__dlygate4sd3_1
Xhold97 hostdisp.top\[57\] vssd1 vssd1 vccd1 vccd1 net361 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold86 hostdisp.top\[69\] vssd1 vssd1 vccd1 vccd1 net350 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_187_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_180_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout53_X net53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2975__B1 net49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3170_ clknet_leaf_30_clk _0146_ net174 vssd1 vssd1 vccd1 vccd1 hostdisp.top\[54\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_174_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2121_ gamelogic.setWord\[3\] net121 vssd1 vssd1 vccd1 vccd1 _0863_ sky130_fd_sc_hd__or2_1
X_2052_ _0835_ vssd1 vssd1 vccd1 vccd1 _0836_ sky130_fd_sc_hd__inv_2
XFILLER_0_178_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_190_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2954_ host_message_reg.setLetter\[1\] net53 net49 gamelogic.setWord\[1\] vssd1 vssd1
+ vccd1 vccd1 _0317_ sky130_fd_sc_hd__o22a_1
XFILLER_0_32_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2885_ dispFSM.guesses\[25\] net86 net62 net481 vssd1 vssd1 vccd1 vccd1 _0252_ sky130_fd_sc_hd__o22a_1
XANTENNA__2430__A2 net73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1905_ _0754_ _0755_ _0756_ _0757_ vssd1 vssd1 vccd1 vccd1 _0758_ sky130_fd_sc_hd__or4b_2
X_1836_ clock_div.count\[17\] _0714_ vssd1 vssd1 vccd1 vccd1 _0717_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_6_Right_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1767_ _0398_ _0662_ vssd1 vssd1 vccd1 vccd1 _0669_ sky130_fd_sc_hd__nor2_1
XFILLER_0_12_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout100_A net104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3506_ clknet_leaf_31_clk hostdisp.next_curr_word\[28\] net172 vssd1 vssd1 vccd1
+ vccd1 hostdisp.curr_word\[28\] sky130_fd_sc_hd__dfstp_1
X_1698_ keypadFSMPlayer.state\[4\] keypadFSMPlayer.state\[0\] _0446_ _0442_ vssd1
+ vssd1 vccd1 vccd1 _0615_ sky130_fd_sc_hd__o31a_1
XFILLER_0_12_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3437_ clknet_leaf_17_clk _0016_ _0044_ vssd1 vssd1 vccd1 vccd1 keypadFSMPlayer.state\[5\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_148_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3368_ clknet_leaf_20_clk _0257_ net204 vssd1 vssd1 vccd1 vccd1 dispFSM.guesses\[22\]
+ sky130_fd_sc_hd__dfstp_1
X_2319_ lcdPlayer.cnt_500hz\[12\] _0973_ _0975_ vssd1 vssd1 vccd1 vccd1 _0095_ sky130_fd_sc_hd__o21a_1
XANTENNA__2288__A_N net106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3299_ clknet_leaf_20_clk _0217_ net210 vssd1 vssd1 vccd1 vccd1 message_reg.state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__2408__S _0934_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2654__C1 _0360_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2957__B1 net48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3356__CLK clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput10 net10 vssd1 vssd1 vccd1 vccd1 gpio_oeb[11] sky130_fd_sc_hd__buf_2
Xoutput21 net21 vssd1 vssd1 vccd1 vccd1 gpio_oeb[29] sky130_fd_sc_hd__buf_2
Xoutput43 net43 vssd1 vssd1 vccd1 vccd1 gpio_out[6] sky130_fd_sc_hd__buf_2
Xoutput32 net32 vssd1 vssd1 vccd1 vccd1 gpio_out[13] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_91_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_28 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_168_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_59_Right_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2670_ _0929_ net66 vssd1 vssd1 vccd1 vccd1 _1236_ sky130_fd_sc_hd__and2_1
XFILLER_0_169_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1621_ _0542_ _0553_ _0555_ vssd1 vssd1 vccd1 vccd1 _0556_ sky130_fd_sc_hd__or3_2
XANTENNA__3217__RESET_B net164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1552_ net232 _0415_ _0435_ _0461_ vssd1 vssd1 vccd1 vccd1 _0500_ sky130_fd_sc_hd__or4_1
XFILLER_0_1_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1483_ _0419_ net128 vssd1 vssd1 vccd1 vccd1 _0435_ sky130_fd_sc_hd__nand2_1
X_3222_ clknet_leaf_10_clk net266 net216 vssd1 vssd1 vccd1 vccd1 keypadFSMHost.strobe_edge
+ sky130_fd_sc_hd__dfrtp_1
X_3153_ clknet_leaf_16_clk _0129_ net222 vssd1 vssd1 vccd1 vccd1 keypadplayer.scan_col\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_68_Right_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2104_ hostdisp.curr_word\[32\] net99 _0855_ net145 vssd1 vssd1 vccd1 vccd1 hostdisp.next_curr_word\[32\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_118_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3084_ clknet_leaf_33_clk net308 net160 vssd1 vssd1 vccd1 vccd1 buffer.temp_guess\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_2035_ net144 net93 net78 net475 vssd1 vssd1 vccd1 vccd1 hostdisp.next_curr_guesses\[41\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_134_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_174_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2651__A2 _1097_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3379__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_77_Right_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_174_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2937_ net426 net90 net64 net430 vssd1 vssd1 vccd1 vccd1 _0304_ sky130_fd_sc_hd__a22o_1
XFILLER_0_57_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_157_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2868_ dispFSM.guesses\[8\] net81 net56 net464 vssd1 vssd1 vccd1 vccd1 _0235_ sky130_fd_sc_hd__o22a_1
X_1819_ clock_div.count\[10\] _0703_ net531 vssd1 vssd1 vccd1 vccd1 _0706_ sky130_fd_sc_hd__a21oi_1
X_2799_ _0385_ gamelogic.setWord\[14\] gamelogic.setWord\[8\] _0377_ vssd1 vssd1 vccd1
+ vccd1 _1345_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_4_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2199__A net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_86_Right_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_175_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_168_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2138__S net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_95_Right_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_192_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_2_Left_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2633__A2 net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3521__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_156_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_156_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_171_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2722_ net145 _0390_ gamelogic.setWord\[4\] _0382_ _1284_ vssd1 vssd1 vccd1 vccd1
+ _1285_ sky130_fd_sc_hd__o221a_1
XFILLER_0_54_352 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2653_ dispFSM.guesses\[31\] net115 net110 dispFSM.guesses\[39\] _1223_ vssd1 vssd1
+ vccd1 vccd1 _1224_ sky130_fd_sc_hd__a221o_1
X_1604_ net229 net6 vssd1 vssd1 vccd1 vccd1 _0539_ sky130_fd_sc_hd__and2b_1
X_2584_ _1156_ _1158_ net106 vssd1 vssd1 vccd1 vccd1 _1159_ sky130_fd_sc_hd__o21ai_1
X_1535_ _0481_ _0482_ _0479_ vssd1 vssd1 vccd1 vccd1 _0483_ sky130_fd_sc_hd__o21a_1
Xfanout129 _0375_ vssd1 vssd1 vccd1 vccd1 net129 sky130_fd_sc_hd__buf_4
Xfanout107 _0759_ vssd1 vssd1 vccd1 vccd1 net107 sky130_fd_sc_hd__clkbuf_2
Xfanout118 _1079_ vssd1 vssd1 vccd1 vccd1 net118 sky130_fd_sc_hd__clkbuf_4
X_1466_ net231 net3 vssd1 vssd1 vccd1 vccd1 _0418_ sky130_fd_sc_hd__and2_1
XFILLER_0_38_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3205_ clknet_leaf_24_clk _0181_ vssd1 vssd1 vccd1 vccd1 net32 sky130_fd_sc_hd__dfxtp_1
X_3136_ clknet_leaf_26_clk net270 vssd1 vssd1 vccd1 vccd1 lcdPlayer.cnt_20ms\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_3067_ clknet_leaf_21_clk _0060_ _0029_ vssd1 vssd1 vccd1 vccd1 dispFSM.msg\[2\]
+ sky130_fd_sc_hd__dfstp_2
X_2018_ hostdisp.curr_guesses\[32\] net93 net78 net484 vssd1 vssd1 vccd1 vccd1 hostdisp.next_curr_guesses\[24\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_49_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_346 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_240 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold161 dispFSM.guesses\[55\] vssd1 vssd1 vccd1 vccd1 net425 sky130_fd_sc_hd__dlygate4sd3_1
Xhold150 hostdisp.curr_guesses\[4\] vssd1 vssd1 vccd1 vccd1 net414 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold172 hostdisp.curr_guesses\[1\] vssd1 vssd1 vccd1 vccd1 net436 sky130_fd_sc_hd__dlygate4sd3_1
Xhold183 hostdisp.top\[43\] vssd1 vssd1 vccd1 vccd1 net447 sky130_fd_sc_hd__dlygate4sd3_1
Xhold194 hostdisp.curr_guesses\[43\] vssd1 vssd1 vccd1 vccd1 net458 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_69_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_44_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_177_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2823__C net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_180_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_188_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_184_Right_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_298 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2606__A2 net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_173 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2705_ net145 gamelogic.setWord\[16\] vssd1 vssd1 vccd1 vccd1 _1269_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_154_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2790__B2 host_message_reg.setLetter\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3417__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2636_ _1204_ _1206_ _1207_ net227 vssd1 vssd1 vccd1 vccd1 _1208_ sky130_fd_sc_hd__o31a_1
XFILLER_0_42_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_65_Left_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_151_Right_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2567_ _0356_ _1064_ vssd1 vssd1 vccd1 vccd1 _1142_ sky130_fd_sc_hd__nor2_1
X_1518_ net232 _0435_ _0458_ vssd1 vssd1 vccd1 vccd1 _0466_ sky130_fd_sc_hd__or3_1
XANTENNA__2542__B2 dispFSM.msg\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2498_ _1073_ _1074_ vssd1 vssd1 vccd1 vccd1 _1076_ sky130_fd_sc_hd__nor2_1
X_1449_ uart_transmitter.bit_index\[0\] vssd1 vssd1 vccd1 vccd1 _0402_ sky130_fd_sc_hd__inv_2
XANTENNA__2477__A net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_165_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_4_clk_A clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_74_Left_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_167_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3119_ clknet_leaf_34_clk _0106_ net158 vssd1 vssd1 vccd1 vccd1 uart_receiver.bit_index\[2\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_66_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_147_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_316 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_83_Left_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2151__S net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_243 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_92_Left_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_158_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3011__A net223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_142_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1466__A net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3470_ clknet_leaf_5_clk _0348_ net192 vssd1 vssd1 vccd1 vccd1 gamelogic.setWord\[32\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_101_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2421_ net514 net72 net69 hostdisp.top\[47\] vssd1 vssd1 vccd1 vccd1 _0139_ sky130_fd_sc_hd__a22o_1
X_2352_ net167 _0944_ _0994_ _0955_ vssd1 vssd1 vccd1 vccd1 _0109_ sky130_fd_sc_hd__a31o_1
XANTENNA__2297__A _0752_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2283_ lcdPlayer.cnt_20ms\[12\] lcdPlayer.cnt_20ms\[9\] lcdPlayer.cnt_20ms\[7\] _0951_
+ vssd1 vssd1 vccd1 vccd1 _0952_ sky130_fd_sc_hd__or4b_1
XFILLER_0_193_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_191_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_191_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_142_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2460__B1 net71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout228_A net7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_379 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1998_ hostdisp.curr_guesses\[12\] net92 net77 net414 vssd1 vssd1 vccd1 vccd1 hostdisp.next_curr_guesses\[4\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_27_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2619_ hostdisp.bottom\[101\] dispFSM.guesses\[13\] net228 vssd1 vssd1 vccd1 vccd1
+ _1192_ sky130_fd_sc_hd__mux2_1
X_3599_ net264 vssd1 vssd1 vccd1 vccd1 gpio_oeb[33] sky130_fd_sc_hd__buf_2
XANTENNA__3234__SET_B net221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_3_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_183_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2146__S net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_174_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_346 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_133_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_94_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_85_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkload6_A clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3262__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2970_ gamelogic.setWord\[9\] net54 net50 gamelogic.setWord\[17\] vssd1 vssd1 vccd1
+ vccd1 _0333_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_103_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1921_ lcdPlayer.nextState\[5\] lcdPlayer.currentState\[5\] _0764_ vssd1 vssd1 vccd1
+ vccd1 _0772_ sky130_fd_sc_hd__mux2_1
X_1852_ _0724_ _0725_ vssd1 vssd1 vccd1 vccd1 clock_div.next_count\[24\] sky130_fd_sc_hd__nor2_1
XFILLER_0_56_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_188_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1783_ _0676_ _0680_ _0681_ _0662_ vssd1 vssd1 vccd1 vccd1 uart_transmitter.tx_serial
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_114_327 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3522_ clknet_leaf_4_clk hostdisp.next_curr_guesses\[4\] net177 vssd1 vssd1 vccd1
+ vccd1 hostdisp.curr_guesses\[4\] sky130_fd_sc_hd__dfstp_1
XPHY_EDGE_ROW_139_Left_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3453_ clknet_leaf_14_clk _0331_ net193 vssd1 vssd1 vccd1 vccd1 gamelogic.setWord\[15\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_122_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2404_ _1027_ keypadplayer.scan_col\[0\] _0934_ vssd1 vssd1 vccd1 vccd1 _0128_ sky130_fd_sc_hd__mux2_1
X_3384_ clknet_leaf_20_clk _0273_ net204 vssd1 vssd1 vccd1 vccd1 dispFSM.guesses\[38\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_110_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2335_ lcdPlayer.cnt_500hz\[18\] _0984_ _0957_ vssd1 vssd1 vccd1 vccd1 _0986_ sky130_fd_sc_hd__a21oi_1
X_2266_ dispFSM.msg\[0\] _0941_ _0942_ net284 vssd1 vssd1 vccd1 vccd1 _0075_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_162_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2197_ net130 gamelogic.setWord\[33\] vssd1 vssd1 vccd1 vccd1 _0901_ sky130_fd_sc_hd__and2_1
XFILLER_0_79_303 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2130__C1 net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout178_A net179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_148_Left_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_121_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_238 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2984__B2 gamelogic.setWord\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout133_X net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_157_Left_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_319 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2200__A3 net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold21 keypadFSMHost.unlocked vssd1 vssd1 vccd1 vccd1 net285 sky130_fd_sc_hd__dlygate4sd3_1
Xhold32 net31 vssd1 vssd1 vccd1 vccd1 net296 sky130_fd_sc_hd__dlygate4sd3_1
Xhold10 _0127_ vssd1 vssd1 vccd1 vccd1 net274 sky130_fd_sc_hd__dlygate4sd3_1
Xhold43 buffer.Rx_byte\[7\] vssd1 vssd1 vccd1 vccd1 net307 sky130_fd_sc_hd__dlygate4sd3_1
Xhold54 _0067_ vssd1 vssd1 vccd1 vccd1 net318 sky130_fd_sc_hd__dlygate4sd3_1
Xhold65 hostdisp.top\[54\] vssd1 vssd1 vccd1 vccd1 net329 sky130_fd_sc_hd__dlygate4sd3_1
Xhold87 message_reg.msg\[3\] vssd1 vssd1 vccd1 vccd1 net351 sky130_fd_sc_hd__dlygate4sd3_1
Xhold76 hostdisp.top\[58\] vssd1 vssd1 vccd1 vccd1 net340 sky130_fd_sc_hd__dlygate4sd3_1
Xhold98 hostdisp.top\[59\] vssd1 vssd1 vccd1 vccd1 net362 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3285__CLK clknet_leaf_30_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_180_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_166_Left_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_39_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2120_ hostdisp.curr_guesses\[2\] net119 _0862_ net131 vssd1 vssd1 vccd1 vccd1 hostdisp.nextBottom\[42\]
+ sky130_fd_sc_hd__o211a_1
X_2051_ _0403_ net96 _0831_ _0834_ vssd1 vssd1 vccd1 vccd1 _0835_ sky130_fd_sc_hd__a211o_2
XFILLER_0_16_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_99 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2953_ host_message_reg.setLetter\[0\] net53 net50 gamelogic.setWord\[0\] vssd1 vssd1
+ vccd1 vccd1 _0316_ sky130_fd_sc_hd__o22a_1
XANTENNA__2415__B1 net69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_290 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1904_ lcdPlayer.cnt_500hz\[8\] lcdPlayer.cnt_500hz\[9\] lcdPlayer.cnt_500hz\[11\]
+ lcdPlayer.cnt_500hz\[10\] vssd1 vssd1 vccd1 vccd1 _0757_ sky130_fd_sc_hd__and4b_1
XFILLER_0_84_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2884_ dispFSM.guesses\[24\] net81 net56 net547 vssd1 vssd1 vccd1 vccd1 _0251_ sky130_fd_sc_hd__o22a_1
X_1835_ clock_div.count\[17\] _0714_ vssd1 vssd1 vccd1 vccd1 _0716_ sky130_fd_sc_hd__nor2_1
XFILLER_0_4_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1766_ uart_transmitter.state\[0\] _0664_ vssd1 vssd1 vccd1 vccd1 _0668_ sky130_fd_sc_hd__or2_1
XANTENNA__3158__CLK clknet_leaf_31_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3505_ clknet_leaf_31_clk hostdisp.next_curr_word\[27\] net173 vssd1 vssd1 vccd1
+ vccd1 hostdisp.curr_word\[27\] sky130_fd_sc_hd__dfstp_1
X_1697_ _0009_ _0010_ _0008_ vssd1 vssd1 vccd1 vccd1 keypadFSMHost.next_state\[0\]
+ sky130_fd_sc_hd__or3_1
XFILLER_0_12_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3436_ clknet_leaf_18_clk _0015_ _0043_ vssd1 vssd1 vccd1 vccd1 keypadFSMPlayer.state\[4\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_110_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3367_ clknet_leaf_20_clk net396 net203 vssd1 vssd1 vccd1 vccd1 dispFSM.guesses\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_2318_ lcdPlayer.cnt_500hz\[12\] _0973_ net74 vssd1 vssd1 vccd1 vccd1 _0975_ sky130_fd_sc_hd__a21oi_1
X_3298_ clknet_leaf_19_clk _0216_ net210 vssd1 vssd1 vccd1 vccd1 message_reg.state\[0\]
+ sky130_fd_sc_hd__dfrtp_2
X_2249_ _0600_ net152 _0937_ vssd1 vssd1 vccd1 vccd1 _0047_ sky130_fd_sc_hd__mux2_1
XFILLER_0_164_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2654__B1 _1086_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_36_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_192_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2957__A1 host_message_reg.setLetter\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput33 net33 vssd1 vssd1 vccd1 vccd1 gpio_out[16] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_130_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput22 net22 vssd1 vssd1 vccd1 vccd1 gpio_oeb[30] sky130_fd_sc_hd__buf_2
Xoutput11 net11 vssd1 vssd1 vccd1 vccd1 gpio_oeb[12] sky130_fd_sc_hd__buf_2
Xoutput9 net9 vssd1 vssd1 vccd1 vccd1 gpio_oeb[10] sky130_fd_sc_hd__buf_2
Xoutput44 net44 vssd1 vssd1 vccd1 vccd1 gpio_out[7] sky130_fd_sc_hd__buf_2
XFILLER_0_9_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_187_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1999__A2 net95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_100_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3300__CLK clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1620_ _0544_ _0552_ vssd1 vssd1 vccd1 vccd1 _0555_ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1551_ _0496_ _0498_ vssd1 vssd1 vccd1 vccd1 _0499_ sky130_fd_sc_hd__xor2_2
XANTENNA__1474__A net4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3450__CLK clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1482_ _0422_ _0426_ _0432_ _0433_ vssd1 vssd1 vccd1 vccd1 _0434_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_185_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3221_ clknet_leaf_10_clk net268 net216 vssd1 vssd1 vccd1 vccd1 keypadFSMHost.strobe_edge1
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_182_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3152_ clknet_leaf_16_clk _0128_ net222 vssd1 vssd1 vccd1 vccd1 keypadplayer.scan_col\[0\]
+ sky130_fd_sc_hd__dfrtp_4
X_2103_ _0855_ vssd1 vssd1 vccd1 vccd1 _0856_ sky130_fd_sc_hd__inv_2
X_3083_ clknet_leaf_33_clk net306 net160 vssd1 vssd1 vccd1 vccd1 buffer.temp_guess\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_2034_ net145 net94 net79 net492 vssd1 vssd1 vccd1 vccd1 hostdisp.next_curr_guesses\[40\]
+ sky130_fd_sc_hd__o22a_1
XANTENNA__2636__B1 net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_174_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2936_ dispFSM.guesses\[76\] net84 net58 net524 vssd1 vssd1 vccd1 vccd1 _0303_ sky130_fd_sc_hd__o22a_1
XFILLER_0_17_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2867_ _0465_ net88 vssd1 vssd1 vccd1 vccd1 _1391_ sky130_fd_sc_hd__or2_1
X_1818_ clock_div.count\[10\] _0703_ _0705_ _0693_ vssd1 vssd1 vccd1 vccd1 clock_div.next_count\[10\]
+ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_157_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2798_ _0377_ gamelogic.setWord\[8\] gamelogic.setWord\[15\] _0386_ vssd1 vssd1 vccd1
+ vccd1 _1344_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_7_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1749_ _0654_ vssd1 vssd1 vccd1 vccd1 _0655_ sky130_fd_sc_hd__inv_2
X_3419_ clknet_leaf_20_clk _0308_ net205 vssd1 vssd1 vccd1 vccd1 dispFSM.guesses\[73\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_168_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_191_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_165_Right_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3570__254 vssd1 vssd1 vccd1 vccd1 net254 _3570__254/LO sky130_fd_sc_hd__conb_1
XFILLER_0_31_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2094__B2 net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_103_Left_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2721_ _0378_ gamelogic.setWord\[1\] gamelogic.setWord\[2\] _0379_ vssd1 vssd1 vccd1
+ vccd1 _1284_ sky130_fd_sc_hd__o22a_1
XPHY_EDGE_ROW_132_Right_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2652_ dispFSM.guesses\[55\] net113 _1085_ dispFSM.guesses\[47\] vssd1 vssd1 vccd1
+ vccd1 _1223_ sky130_fd_sc_hd__a22o_1
XFILLER_0_89_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1603_ keypadFSMHost.strobe_edge1 keypadFSMHost.strobe_edge vssd1 vssd1 vccd1 vccd1
+ _0538_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_10_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2583_ _1083_ _1123_ _1155_ _1157_ vssd1 vssd1 vccd1 vccd1 _1158_ sky130_fd_sc_hd__or4_1
X_1534_ keypadplayer.scan_col\[0\] net154 keypadFSMPlayer.prev_key\[0\] vssd1 vssd1
+ vccd1 vccd1 _0482_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_129_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout119 _0859_ vssd1 vssd1 vccd1 vccd1 net119 sky130_fd_sc_hd__buf_2
Xfanout108 _1106_ vssd1 vssd1 vccd1 vccd1 net108 sky130_fd_sc_hd__clkbuf_4
XANTENNA__3020__RESET_B net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1465_ net232 net6 net231 vssd1 vssd1 vccd1 vccd1 _0417_ sky130_fd_sc_hd__o21a_1
X_3204_ clknet_leaf_20_clk _0180_ vssd1 vssd1 vccd1 vccd1 net31 sky130_fd_sc_hd__dfxtp_1
X_3135_ clknet_leaf_27_clk _0111_ vssd1 vssd1 vccd1 vccd1 lcdPlayer.cnt_20ms\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_3066_ clknet_leaf_19_clk _0059_ _0028_ vssd1 vssd1 vccd1 vccd1 dispFSM.msg\[1\]
+ sky130_fd_sc_hd__dfstp_1
X_2017_ net433 net95 net80 net439 vssd1 vssd1 vccd1 vccd1 hostdisp.next_curr_guesses\[23\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__2085__B2 net140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout160_A net225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_136 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_147_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3496__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_314 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2919_ dispFSM.guesses\[59\] net81 net57 net506 vssd1 vssd1 vccd1 vccd1 _0286_ sky130_fd_sc_hd__o22a_1
XFILLER_0_162_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_118_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_252 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold140 keypadFSMHost.prev_key\[6\] vssd1 vssd1 vccd1 vccd1 net404 sky130_fd_sc_hd__dlygate4sd3_1
Xhold162 dispFSM.guesses\[77\] vssd1 vssd1 vccd1 vccd1 net426 sky130_fd_sc_hd__dlygate4sd3_1
Xhold151 hostdisp.top\[71\] vssd1 vssd1 vccd1 vccd1 net415 sky130_fd_sc_hd__dlygate4sd3_1
Xhold173 clock_div.count\[1\] vssd1 vssd1 vccd1 vccd1 net437 sky130_fd_sc_hd__dlygate4sd3_1
Xhold184 clock_div.count\[2\] vssd1 vssd1 vccd1 vccd1 net448 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2560__A2 net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold195 dispFSM.guesses\[48\] vssd1 vssd1 vccd1 vccd1 net459 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2149__S net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_177_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_180_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_312 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3219__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_188_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2551__A2 _1095_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3369__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_188_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_111_Left_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_106_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2067__B2 gamelogic.letter\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2704_ _0384_ gamelogic.setWord\[21\] gamelogic.setWord\[22\] _0385_ _1267_ vssd1
+ vssd1 vccd1 vccd1 _1268_ sky130_fd_sc_hd__o221a_1
XANTENNA__3272__RESET_B net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_120_Left_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2635_ dispFSM.guesses\[54\] net113 net111 dispFSM.guesses\[46\] _1203_ vssd1 vssd1
+ vccd1 vccd1 _1207_ sky130_fd_sc_hd__a221o_1
XFILLER_0_42_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2542__A2 _1081_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2566_ hostdisp.bottom\[75\] net112 _1098_ hostdisp.top\[43\] vssd1 vssd1 vccd1 vccd1
+ _1141_ sky130_fd_sc_hd__a22o_1
X_1517_ dispFSM.msg\[5\] _0455_ _0456_ _0465_ vssd1 vssd1 vccd1 vccd1 _0063_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_113_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2497_ _1074_ vssd1 vssd1 vccd1 vccd1 _1075_ sky130_fd_sc_hd__inv_2
X_1448_ uart_transmitter.bit_index\[1\] vssd1 vssd1 vccd1 vccd1 _0401_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_165_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3118_ clknet_leaf_33_clk _0105_ net158 vssd1 vssd1 vccd1 vccd1 uart_receiver.bit_index\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_66_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3049_ clknet_leaf_7_clk clock_div.next_count\[29\] net195 vssd1 vssd1 vccd1 vccd1
+ clock_div.count\[29\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__2058__B2 gamelogic.letter\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_150_328 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_255 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2533__A2 net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_183_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_142_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_72_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_336 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout90 _0939_ vssd1 vssd1 vccd1 vccd1 net90 sky130_fd_sc_hd__buf_2
XFILLER_0_24_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1466__B net3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2420_ hostdisp.curr_word\[6\] net72 net69 hostdisp.top\[46\] vssd1 vssd1 vccd1 vccd1
+ _0138_ sky130_fd_sc_hd__a22o_1
XFILLER_0_177_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3191__CLK clknet_leaf_31_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2524__A2 net114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2351_ lcdPlayer.cnt_20ms\[1\] lcdPlayer.cnt_20ms\[0\] lcdPlayer.cnt_20ms\[2\] vssd1
+ vssd1 vccd1 vccd1 _0994_ sky130_fd_sc_hd__a21o_1
X_2282_ lcdPlayer.cnt_20ms\[6\] lcdPlayer.cnt_20ms\[8\] lcdPlayer.cnt_20ms\[10\] lcdPlayer.cnt_20ms\[11\]
+ vssd1 vssd1 vccd1 vccd1 _0951_ sky130_fd_sc_hd__and4b_1
XFILLER_0_193_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_31 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1997_ hostdisp.curr_guesses\[11\] net91 net76 net424 vssd1 vssd1 vccd1 vccd1 hostdisp.next_curr_guesses\[3\]
+ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout123_A net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3534__CLK clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3598_ net24 vssd1 vssd1 vccd1 vccd1 net23 sky130_fd_sc_hd__clkbuf_1
X_2618_ net226 hostdisp.top\[53\] vssd1 vssd1 vccd1 vccd1 _1191_ sky130_fd_sc_hd__or2_1
X_2549_ net282 net106 _1125_ net188 vssd1 vssd1 vccd1 vccd1 _0175_ sky130_fd_sc_hd__o211a_1
XFILLER_0_167_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2494__Y _1072_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_183_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_26_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2951__A net104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2162__S net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_133_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3290__Q hostdisp.bottom\[101\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3407__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_85_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1920_ _0768_ _0184_ vssd1 vssd1 vccd1 vccd1 _0771_ sky130_fd_sc_hd__nand2_1
X_1851_ clock_div.count\[23\] clock_div.count\[24\] _0723_ vssd1 vssd1 vccd1 vccd1
+ _0725_ sky130_fd_sc_hd__and3_1
XANTENNA__3557__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1477__A net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1782_ message_reg.state\[0\] _0370_ uart_transmitter.state\[0\] vssd1 vssd1 vccd1
+ vccd1 _0681_ sky130_fd_sc_hd__o21a_1
XFILLER_0_114_339 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3521_ clknet_leaf_2_clk hostdisp.next_curr_guesses\[3\] net180 vssd1 vssd1 vccd1
+ vccd1 hostdisp.curr_guesses\[3\] sky130_fd_sc_hd__dfstp_1
XFILLER_0_141_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_3_clk_A clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3452_ clknet_leaf_5_clk _0330_ net193 vssd1 vssd1 vccd1 vccd1 gamelogic.setWord\[14\]
+ sky130_fd_sc_hd__dfstp_1
X_2403_ keypadplayer.scan_col\[0\] _0414_ net148 vssd1 vssd1 vccd1 vccd1 _1027_ sky130_fd_sc_hd__and3b_1
X_3383_ clknet_leaf_21_clk net374 net202 vssd1 vssd1 vccd1 vccd1 dispFSM.guesses\[37\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__1924__B net106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2334_ net275 _0982_ _0985_ vssd1 vssd1 vccd1 vccd1 _0100_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_110_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2265_ _0370_ net86 message_reg.state\[0\] vssd1 vssd1 vccd1 vccd1 _0942_ sky130_fd_sc_hd__a21o_2
XFILLER_0_137_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2196_ net134 hostdisp.curr_guesses\[40\] net124 _0900_ vssd1 vssd1 vccd1 vccd1 hostdisp.nextBottom\[80\]
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_46_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_315 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_162_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_121_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2433__B2 _0828_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout126_X net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold11 lcdPlayer.cnt_500hz\[17\] vssd1 vssd1 vccd1 vccd1 net275 sky130_fd_sc_hd__dlygate4sd3_1
Xhold22 net45 vssd1 vssd1 vccd1 vccd1 net286 sky130_fd_sc_hd__dlygate4sd3_1
Xhold44 _0074_ vssd1 vssd1 vccd1 vccd1 net308 sky130_fd_sc_hd__dlygate4sd3_1
Xhold33 buffer.Rx_byte\[5\] vssd1 vssd1 vccd1 vccd1 net297 sky130_fd_sc_hd__dlygate4sd3_1
Xhold55 lcdPlayer.cnt_500hz\[7\] vssd1 vssd1 vccd1 vccd1 net319 sky130_fd_sc_hd__dlygate4sd3_1
Xhold99 clock_div.count\[26\] vssd1 vssd1 vccd1 vccd1 net363 sky130_fd_sc_hd__dlygate4sd3_1
Xhold88 message_reg.msg\[5\] vssd1 vssd1 vccd1 vccd1 net352 sky130_fd_sc_hd__dlygate4sd3_1
Xhold77 hostdisp.top\[62\] vssd1 vssd1 vccd1 vccd1 net341 sky130_fd_sc_hd__dlygate4sd3_1
Xhold66 hostdisp.top\[72\] vssd1 vssd1 vccd1 vccd1 net330 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_180_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2157__S net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2975__A2 net53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2620__S net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_150_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3017__A net223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2050_ net145 _0831_ _0834_ hostdisp.curr_word\[0\] net98 vssd1 vssd1 vccd1 vccd1
+ hostdisp.next_curr_word\[0\] sky130_fd_sc_hd__o32a_1
XFILLER_0_178_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_179_Right_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2952_ net97 net54 vssd1 vssd1 vccd1 vccd1 _1395_ sky130_fd_sc_hd__nand2_1
XFILLER_0_29_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1903_ lcdPlayer.cnt_500hz\[13\] lcdPlayer.cnt_500hz\[12\] lcdPlayer.cnt_500hz\[14\]
+ vssd1 vssd1 vccd1 vccd1 _0756_ sky130_fd_sc_hd__or3b_1
X_2883_ net406 net88 net65 net441 vssd1 vssd1 vccd1 vccd1 _0250_ sky130_fd_sc_hd__a22o_1
XFILLER_0_32_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1834_ _0714_ _0715_ vssd1 vssd1 vccd1 vccd1 clock_div.next_count\[16\] sky130_fd_sc_hd__nor2_1
XFILLER_0_4_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1765_ uart_transmitter.state\[0\] uart_transmitter.bit_index\[2\] _0665_ _0662_
+ vssd1 vssd1 vccd1 vccd1 _0667_ sky130_fd_sc_hd__a31oi_1
XANTENNA__2718__A2 gamelogic.setWord\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3195__Q hostdisp.top\[79\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3504_ clknet_leaf_31_clk hostdisp.next_curr_word\[26\] net173 vssd1 vssd1 vccd1
+ vccd1 hostdisp.curr_word\[26\] sky130_fd_sc_hd__dfstp_1
X_3435_ clknet_leaf_17_clk _0014_ _0042_ vssd1 vssd1 vccd1 vccd1 keypadFSMPlayer.state\[3\]
+ sky130_fd_sc_hd__dfrtp_2
X_1696_ keypadFSMHost.state\[3\] _0565_ _0605_ _0614_ vssd1 vssd1 vccd1 vccd1 _0008_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_148_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3366_ clknet_leaf_21_clk _0255_ net203 vssd1 vssd1 vccd1 vccd1 dispFSM.guesses\[20\]
+ sky130_fd_sc_hd__dfstp_1
X_3297_ clknet_leaf_34_clk uart_receiver.next_state\[2\] net158 vssd1 vssd1 vccd1
+ vccd1 uart_receiver.state\[2\] sky130_fd_sc_hd__dfrtp_1
X_2317_ lcdPlayer.cnt_500hz\[11\] _0971_ _0974_ vssd1 vssd1 vccd1 vccd1 _0094_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout190_A net225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2248_ _0935_ keypadHostt.scan_col\[0\] _0937_ vssd1 vssd1 vccd1 vccd1 _0046_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2179_ gamelogic.setWord\[32\] hostdisp.curr_guesses\[32\] net124 vssd1 vssd1 vccd1
+ vccd1 _0892_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_146_Right_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_36_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_192_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_180_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2957__A2 net52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_192_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_189_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2590__B1 _1095_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput12 net12 vssd1 vssd1 vccd1 vccd1 gpio_oeb[13] sky130_fd_sc_hd__buf_2
Xoutput23 net23 vssd1 vssd1 vccd1 vccd1 gpio_oeb[31] sky130_fd_sc_hd__buf_2
Xoutput34 net34 vssd1 vssd1 vccd1 vccd1 gpio_out[17] sky130_fd_sc_hd__buf_2
Xoutput45 net45 vssd1 vssd1 vccd1 vccd1 gpio_out[8] sky130_fd_sc_hd__buf_2
XANTENNA__3252__CLK clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_113_Right_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2615__S net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_2_0__f_clk_X clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1550_ keypadFSMPlayer.state\[5\] _0497_ _0492_ _0490_ _0469_ vssd1 vssd1 vccd1 vccd1
+ _0498_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_151_264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1481_ _0417_ _0420_ net128 _0431_ vssd1 vssd1 vccd1 vccd1 _0433_ sky130_fd_sc_hd__and4_1
XFILLER_0_185_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3220_ clknet_leaf_31_clk _0196_ net172 vssd1 vssd1 vccd1 vccd1 gamelogic.indexCorrect\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_94_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3151_ clknet_leaf_26_clk net274 vssd1 vssd1 vccd1 vccd1 lcdPlayer.cnt_20ms\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_175_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1687__A2 keypadFSMHost.state\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2102_ _0853_ _0854_ vssd1 vssd1 vccd1 vccd1 _0855_ sky130_fd_sc_hd__nand2_2
X_3082_ clknet_leaf_33_clk net298 net160 vssd1 vssd1 vccd1 vccd1 buffer.temp_guess\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_178_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2033_ hostdisp.curr_guesses\[47\] net95 net80 net393 vssd1 vssd1 vccd1 vccd1 hostdisp.next_curr_guesses\[39\]
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_109_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_185_Left_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_174_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2935_ dispFSM.guesses\[75\] net82 net57 net474 vssd1 vssd1 vccd1 vccd1 _0302_ sky130_fd_sc_hd__o22a_1
XFILLER_0_174_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2866_ _0465_ net88 vssd1 vssd1 vccd1 vccd1 _1390_ sky130_fd_sc_hd__nor2_1
X_1817_ clock_div.count\[10\] _0703_ vssd1 vssd1 vccd1 vccd1 _0705_ sky130_fd_sc_hd__nand2_1
Xhold300 clock_div.count\[14\] vssd1 vssd1 vccd1 vccd1 net564 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3275__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2797_ gamelogic.letter\[2\] gamelogic.setWord\[10\] vssd1 vssd1 vccd1 vccd1 _1343_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_25_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_142_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1748_ uart_receiver.clk_count\[6\] uart_receiver.clk_count\[7\] _0649_ vssd1 vssd1
+ vccd1 vccd1 _0654_ sky130_fd_sc_hd__and3_1
X_1679_ _0601_ vssd1 vssd1 vccd1 vccd1 _0602_ sky130_fd_sc_hd__inv_2
XFILLER_0_110_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3418_ clknet_leaf_23_clk _0307_ net187 vssd1 vssd1 vccd1 vccd1 dispFSM.guesses\[72\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA_input8_A nrst vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3349_ clknet_leaf_24_clk _0238_ net187 vssd1 vssd1 vccd1 vccd1 dispFSM.guesses\[3\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_168_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2627__B2 _1097_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2627__A1 _1096_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_184_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_192_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_47_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2720_ _0385_ gamelogic.setWord\[6\] _0392_ _1277_ _1278_ vssd1 vssd1 vccd1 vccd1
+ _1283_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_66_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2651_ hostdisp.top\[55\] _1097_ _1219_ _1221_ vssd1 vssd1 vccd1 vccd1 _1222_ sky130_fd_sc_hd__a211o_1
XFILLER_0_54_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1602_ keypadFSMHost.strobe_edge1 keypadFSMHost.strobe_edge vssd1 vssd1 vccd1 vccd1
+ _0537_ sky130_fd_sc_hd__and2b_2
XFILLER_0_22_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2554__B1 net109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2582_ net138 net139 _1057_ _1082_ vssd1 vssd1 vccd1 vccd1 _1157_ sky130_fd_sc_hd__and4b_1
X_1533_ keypadFSMPlayer.prev_key\[0\] keypadplayer.scan_col\[0\] net154 vssd1 vssd1
+ vccd1 vccd1 _0481_ sky130_fd_sc_hd__and3_1
XFILLER_0_1_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1464_ net229 net232 vssd1 vssd1 vccd1 vccd1 _0416_ sky130_fd_sc_hd__nand2_1
Xfanout109 _1087_ vssd1 vssd1 vccd1 vccd1 net109 sky130_fd_sc_hd__buf_4
X_3203_ clknet_leaf_24_clk _0179_ vssd1 vssd1 vccd1 vccd1 net30 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3134_ clknet_leaf_27_clk _0110_ vssd1 vssd1 vccd1 vccd1 lcdPlayer.cnt_20ms\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_3065_ clknet_leaf_15_clk _0058_ _0027_ vssd1 vssd1 vccd1 vccd1 dispFSM.msg\[0\]
+ sky130_fd_sc_hd__dfstp_2
X_2016_ hostdisp.curr_guesses\[30\] net94 net79 net500 vssd1 vssd1 vccd1 vccd1 hostdisp.next_curr_guesses\[22\]
+ sky130_fd_sc_hd__o22a_1
XANTENNA__2085__A2 net97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_148 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_147_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_174_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_147_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2918_ dispFSM.guesses\[58\] net84 net61 net550 vssd1 vssd1 vccd1 vccd1 _0285_ sky130_fd_sc_hd__o22a_1
XFILLER_0_70_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1596__A1 net4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_30_clk clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_30_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_115_264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2849_ _0822_ _1379_ _1381_ net454 vssd1 vssd1 vccd1 vccd1 _0226_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA_fanout206_X net206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold130 hostdisp.next_curr_guesses\[39\] vssd1 vssd1 vccd1 vccd1 net394 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold152 _0163_ vssd1 vssd1 vccd1 vccd1 net416 sky130_fd_sc_hd__dlygate4sd3_1
Xhold141 dispFSM.guesses\[3\] vssd1 vssd1 vccd1 vccd1 net405 sky130_fd_sc_hd__dlygate4sd3_1
Xhold174 clock_div.next_count\[1\] vssd1 vssd1 vccd1 vccd1 net438 sky130_fd_sc_hd__dlygate4sd3_1
Xhold185 clock_div.count\[24\] vssd1 vssd1 vccd1 vccd1 net449 sky130_fd_sc_hd__dlygate4sd3_1
Xhold163 lcdPlayer.cnt_20ms\[14\] vssd1 vssd1 vccd1 vccd1 net427 sky130_fd_sc_hd__dlygate4sd3_1
Xhold196 dispFSM.guesses\[71\] vssd1 vssd1 vccd1 vccd1 net460 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3440__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_21_clk clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_21_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_36_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_151 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_136_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_324 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_234 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2000__A2 net94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2536__B1 _1097_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_188_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_9_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_182_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_106_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_12_clk clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_12_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_42_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2703_ gamelogic.letter\[1\] _0389_ gamelogic.setWord\[18\] _0379_ vssd1 vssd1 vccd1
+ vccd1 _1267_ sky130_fd_sc_hd__o22a_1
XFILLER_0_54_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2634_ dispFSM.guesses\[70\] _1072_ net105 dispFSM.guesses\[22\] _1205_ vssd1 vssd1
+ vccd1 vccd1 _1206_ sky130_fd_sc_hd__a221o_1
X_2565_ net286 net107 _1140_ net183 vssd1 vssd1 vccd1 vccd1 _0176_ sky130_fd_sc_hd__o211a_1
XANTENNA__2527__B1 _1104_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1516_ _0437_ _0443_ vssd1 vssd1 vccd1 vccd1 _0465_ sky130_fd_sc_hd__and2_1
XFILLER_0_10_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3313__CLK clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2496_ lcdPlayer.nextState\[5\] lcdPlayer.nextState\[4\] _1068_ vssd1 vssd1 vccd1
+ vccd1 _1074_ sky130_fd_sc_hd__nand3_2
X_1447_ net208 vssd1 vssd1 vccd1 vccd1 _0017_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_165_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3117_ clknet_leaf_34_clk _0104_ net158 vssd1 vssd1 vccd1 vccd1 uart_receiver.bit_index\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_179_234 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3463__CLK clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3048_ clknet_leaf_7_clk clock_div.next_count\[28\] net195 vssd1 vssd1 vccd1 vccd1
+ clock_div.count\[28\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_77_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_124_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_254 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_175 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3329__RESET_B net164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2949__A host_message_reg.Cstate vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout69_X net69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_183_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout80 _0825_ vssd1 vssd1 vccd1 vccd1 net80 sky130_fd_sc_hd__buf_2
XFILLER_0_126_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout91 net92 vssd1 vssd1 vccd1 vccd1 net91 sky130_fd_sc_hd__buf_2
XFILLER_0_153_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_153_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2350_ net167 _0943_ _0993_ _0955_ vssd1 vssd1 vccd1 vccd1 _0108_ sky130_fd_sc_hd__a31o_1
X_2281_ lcdPlayer.cnt_20ms\[20\] lcdPlayer.cnt_20ms\[19\] lcdPlayer.cnt_20ms\[18\]
+ lcdPlayer.cnt_20ms\[17\] vssd1 vssd1 vccd1 vccd1 _0950_ sky130_fd_sc_hd__or4b_1
XANTENNA__3486__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_1_clk clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_1_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_59_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2445__C1 _1034_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2460__A2 net75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1996_ hostdisp.curr_guesses\[10\] net92 net76 net410 vssd1 vssd1 vccd1 vccd1 hostdisp.next_curr_guesses\[2\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_15_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_171_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3597_ net157 vssd1 vssd1 vccd1 vccd1 net22 sky130_fd_sc_hd__clkbuf_1
X_2617_ net226 hostdisp.top\[77\] _1095_ vssd1 vssd1 vccd1 vccd1 _1190_ sky130_fd_sc_hd__o21a_1
X_2548_ net111 _1122_ _1124_ _1115_ _1121_ vssd1 vssd1 vccd1 vccd1 _1125_ sky130_fd_sc_hd__a2111o_1
X_2479_ lcdPlayer.nextState\[5\] lcdPlayer.nextState\[4\] vssd1 vssd1 vccd1 vccd1
+ _1058_ sky130_fd_sc_hd__or2_1
XFILLER_0_167_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2436__C1 net70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3209__CLK clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2451__A2 net67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_175_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload0 clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clkload0/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_80_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_133_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2978__B1 net50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_60_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1850_ clock_div.count\[23\] _0723_ net449 vssd1 vssd1 vccd1 vccd1 _0724_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_126_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_7_Left_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1477__B net6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1781_ _0401_ _0677_ _0679_ vssd1 vssd1 vccd1 vccd1 _0680_ sky130_fd_sc_hd__a21o_1
XFILLER_0_24_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3520_ clknet_leaf_2_clk hostdisp.next_curr_guesses\[2\] net180 vssd1 vssd1 vccd1
+ vccd1 hostdisp.curr_guesses\[2\] sky130_fd_sc_hd__dfstp_1
XFILLER_0_97_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3451_ clknet_leaf_13_clk _0329_ net198 vssd1 vssd1 vccd1 vccd1 gamelogic.setWord\[13\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_122_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3382_ clknet_leaf_22_clk _0271_ net188 vssd1 vssd1 vccd1 vccd1 dispFSM.guesses\[36\]
+ sky130_fd_sc_hd__dfstp_1
X_2402_ _0357_ _1025_ _1026_ vssd1 vssd1 vccd1 vccd1 _0127_ sky130_fd_sc_hd__a21oi_1
X_2333_ net74 _0984_ vssd1 vssd1 vccd1 vccd1 _0985_ sky130_fd_sc_hd__nor2_1
X_2264_ message_reg.state\[0\] _0370_ net89 vssd1 vssd1 vccd1 vccd1 _0941_ sky130_fd_sc_hd__and3b_2
XPHY_EDGE_ROW_127_Right_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1469__B1 net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2195_ net134 _0376_ vssd1 vssd1 vccd1 vccd1 _0900_ sky130_fd_sc_hd__nor2_1
XFILLER_0_79_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_189_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2969__B1 net49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3501__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_173_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_284 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1979_ _0365_ gamelogic.state\[2\] vssd1 vssd1 vccd1 vccd1 _0812_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout119_X net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold23 lcdPlayer.cnt_500hz\[15\] vssd1 vssd1 vccd1 vccd1 net287 sky130_fd_sc_hd__dlygate4sd3_1
Xhold12 lcdPlayer.cnt_500hz\[0\] vssd1 vssd1 vccd1 vccd1 net276 sky130_fd_sc_hd__dlygate4sd3_1
Xhold45 hostdisp.top\[52\] vssd1 vssd1 vccd1 vccd1 net309 sky130_fd_sc_hd__dlygate4sd3_1
Xhold56 lcdPlayer.cnt_500hz\[16\] vssd1 vssd1 vccd1 vccd1 net320 sky130_fd_sc_hd__dlygate4sd3_1
Xhold34 _0072_ vssd1 vssd1 vccd1 vccd1 net298 sky130_fd_sc_hd__dlygate4sd3_1
Xhold78 keypadFSMPlayer.prev_key\[3\] vssd1 vssd1 vccd1 vccd1 net342 sky130_fd_sc_hd__dlygate4sd3_1
Xhold89 uart_transmitter.clk_count\[7\] vssd1 vssd1 vccd1 vccd1 net353 sky130_fd_sc_hd__dlygate4sd3_1
Xhold67 hostdisp.top\[65\] vssd1 vssd1 vccd1 vccd1 net331 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_180_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3181__CLK clknet_leaf_30_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1578__A dispFSM.msg\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2173__S net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3566__Q hostdisp.Cstate vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_191_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_150_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_89_Left_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3524__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_98_Left_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_190_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2951_ net104 net55 vssd1 vssd1 vccd1 vccd1 _1394_ sky130_fd_sc_hd__nor2_4
XFILLER_0_139_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1902_ lcdPlayer.cnt_500hz\[5\] lcdPlayer.cnt_500hz\[7\] lcdPlayer.cnt_500hz\[6\]
+ vssd1 vssd1 vccd1 vccd1 _0755_ sky130_fd_sc_hd__or3_1
X_2882_ dispFSM.guesses\[22\] net87 net62 net562 vssd1 vssd1 vccd1 vccd1 _0249_ sky130_fd_sc_hd__o22a_1
XFILLER_0_120_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_0_clk_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1833_ net379 _0712_ _0693_ vssd1 vssd1 vccd1 vccd1 _0715_ sky130_fd_sc_hd__o21ai_1
X_1764_ _0665_ vssd1 vssd1 vccd1 vccd1 _0666_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3503_ clknet_leaf_30_clk hostdisp.next_curr_word\[25\] net173 vssd1 vssd1 vccd1
+ vccd1 hostdisp.curr_word\[25\] sky130_fd_sc_hd__dfstp_1
X_3434_ clknet_leaf_17_clk _0013_ _0041_ vssd1 vssd1 vccd1 vccd1 keypadFSMPlayer.state\[2\]
+ sky130_fd_sc_hd__dfrtp_2
X_1695_ keypadFSMHost.state\[1\] _0612_ _0613_ vssd1 vssd1 vccd1 vccd1 _0614_ sky130_fd_sc_hd__or3_1
XFILLER_0_148_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkload18_A clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3365_ clknet_leaf_24_clk _0254_ net183 vssd1 vssd1 vccd1 vccd1 dispFSM.guesses\[19\]
+ sky130_fd_sc_hd__dfstp_1
X_3296_ clknet_leaf_34_clk uart_receiver.next_state\[1\] net158 vssd1 vssd1 vccd1
+ vccd1 uart_receiver.state\[1\] sky130_fd_sc_hd__dfrtp_1
X_2316_ net74 _0973_ vssd1 vssd1 vccd1 vccd1 _0974_ sky130_fd_sc_hd__nor2_1
X_2247_ net230 _0546_ _0693_ vssd1 vssd1 vccd1 vccd1 _0937_ sky130_fd_sc_hd__or3_2
XFILLER_0_164_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout183_A net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2654__A2 _1078_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2178_ gamelogic.setWord\[23\] _0891_ net136 vssd1 vssd1 vccd1 vccd1 hostdisp.nextBottom\[71\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_189_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_116 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput13 net13 vssd1 vssd1 vccd1 vccd1 gpio_oeb[16] sky130_fd_sc_hd__buf_2
Xoutput24 net157 vssd1 vssd1 vccd1 vccd1 gpio_oeb[32] sky130_fd_sc_hd__buf_2
Xoutput35 net35 vssd1 vssd1 vccd1 vccd1 gpio_out[18] sky130_fd_sc_hd__buf_2
Xoutput46 net46 vssd1 vssd1 vccd1 vccd1 gpio_out[9] sky130_fd_sc_hd__buf_2
XANTENNA_fanout96_A _0626_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3547__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_2_clk_A clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3525__RESET_B net206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_19_Right_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_168_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_183_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_139_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2030__B1 net77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3077__CLK clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_28_Right_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1480_ net232 _0428_ vssd1 vssd1 vccd1 vccd1 _0432_ sky130_fd_sc_hd__nand2_1
XFILLER_0_94_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3150_ clknet_leaf_26_clk _0126_ vssd1 vssd1 vccd1 vccd1 lcdPlayer.cnt_20ms\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_3081_ clknet_leaf_33_clk _0071_ net160 vssd1 vssd1 vccd1 vccd1 buffer.temp_guess\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_2101_ hostdisp.curr_word\[32\] net99 net75 _0852_ gamelogic.indexCorrect\[4\] vssd1
+ vssd1 vccd1 vccd1 _0854_ sky130_fd_sc_hd__o2111a_1
X_2032_ hostdisp.curr_guesses\[46\] net94 net79 net465 vssd1 vssd1 vccd1 vccd1 hostdisp.next_curr_guesses\[38\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_168_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_109_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_37_Right_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_159_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_186_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2934_ dispFSM.guesses\[74\] net83 net61 net480 vssd1 vssd1 vccd1 vccd1 _0301_ sky130_fd_sc_hd__o22a_1
XFILLER_0_17_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2865_ net66 _1389_ vssd1 vssd1 vccd1 vccd1 _0234_ sky130_fd_sc_hd__and2_1
X_1816_ _0693_ _0702_ _0704_ vssd1 vssd1 vccd1 vccd1 clock_div.next_count\[9\] sky130_fd_sc_hd__and3_1
XFILLER_0_4_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_46_Right_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_142_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_107 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold301 hostdisp.top\[79\] vssd1 vssd1 vccd1 vccd1 net565 sky130_fd_sc_hd__dlygate4sd3_1
X_2796_ _0364_ gamelogic.state\[1\] gamelogic.state\[2\] _1248_ gamelogic.state\[3\]
+ vssd1 vssd1 vccd1 vccd1 _1342_ sky130_fd_sc_hd__a311o_1
X_1747_ uart_receiver.clk_count\[6\] _0649_ uart_receiver.clk_count\[7\] vssd1 vssd1
+ vccd1 vccd1 _0653_ sky130_fd_sc_hd__a21o_1
X_1678_ _0559_ _0599_ _0556_ vssd1 vssd1 vccd1 vccd1 _0601_ sky130_fd_sc_hd__a21oi_4
X_3417_ clknet_leaf_21_clk _0306_ net210 vssd1 vssd1 vccd1 vccd1 dispFSM.guesses\[71\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3348_ clknet_leaf_24_clk _0237_ net188 vssd1 vssd1 vccd1 vccd1 dispFSM.guesses\[2\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_0_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_175_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_168_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3279_ clknet_leaf_14_clk hostdisp.nextBottom\[77\] net207 vssd1 vssd1 vccd1 vccd1
+ hostdisp.bottom\[77\] sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_55_Right_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2088__B1 net75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_192_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_64_Right_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_210 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3611__242 vssd1 vssd1 vccd1 vccd1 _3611__242/HI net242 sky130_fd_sc_hd__conb_1
XANTENNA__2563__B2 net108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_73_Right_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_186_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_82_Right_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_183_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_130 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2650_ hostdisp.top\[47\] _1098_ _1217_ _1220_ net226 vssd1 vssd1 vccd1 vccd1 _1221_
+ sky130_fd_sc_hd__a2111o_1
X_1601_ keypadFSMPlayer.unlocked keypadplayer.scan_col\[0\] net154 _0536_ net332 vssd1
+ vssd1 vccd1 vccd1 _0050_ sky130_fd_sc_hd__a32o_1
XANTENNA__2003__B1 net79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_156_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2581_ lcdPlayer.nextState\[3\] _1059_ _1057_ lcdPlayer.nextState\[2\] vssd1 vssd1
+ vccd1 vccd1 _1156_ sky130_fd_sc_hd__o211a_1
X_1532_ keypadFSMPlayer.prev_key\[3\] _0361_ net155 vssd1 vssd1 vccd1 vccd1 _0480_
+ sky130_fd_sc_hd__or3b_1
X_1463_ net146 net147 vssd1 vssd1 vccd1 vccd1 _0415_ sky130_fd_sc_hd__or2_2
XFILLER_0_129_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3202_ clknet_leaf_24_clk _0178_ vssd1 vssd1 vccd1 vccd1 net29 sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_91_Right_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3133_ clknet_leaf_27_clk _0109_ vssd1 vssd1 vccd1 vccd1 lcdPlayer.cnt_20ms\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_179_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3064_ clknet_leaf_15_clk _0057_ _0026_ vssd1 vssd1 vccd1 vccd1 keypadFSMPlayer.prev_key\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_145_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2015_ net391 net95 net80 net400 vssd1 vssd1 vccd1 vccd1 hostdisp.next_curr_guesses\[21\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_159_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_174_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_159_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3242__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2917_ dispFSM.guesses\[57\] net86 net62 net563 vssd1 vssd1 vccd1 vccd1 _0284_ sky130_fd_sc_hd__o22a_1
XFILLER_0_9_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_118_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2848_ _1380_ _1381_ vssd1 vssd1 vccd1 vccd1 _0225_ sky130_fd_sc_hd__and2_1
X_2779_ host_message_reg.setLetter\[2\] _1290_ _1329_ _1330_ vssd1 vssd1 vccd1 vccd1
+ _0207_ sky130_fd_sc_hd__o22a_1
XFILLER_0_115_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold120 dispFSM.guesses\[47\] vssd1 vssd1 vccd1 vccd1 net384 sky130_fd_sc_hd__dlygate4sd3_1
Xhold142 dispFSM.guesses\[23\] vssd1 vssd1 vccd1 vccd1 net406 sky130_fd_sc_hd__dlygate4sd3_1
Xhold131 dispFSM.guesses\[21\] vssd1 vssd1 vccd1 vccd1 net395 sky130_fd_sc_hd__dlygate4sd3_1
Xhold153 lcdPlayer.cnt_20ms\[17\] vssd1 vssd1 vccd1 vccd1 net417 sky130_fd_sc_hd__dlygate4sd3_1
Xhold186 dispFSM.guesses\[31\] vssd1 vssd1 vccd1 vccd1 net450 sky130_fd_sc_hd__dlygate4sd3_1
Xhold175 hostdisp.curr_guesses\[23\] vssd1 vssd1 vccd1 vccd1 net439 sky130_fd_sc_hd__dlygate4sd3_1
Xhold164 hostdisp.curr_guesses\[47\] vssd1 vssd1 vccd1 vccd1 net428 sky130_fd_sc_hd__dlygate4sd3_1
Xhold197 clock_div.count\[4\] vssd1 vssd1 vccd1 vccd1 net461 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_186_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_129_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2446__S net67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout59_A _1391_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_165_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_52_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2784__B2 host_message_reg.setLetter\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_136_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2536__A1 hostdisp.bottom\[49\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_246 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_188_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3265__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_25_Left_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_379 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_171_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2702_ _0384_ gamelogic.setWord\[21\] gamelogic.setWord\[22\] _0385_ _1265_ vssd1
+ vssd1 vccd1 vccd1 _1266_ sky130_fd_sc_hd__a221o_1
XFILLER_0_42_325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2633_ dispFSM.guesses\[30\] net115 _1086_ dispFSM.guesses\[78\] vssd1 vssd1 vccd1
+ vccd1 _1205_ sky130_fd_sc_hd__a22o_1
XFILLER_0_2_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2564_ _0764_ _1131_ _1137_ _1139_ vssd1 vssd1 vccd1 vccd1 _1140_ sky130_fd_sc_hd__or4_1
X_1515_ _0459_ _0463_ _0464_ _0457_ vssd1 vssd1 vccd1 vccd1 _0064_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_10_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_34_Left_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2495_ net138 _0356_ vssd1 vssd1 vccd1 vccd1 _1073_ sky130_fd_sc_hd__or2_1
X_1446_ net442 vssd1 vssd1 vccd1 vccd1 _0400_ sky130_fd_sc_hd__inv_2
XFILLER_0_156_42 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2477__D _0822_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_165_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3116_ clknet_leaf_19_clk uart_transmitter.next_state\[2\] net210 vssd1 vssd1 vccd1
+ vccd1 uart_transmitter.state\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_65_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_179_246 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3047_ clknet_leaf_7_clk clock_div.next_count\[27\] net195 vssd1 vssd1 vccd1 vccd1
+ clock_div.count\[27\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_124_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_43_Left_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_266 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_176_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_269 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3511__SET_B net164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_52_Left_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3369__RESET_B net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3288__CLK clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_183_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_61_Left_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_185_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_193_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2757__A1 host_message_reg.setLetter\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout70 net71 vssd1 vssd1 vccd1 vccd1 net70 sky130_fd_sc_hd__buf_2
XFILLER_0_36_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout81 net82 vssd1 vssd1 vccd1 vccd1 net81 sky130_fd_sc_hd__buf_2
Xfanout92 _0824_ vssd1 vssd1 vccd1 vccd1 net92 sky130_fd_sc_hd__clkbuf_4
XANTENNA__2205__A net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_108_Right_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_70_Left_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_153_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2280_ lcdPlayer.cnt_20ms\[15\] lcdPlayer.cnt_20ms\[14\] lcdPlayer.cnt_20ms\[13\]
+ lcdPlayer.cnt_20ms\[16\] vssd1 vssd1 vccd1 vccd1 _0949_ sky130_fd_sc_hd__or4b_1
XFILLER_0_193_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1995_ hostdisp.curr_guesses\[9\] net94 net78 net436 vssd1 vssd1 vccd1 vccd1 hostdisp.next_curr_guesses\[1\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_125_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2616_ net226 hostdisp.top\[45\] _1098_ vssd1 vssd1 vccd1 vccd1 _1189_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_171_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3596_ net156 vssd1 vssd1 vccd1 vccd1 net21 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3430__CLK clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2547_ lcdPlayer.nextState\[2\] _0356_ _1123_ _0758_ _0752_ vssd1 vssd1 vccd1 vccd1
+ _1124_ sky130_fd_sc_hd__a311o_1
XFILLER_0_55_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2478_ lcdPlayer.nextState\[5\] lcdPlayer.nextState\[4\] vssd1 vssd1 vccd1 vccd1
+ _1057_ sky130_fd_sc_hd__nor2_1
X_1429_ gamelogic.setWord\[37\] vssd1 vssd1 vccd1 vccd1 _0383_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_183_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2436__B1 _0828_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_182_208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload1 clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clkload1/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_33_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_143_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_374 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2124__C1 net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1780_ uart_transmitter.bit_index\[1\] _0678_ uart_transmitter.bit_index\[2\] vssd1
+ vssd1 vccd1 vccd1 _0679_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_24_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_188_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3453__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3450_ clknet_leaf_3_clk _0328_ net177 vssd1 vssd1 vccd1 vccd1 gamelogic.setWord\[12\]
+ sky130_fd_sc_hd__dfstp_1
X_2401_ lcdPlayer.cnt_20ms\[20\] lcdPlayer.cnt_20ms\[19\] _1022_ _0017_ vssd1 vssd1
+ vccd1 vccd1 _1026_ sky130_fd_sc_hd__a31o_1
X_3381_ clknet_leaf_25_clk _0270_ net183 vssd1 vssd1 vccd1 vccd1 dispFSM.guesses\[35\]
+ sky130_fd_sc_hd__dfstp_1
X_2332_ lcdPlayer.cnt_500hz\[17\] lcdPlayer.cnt_500hz\[16\] _0980_ vssd1 vssd1 vccd1
+ vccd1 _0984_ sky130_fd_sc_hd__and3_1
XFILLER_0_41_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2263_ keypadFSMPlayer.state\[4\] keypadFSMPlayer.state\[0\] _0444_ _0446_ vssd1
+ vssd1 vccd1 vccd1 _0940_ sky130_fd_sc_hd__or4_4
XFILLER_0_137_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_108_Left_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_42 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1469__A1 net4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2194_ gamelogic.setWord\[31\] _0899_ net133 vssd1 vssd1 vccd1 vccd1 hostdisp.nextBottom\[79\]
+ sky130_fd_sc_hd__mux2_1
XANTENNA__2130__A2 net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2418__B1 net69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_121_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_157_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_117_Left_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_173_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1978_ _0618_ _0811_ vssd1 vssd1 vccd1 vccd1 uart_receiver.temp_byte\[7\] sky130_fd_sc_hd__and2_1
XANTENNA_fanout226_A net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_294 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3579_ net156 vssd1 vssd1 vccd1 vccd1 net11 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_126_Left_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold13 hostdisp.top\[45\] vssd1 vssd1 vccd1 vccd1 net277 sky130_fd_sc_hd__dlygate4sd3_1
Xhold24 clock_div.count\[6\] vssd1 vssd1 vccd1 vccd1 net288 sky130_fd_sc_hd__dlygate4sd3_1
Xhold46 lcdPlayer.cnt_500hz\[20\] vssd1 vssd1 vccd1 vccd1 net310 sky130_fd_sc_hd__dlygate4sd3_1
Xhold35 net32 vssd1 vssd1 vccd1 vccd1 net299 sky130_fd_sc_hd__dlygate4sd3_1
Xhold68 keypadFSMPlayer.prev_key\[0\] vssd1 vssd1 vccd1 vccd1 net332 sky130_fd_sc_hd__dlygate4sd3_1
Xhold57 dispFSM.guesses\[5\] vssd1 vssd1 vccd1 vccd1 net321 sky130_fd_sc_hd__dlygate4sd3_1
Xhold79 hostdisp.top\[68\] vssd1 vssd1 vccd1 vccd1 net343 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_180_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3326__CLK clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3476__CLK clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_193_Right_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_191_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2042__X _0827_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2648__B1 net108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_186_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2950_ host_message_reg.Cstate keypadFSMHost.state\[4\] keypadFSMHost.state\[0\]
+ _0595_ vssd1 vssd1 vccd1 vccd1 _1393_ sky130_fd_sc_hd__or4_2
XFILLER_0_29_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2881_ net395 net90 net64 net446 vssd1 vssd1 vccd1 vccd1 _0248_ sky130_fd_sc_hd__a22o_1
X_1901_ lcdPlayer.cnt_500hz\[15\] lcdPlayer.cnt_500hz\[20\] _0753_ vssd1 vssd1 vccd1
+ vccd1 _0754_ sky130_fd_sc_hd__or3_1
X_1832_ clock_div.count\[13\] clock_div.count\[14\] _0685_ _0709_ vssd1 vssd1 vccd1
+ vccd1 _0714_ sky130_fd_sc_hd__and4_1
XFILLER_0_123_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_160_Right_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1763_ uart_transmitter.bit_index\[1\] uart_transmitter.bit_index\[0\] _0664_ vssd1
+ vssd1 vccd1 vccd1 _0665_ sky130_fd_sc_hd__and3_1
XFILLER_0_40_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1694_ _0583_ _0584_ _0369_ vssd1 vssd1 vccd1 vccd1 _0613_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_52_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3502_ clknet_leaf_3_clk hostdisp.next_curr_word\[24\] net172 vssd1 vssd1 vccd1 vccd1
+ hostdisp.curr_word\[24\] sky130_fd_sc_hd__dfstp_1
X_3433_ clknet_leaf_17_clk _0012_ _0040_ vssd1 vssd1 vccd1 vccd1 keypadFSMPlayer.state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3589__261 vssd1 vssd1 vccd1 vccd1 net261 _3589__261/LO sky130_fd_sc_hd__conb_1
X_3364_ clknet_leaf_24_clk _0253_ net187 vssd1 vssd1 vccd1 vccd1 dispFSM.guesses\[18\]
+ sky130_fd_sc_hd__dfstp_1
X_3295_ clknet_leaf_34_clk uart_receiver.next_state\[0\] net158 vssd1 vssd1 vccd1
+ vccd1 uart_receiver.state\[0\] sky130_fd_sc_hd__dfstp_1
X_2315_ lcdPlayer.cnt_500hz\[11\] _0971_ vssd1 vssd1 vccd1 vccd1 _0973_ sky130_fd_sc_hd__and2_1
X_2246_ net230 _0693_ vssd1 vssd1 vccd1 vccd1 _0936_ sky130_fd_sc_hd__nor2_1
XANTENNA__2639__B1 _1096_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3349__CLK clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2177_ gamelogic.setWord\[31\] hostdisp.curr_guesses\[31\] net126 vssd1 vssd1 vccd1
+ vccd1 _0891_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout176_A net179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3499__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_128 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2811__B1 _1275_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_180_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2590__A2 net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput14 net14 vssd1 vssd1 vccd1 vccd1 gpio_oeb[17] sky130_fd_sc_hd__buf_2
Xoutput25 net25 vssd1 vssd1 vccd1 vccd1 gpio_oeb[6] sky130_fd_sc_hd__buf_2
Xoutput36 net36 vssd1 vssd1 vccd1 vccd1 gpio_out[25] sky130_fd_sc_hd__buf_2
XFILLER_0_3_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3605__239 vssd1 vssd1 vccd1 vccd1 _3605__239/HI net239 sky130_fd_sc_hd__conb_1
XFILLER_0_58_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_168_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_150 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_191_380 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_139_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3080_ clknet_leaf_35_clk net280 net161 vssd1 vssd1 vccd1 vccd1 buffer.temp_guess\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_2100_ hostdisp.curr_word\[33\] hostdisp.curr_word\[34\] hostdisp.curr_word\[35\]
+ _0412_ net99 vssd1 vssd1 vccd1 vccd1 _0853_ sky130_fd_sc_hd__a41o_1
X_2031_ net401 net95 _0825_ net431 vssd1 vssd1 vccd1 vccd1 hostdisp.next_curr_guesses\[37\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_27_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_109_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2097__B2 gamelogic.letter\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_186_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2933_ dispFSM.guesses\[73\] net86 net63 net536 vssd1 vssd1 vccd1 vccd1 _0300_ sky130_fd_sc_hd__o22a_1
XFILLER_0_57_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2864_ net140 buffer.temp_guess\[7\] _0918_ vssd1 vssd1 vccd1 vccd1 _1389_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1815_ _0703_ vssd1 vssd1 vccd1 vccd1 _0704_ sky130_fd_sc_hd__inv_2
XFILLER_0_150_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2795_ host_message_reg.setLetter\[7\] _1336_ vssd1 vssd1 vccd1 vccd1 _0212_ sky130_fd_sc_hd__and2_1
XFILLER_0_142_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold302 gamelogic.setWord\[5\] vssd1 vssd1 vccd1 vccd1 net566 sky130_fd_sc_hd__dlygate4sd3_1
X_1746_ net323 _0649_ _0652_ vssd1 vssd1 vccd1 vccd1 uart_receiver.next_clk_count\[6\]
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_102_119 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2572__A2 net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1677_ _0599_ vssd1 vssd1 vccd1 vccd1 _0600_ sky130_fd_sc_hd__inv_2
XFILLER_0_110_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3416_ clknet_leaf_20_clk _0305_ net203 vssd1 vssd1 vccd1 vccd1 dispFSM.guesses\[70\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_0_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_90_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3171__CLK clknet_leaf_30_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3347_ clknet_leaf_21_clk _0236_ net204 vssd1 vssd1 vccd1 vccd1 dispFSM.guesses\[1\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_168_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3278_ clknet_leaf_3_clk hostdisp.nextBottom\[76\] net177 vssd1 vssd1 vccd1 vccd1
+ hostdisp.bottom\[76\] sky130_fd_sc_hd__dfrtp_1
X_2229_ _0364_ _0923_ vssd1 vssd1 vccd1 vccd1 _0924_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout179_X net179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_191_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_192_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_179_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_288 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3514__CLK clknet_leaf_31_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_186_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2079__B2 gamelogic.letter\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_55_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3044__CLK clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_30_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1600_ net367 net148 _0535_ vssd1 vssd1 vccd1 vccd1 _0051_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_156_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3194__CLK clknet_leaf_31_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2554__A2 net114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2580_ _1061_ _1075_ _1094_ vssd1 vssd1 vccd1 vccd1 _1155_ sky130_fd_sc_hd__or3_1
X_1531_ keypadFSMPlayer.prev_key\[4\] _0425_ vssd1 vssd1 vccd1 vccd1 _0479_ sky130_fd_sc_hd__xor2_1
X_1462_ net146 net147 vssd1 vssd1 vccd1 vccd1 _0414_ sky130_fd_sc_hd__nor2_1
XFILLER_0_1_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3201_ clknet_leaf_25_clk _0177_ vssd1 vssd1 vccd1 vccd1 net46 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_180_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3132_ clknet_leaf_27_clk _0108_ vssd1 vssd1 vccd1 vccd1 lcdPlayer.cnt_20ms\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_3063_ clknet_leaf_16_clk _0056_ _0025_ vssd1 vssd1 vccd1 vccd1 keypadFSMPlayer.prev_key\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_2014_ hostdisp.curr_guesses\[28\] net92 net77 net489 vssd1 vssd1 vccd1 vccd1 hostdisp.next_curr_guesses\[20\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_89_264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_159_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_174_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_162_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2916_ dispFSM.guesses\[56\] net81 net56 net459 vssd1 vssd1 vccd1 vccd1 _0283_ sky130_fd_sc_hd__o22a_1
XFILLER_0_155_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2847_ _0821_ _1379_ _1378_ vssd1 vssd1 vccd1 vccd1 _1381_ sky130_fd_sc_hd__a21o_1
XFILLER_0_72_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2778_ host_message_reg.setLetter\[2\] _0601_ _1310_ _0597_ vssd1 vssd1 vccd1 vccd1
+ _1330_ sky130_fd_sc_hd__a211o_1
Xhold110 _0272_ vssd1 vssd1 vccd1 vccd1 net374 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_2_1__f_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold121 _0274_ vssd1 vssd1 vccd1 vccd1 net385 sky130_fd_sc_hd__dlygate4sd3_1
Xhold143 _0258_ vssd1 vssd1 vccd1 vccd1 net407 sky130_fd_sc_hd__dlygate4sd3_1
Xhold132 _0256_ vssd1 vssd1 vccd1 vccd1 net396 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_1_clk_A clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1729_ _0627_ _0637_ _0640_ _0641_ vssd1 vssd1 vccd1 vccd1 _0642_ sky130_fd_sc_hd__o31a_1
XFILLER_0_79_94 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold165 clock_div.count\[15\] vssd1 vssd1 vccd1 vccd1 net429 sky130_fd_sc_hd__dlygate4sd3_1
Xhold176 clock_div.count\[27\] vssd1 vssd1 vccd1 vccd1 net440 sky130_fd_sc_hd__dlygate4sd3_1
Xhold154 lcdPlayer.cnt_20ms\[16\] vssd1 vssd1 vccd1 vccd1 net418 sky130_fd_sc_hd__dlygate4sd3_1
Xhold198 hostdisp.curr_guesses\[33\] vssd1 vssd1 vccd1 vccd1 net462 sky130_fd_sc_hd__dlygate4sd3_1
Xhold187 _0266_ vssd1 vssd1 vccd1 vccd1 net451 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3067__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_52_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_258 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2536__A2 net114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_188_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_147_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2701_ _0382_ gamelogic.setWord\[20\] vssd1 vssd1 vccd1 vccd1 _1265_ sky130_fd_sc_hd__nor2_1
XFILLER_0_42_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2632_ dispFSM.guesses\[62\] net117 _1084_ dispFSM.guesses\[6\] vssd1 vssd1 vccd1
+ vccd1 _1204_ sky130_fd_sc_hd__a22o_1
X_2563_ lcdPlayer.nextState\[2\] _1123_ _1138_ net108 vssd1 vssd1 vccd1 vccd1 _1139_
+ sky130_fd_sc_hd__a22o_1
X_1514_ _0444_ _0445_ vssd1 vssd1 vccd1 vccd1 _0464_ sky130_fd_sc_hd__nor2_1
XFILLER_0_120_291 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2494_ _1070_ _1071_ vssd1 vssd1 vccd1 vccd1 _1072_ sky130_fd_sc_hd__nor2_4
X_1445_ uart_transmitter.state\[1\] vssd1 vssd1 vccd1 vccd1 _0399_ sky130_fd_sc_hd__inv_2
XFILLER_0_10_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3115_ clknet_leaf_20_clk uart_transmitter.next_state\[1\] net210 vssd1 vssd1 vccd1
+ vccd1 uart_transmitter.state\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_4_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3046_ clknet_leaf_7_clk clock_div.next_count\[26\] net195 vssd1 vssd1 vccd1 vccd1
+ clock_div.count\[26\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_179_258 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_124_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_176_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2949__C keypadFSMHost.state\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_183_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2206__A1 net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout60 net63 vssd1 vssd1 vccd1 vccd1 net60 sky130_fd_sc_hd__buf_2
Xfanout71 _1032_ vssd1 vssd1 vccd1 vccd1 net71 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_36_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout82 _0940_ vssd1 vssd1 vccd1 vccd1 net82 sky130_fd_sc_hd__buf_2
XFILLER_0_153_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2205__B gamelogic.setWord\[37\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout93 net94 vssd1 vssd1 vccd1 vccd1 net93 sky130_fd_sc_hd__buf_2
XFILLER_0_119_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_153_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3382__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2445__B2 _0830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2445__A1 net130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1994_ hostdisp.curr_guesses\[8\] net93 net78 net420 vssd1 vssd1 vccd1 vccd1 hostdisp.next_curr_guesses\[0\]
+ sky130_fd_sc_hd__o22a_1
XANTENNA_clkbuf_leaf_14_clk_X clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2115__B net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload30 clknet_leaf_18_clk vssd1 vssd1 vccd1 vccd1 clkload30/Y sky130_fd_sc_hd__inv_6
X_2615_ hostdisp.bottom\[101\] dispFSM.guesses\[5\] net228 vssd1 vssd1 vccd1 vccd1
+ _1188_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_171_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3595_ net156 vssd1 vssd1 vccd1 vccd1 net20 sky130_fd_sc_hd__clkbuf_1
XANTENNA_clkbuf_leaf_29_clk_X clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_386 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2546_ lcdPlayer.nextState\[3\] lcdPlayer.nextState\[1\] _1057_ vssd1 vssd1 vccd1
+ vccd1 _1123_ sky130_fd_sc_hd__and3b_1
X_2477_ net129 net357 net103 _0822_ vssd1 vssd1 vccd1 vccd1 _0172_ sky130_fd_sc_hd__or4_1
X_1428_ net142 vssd1 vssd1 vccd1 vccd1 _0382_ sky130_fd_sc_hd__inv_2
XFILLER_0_48_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2684__A1 gamelogic.indexCorrect\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3029_ clknet_leaf_7_clk clock_div.next_count\[9\] net214 vssd1 vssd1 vccd1 vccd1
+ clock_div.count\[9\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__2436__A1 net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_174_Right_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_190_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload2 clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clkload2/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_73_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2187__S net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2427__B2 _0828_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_141_Right_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_60_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_181_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2503__X _1081_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2400_ net168 _1024_ _1025_ vssd1 vssd1 vccd1 vccd1 _0126_ sky130_fd_sc_hd__and3_1
X_3380_ clknet_leaf_24_clk _0269_ net189 vssd1 vssd1 vccd1 vccd1 dispFSM.guesses\[34\]
+ sky130_fd_sc_hd__dfstp_1
X_2331_ net320 _0980_ _0983_ vssd1 vssd1 vccd1 vccd1 _0099_ sky130_fd_sc_hd__o21a_1
X_2262_ _0372_ _0374_ _0443_ _0445_ vssd1 vssd1 vccd1 vccd1 _0939_ sky130_fd_sc_hd__and4_1
X_2193_ gamelogic.setWord\[39\] hostdisp.curr_guesses\[39\] net126 vssd1 vssd1 vccd1
+ vccd1 _0899_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_54 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2969__A2 net53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2418__B2 hostdisp.top\[44\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_157_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_121_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2126__A net130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_173_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3278__CLK clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1977_ buffer.Rx_byte\[7\] net2 _0623_ vssd1 vssd1 vccd1 vccd1 _0811_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout121_A net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout219_A net221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3578_ net156 vssd1 vssd1 vccd1 vccd1 net10 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_93_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2529_ hostdisp.top\[56\] dispFSM.msg\[0\] net226 vssd1 vssd1 vccd1 vccd1 _1107_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold14 lcdPlayer.cnt_20ms\[18\] vssd1 vssd1 vccd1 vccd1 net278 sky130_fd_sc_hd__dlygate4sd3_1
Xhold25 message_reg.msg\[6\] vssd1 vssd1 vccd1 vccd1 net289 sky130_fd_sc_hd__dlygate4sd3_1
Xhold36 buffer.Rx_byte\[2\] vssd1 vssd1 vccd1 vccd1 net300 sky130_fd_sc_hd__dlygate4sd3_1
Xhold47 gamelogic.red vssd1 vssd1 vccd1 vccd1 net311 sky130_fd_sc_hd__dlygate4sd3_1
Xhold69 _0050_ vssd1 vssd1 vccd1 vccd1 net333 sky130_fd_sc_hd__dlygate4sd3_1
Xhold58 _0240_ vssd1 vssd1 vccd1 vccd1 net322 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_39_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_22_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_191_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2593__B1 net110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_186_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_186_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2880_ dispFSM.guesses\[20\] net83 net60 net471 vssd1 vssd1 vccd1 vccd1 _0247_ sky130_fd_sc_hd__o22a_1
X_1900_ lcdPlayer.cnt_500hz\[17\] lcdPlayer.cnt_500hz\[16\] lcdPlayer.cnt_500hz\[19\]
+ lcdPlayer.cnt_500hz\[18\] vssd1 vssd1 vccd1 vccd1 _0753_ sky130_fd_sc_hd__or4_1
XFILLER_0_84_343 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1831_ net429 _0711_ _0713_ _0693_ vssd1 vssd1 vccd1 vccd1 clock_div.next_count\[15\]
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_44_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1762_ uart_transmitter.clk_count\[8\] uart_transmitter.clk_count\[9\] _0663_ uart_transmitter.clk_count\[10\]
+ vssd1 vssd1 vccd1 vccd1 _0664_ sky130_fd_sc_hd__o31a_1
XFILLER_0_114_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2584__B1 net106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1693_ keypadFSMHost.state\[0\] _0579_ _0580_ _0581_ vssd1 vssd1 vccd1 vccd1 _0612_
+ sky130_fd_sc_hd__or4_2
X_3501_ clknet_leaf_14_clk hostdisp.next_curr_word\[23\] net201 vssd1 vssd1 vccd1
+ vccd1 hostdisp.curr_word\[23\] sky130_fd_sc_hd__dfrtp_1
X_3432_ clknet_leaf_18_clk _0011_ _0039_ vssd1 vssd1 vccd1 vccd1 keypadFSMPlayer.state\[0\]
+ sky130_fd_sc_hd__dfstp_1
X_3363_ clknet_leaf_20_clk _0252_ net204 vssd1 vssd1 vccd1 vccd1 dispFSM.guesses\[17\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__3023__RESET_B net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2314_ lcdPlayer.cnt_500hz\[10\] _0969_ _0972_ _0956_ vssd1 vssd1 vccd1 vccd1 _0093_
+ sky130_fd_sc_hd__o211a_1
X_3294_ clknet_leaf_35_clk _0215_ net162 vssd1 vssd1 vccd1 vccd1 gamelogic.rights\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_2245_ keypadHostt.scan_col\[0\] net152 _0362_ _0363_ vssd1 vssd1 vccd1 vccd1 _0935_
+ sky130_fd_sc_hd__and4b_1
X_2176_ gamelogic.setWord\[22\] _0890_ net134 vssd1 vssd1 vccd1 vccd1 hostdisp.nextBottom\[70\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_189_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_164_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout169_A net225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_192_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_180_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2575__B1 net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_160_267 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput15 net15 vssd1 vssd1 vccd1 vccd1 gpio_oeb[18] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_1_Right_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput26 net26 vssd1 vssd1 vccd1 vccd1 gpio_oeb[7] sky130_fd_sc_hd__buf_2
Xoutput37 net37 vssd1 vssd1 vccd1 vccd1 gpio_out[26] sky130_fd_sc_hd__buf_2
XFILLER_0_11_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_183_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2030__A2 net92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3484__SET_B net164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2566__B1 _1098_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_172 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2500__Y _1078_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2030_ hostdisp.curr_guesses\[44\] net92 net77 net553 vssd1 vssd1 vccd1 vccd1 hostdisp.next_curr_guesses\[36\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_178_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_145_Left_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_109_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2849__A1_N _0822_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_186_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2932_ dispFSM.guesses\[72\] net82 net56 net483 vssd1 vssd1 vccd1 vccd1 _0299_ sky130_fd_sc_hd__o22a_1
XFILLER_0_186_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_162 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2863_ net66 _1388_ vssd1 vssd1 vccd1 vccd1 _0233_ sky130_fd_sc_hd__and2_1
X_1814_ clock_div.count\[7\] clock_div.count\[8\] clock_div.count\[9\] _0700_ vssd1
+ vssd1 vccd1 vccd1 _0703_ sky130_fd_sc_hd__and4_2
XPHY_EDGE_ROW_154_Left_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2794_ _0605_ _1340_ _1341_ _1289_ _1338_ vssd1 vssd1 vccd1 vccd1 _0211_ sky130_fd_sc_hd__a311o_1
XANTENNA__2123__B net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1745_ uart_receiver.clk_count\[6\] _0649_ _0641_ vssd1 vssd1 vccd1 vccd1 _0652_
+ sky130_fd_sc_hd__o21ai_1
XANTENNA__2557__B1 _1086_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold303 lcdPlayer.cnt_20ms\[3\] vssd1 vssd1 vccd1 vccd1 net567 sky130_fd_sc_hd__dlygate4sd3_1
X_1676_ keypadHostt.scan_col\[0\] net152 keypadHostt.scan_col\[3\] _0363_ vssd1 vssd1
+ vccd1 vccd1 _0599_ sky130_fd_sc_hd__or4_2
XFILLER_0_7_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3316__CLK clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3415_ clknet_leaf_21_clk _0304_ net202 vssd1 vssd1 vccd1 vccd1 dispFSM.guesses\[69\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_110_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_90_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3346_ clknet_leaf_25_clk _0235_ net182 vssd1 vssd1 vccd1 vccd1 dispFSM.guesses\[0\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_168_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_163_Left_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3466__CLK clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3277_ clknet_leaf_0_clk hostdisp.nextBottom\[75\] net170 vssd1 vssd1 vccd1 vccd1
+ hostdisp.bottom\[75\] sky130_fd_sc_hd__dfrtp_1
X_2228_ gamelogic.state\[1\] _0922_ vssd1 vssd1 vccd1 vccd1 _0923_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_127_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2159_ gamelogic.setWord\[22\] hostdisp.curr_guesses\[22\] net124 vssd1 vssd1 vccd1
+ vccd1 _0882_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_165_304 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_179_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_33_clk clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_33_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_192_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_180_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_172_Left_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_181_Left_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2720__B1 _0392_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_186_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_168_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_315 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_190_Left_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_168_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_24_clk clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_24_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_66_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2224__A net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2003__A2 net94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2539__B1 net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3339__CLK clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_176 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_156_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1530_ net146 net155 keypadFSMPlayer.prev_key\[3\] vssd1 vssd1 vccd1 vccd1 _0478_
+ sky130_fd_sc_hd__a21bo_1
XFILLER_0_22_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1461_ net1 vssd1 vssd1 vccd1 vccd1 net24 sky130_fd_sc_hd__inv_2
XANTENNA__3489__CLK clknet_leaf_30_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3200_ clknet_leaf_25_clk _0176_ vssd1 vssd1 vccd1 vccd1 net45 sky130_fd_sc_hd__dfxtp_1
X_3131_ clknet_leaf_27_clk _0107_ vssd1 vssd1 vccd1 vccd1 lcdPlayer.cnt_20ms\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_173_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3062_ clknet_leaf_12_clk _0055_ _0024_ vssd1 vssd1 vccd1 vccd1 keypadFSMPlayer.prev_key\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_145_34 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_43 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2475__C1 _1034_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2013_ hostdisp.curr_guesses\[27\] net91 net76 net544 vssd1 vssd1 vccd1 vccd1 hostdisp.next_curr_guesses\[19\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_159_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_174_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_15_clk clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_15_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_9_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2915_ net425 net88 net65 net384 vssd1 vssd1 vccd1 vccd1 _0282_ sky130_fd_sc_hd__a22o_1
XFILLER_0_45_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2846_ gamelogic.incorrect\[0\] _0821_ gamelogic.incorrect\[1\] vssd1 vssd1 vccd1
+ vccd1 _1380_ sky130_fd_sc_hd__a21o_1
XFILLER_0_170_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2777_ _1327_ _1328_ vssd1 vssd1 vccd1 vccd1 _1329_ sky130_fd_sc_hd__nor2_1
XFILLER_0_115_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold100 gamelogic.green vssd1 vssd1 vccd1 vccd1 net364 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_78_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold144 keypadFSMHost.prev_key\[0\] vssd1 vssd1 vccd1 vccd1 net408 sky130_fd_sc_hd__dlygate4sd3_1
Xhold111 clock_div.count\[3\] vssd1 vssd1 vccd1 vccd1 net375 sky130_fd_sc_hd__dlygate4sd3_1
Xhold122 keypadFSMPlayer.prev_key\[4\] vssd1 vssd1 vccd1 vccd1 net386 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout201_A net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1728_ _0633_ _0640_ vssd1 vssd1 vccd1 vccd1 _0641_ sky130_fd_sc_hd__or2_2
Xhold133 hostdisp.top\[40\] vssd1 vssd1 vccd1 vccd1 net397 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_73 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1659_ keypadFSMPlayer.state\[3\] _0452_ _0588_ _0451_ vssd1 vssd1 vccd1 vccd1 _0014_
+ sky130_fd_sc_hd__a22o_1
Xhold177 dispFSM.guesses\[15\] vssd1 vssd1 vccd1 vccd1 net441 sky130_fd_sc_hd__dlygate4sd3_1
Xhold166 dispFSM.guesses\[69\] vssd1 vssd1 vccd1 vccd1 net430 sky130_fd_sc_hd__dlygate4sd3_1
Xhold155 dispFSM.guesses\[2\] vssd1 vssd1 vccd1 vccd1 net419 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_186_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold199 hostdisp.curr_guesses\[25\] vssd1 vssd1 vccd1 vccd1 net463 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold188 lcdPlayer.cnt_500hz\[18\] vssd1 vssd1 vccd1 vccd1 net452 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_input6_A gpio_in[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_186_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_129_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1912__S net106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3329_ clknet_leaf_33_clk gamelogic.nextState\[3\] net164 vssd1 vssd1 vccd1 vccd1
+ gamelogic.state\[3\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_44_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_52_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2044__A net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_188_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_188_Right_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_147_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_224 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2472__A2 net73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2506__X _1084_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3161__CLK clknet_leaf_30_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2700_ net140 gamelogic.setWord\[23\] vssd1 vssd1 vccd1 vccd1 _1264_ sky130_fd_sc_hd__or2_1
X_2631_ dispFSM.guesses\[14\] _1078_ net110 dispFSM.guesses\[38\] vssd1 vssd1 vccd1
+ vccd1 _1203_ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2562_ hostdisp.top\[58\] dispFSM.msg\[2\] net227 vssd1 vssd1 vccd1 vccd1 _1138_
+ sky130_fd_sc_hd__mux2_1
X_1513_ _0455_ _0457_ _0462_ _0429_ vssd1 vssd1 vccd1 vccd1 _0463_ sky130_fd_sc_hd__o2bb2a_1
X_2493_ _1061_ _1068_ vssd1 vssd1 vccd1 vccd1 _1071_ sky130_fd_sc_hd__nand2_2
X_1444_ uart_transmitter.state\[0\] vssd1 vssd1 vccd1 vccd1 _0398_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_4_clk clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_4_clk
+ sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_155_Right_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3114_ clknet_leaf_19_clk uart_transmitter.next_state\[0\] net211 vssd1 vssd1 vccd1
+ vccd1 uart_transmitter.state\[0\] sky130_fd_sc_hd__dfstp_1
X_3045_ clknet_leaf_7_clk clock_div.next_count\[25\] net195 vssd1 vssd1 vccd1 vccd1
+ clock_div.count\[25\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_77_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_124_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3504__CLK clknet_leaf_31_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_187_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_176_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2829_ gamelogic.correct\[0\] gamelogic.rights\[0\] _0815_ vssd1 vssd1 vccd1 vccd1
+ _1367_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_135_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_96_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_122_Right_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3184__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2045__Y _0830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout50 _1395_ vssd1 vssd1 vccd1 vccd1 net50 sky130_fd_sc_hd__clkbuf_2
Xfanout61 net63 vssd1 vssd1 vccd1 vccd1 net61 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout83 net84 vssd1 vssd1 vccd1 vccd1 net83 sky130_fd_sc_hd__buf_2
XFILLER_0_36_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout72 net73 vssd1 vssd1 vccd1 vccd1 net72 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_153_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout94 _0824_ vssd1 vssd1 vccd1 vccd1 net94 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_36_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_112_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3527__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3620__X net38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_176_207 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2445__A2 host_message_reg.setLetter\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_0_clk_A clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_184_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1993_ net97 net93 vssd1 vssd1 vccd1 vccd1 _0826_ sky130_fd_sc_hd__nand2_1
XFILLER_0_129_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_71_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload20 clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 clkload20/Y sky130_fd_sc_hd__clkinv_1
XFILLER_0_125_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload31 clknet_leaf_19_clk vssd1 vssd1 vccd1 vccd1 clkload31/Y sky130_fd_sc_hd__inv_12
XFILLER_0_2_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2614_ net226 hostdisp.top\[69\] vssd1 vssd1 vccd1 vccd1 _1187_ sky130_fd_sc_hd__or2_1
XFILLER_0_100_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3594_ net157 vssd1 vssd1 vccd1 vccd1 net19 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_171_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2545_ hostdisp.bottom\[65\] dispFSM.guesses\[41\] net231 vssd1 vssd1 vccd1 vccd1
+ _1122_ sky130_fd_sc_hd__mux2_1
X_2476_ hostdisp.curr_word\[39\] net72 net69 net565 vssd1 vssd1 vccd1 vccd1 _0171_
+ sky130_fd_sc_hd__a22o_1
X_1427_ gamelogic.setWord\[36\] vssd1 vssd1 vccd1 vccd1 _0381_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout199_A net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3028_ clknet_leaf_8_clk clock_div.next_count\[8\] net214 vssd1 vssd1 vccd1 vccd1
+ clock_div.count\[8\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__2436__A2 host_message_reg.setLetter\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3599__264 vssd1 vssd1 vccd1 vccd1 net264 _3599__264/LO sky130_fd_sc_hd__conb_1
XFILLER_0_175_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_190_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload3 clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 clkload3/Y sky130_fd_sc_hd__clkinv_8
XFILLER_0_190_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_144_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2675__A2 net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout67_X net67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2427__A2 net70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_238 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_2_3__f_clk_X clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2330_ net74 _0982_ vssd1 vssd1 vccd1 vccd1 _0983_ sky130_fd_sc_hd__nor2_1
X_2261_ net307 buffer.temp_guess\[7\] net127 vssd1 vssd1 vccd1 vccd1 _0074_ sky130_fd_sc_hd__mux2_1
XANTENNA__1469__A3 net6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2192_ gamelogic.setWord\[30\] _0898_ net134 vssd1 vssd1 vccd1 vccd1 hostdisp.nextBottom\[78\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3229__RESET_B net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_190 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_210 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1976_ _0618_ _0810_ vssd1 vssd1 vccd1 vccd1 uart_receiver.temp_byte\[6\] sky130_fd_sc_hd__and2_1
XFILLER_0_15_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout114_A _1076_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3577_ net156 vssd1 vssd1 vccd1 vccd1 net9 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_60_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2528_ _1073_ _1093_ vssd1 vssd1 vccd1 vccd1 _1106_ sky130_fd_sc_hd__nor2_2
Xhold26 uart_transmitter.clk_count\[1\] vssd1 vssd1 vccd1 vccd1 net290 sky130_fd_sc_hd__dlygate4sd3_1
Xhold15 buffer.Rx_byte\[3\] vssd1 vssd1 vccd1 vccd1 net279 sky130_fd_sc_hd__dlygate4sd3_1
Xhold37 _0069_ vssd1 vssd1 vccd1 vccd1 net301 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2106__B2 gamelogic.letter\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2459_ net354 net71 _1052_ _0828_ vssd1 vssd1 vccd1 vccd1 _0158_ sky130_fd_sc_hd__a22o_1
Xhold59 uart_receiver.clk_count\[6\] vssd1 vssd1 vccd1 vccd1 net323 sky130_fd_sc_hd__dlygate4sd3_1
Xhold48 hostdisp.top\[73\] vssd1 vssd1 vccd1 vccd1 net312 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_148_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_22_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_49_Left_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_191_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3372__CLK clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_58_Left_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2648__A2 _1085_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_67_Left_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1830_ _0712_ vssd1 vssd1 vccd1 vccd1 _0713_ sky130_fd_sc_hd__inv_2
XANTENNA__2033__B1 net80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1761_ uart_transmitter.clk_count\[6\] uart_transmitter.clk_count\[7\] uart_transmitter.clk_count\[4\]
+ uart_transmitter.clk_count\[5\] vssd1 vssd1 vccd1 vccd1 _0663_ sky130_fd_sc_hd__or4_1
X_3500_ clknet_leaf_4_clk hostdisp.next_curr_word\[22\] net194 vssd1 vssd1 vccd1 vccd1
+ hostdisp.curr_word\[22\] sky130_fd_sc_hd__dfstp_1
X_1692_ _0010_ _0007_ vssd1 vssd1 vccd1 vccd1 keypadFSMHost.next_state\[1\] sky130_fd_sc_hd__or2_1
X_3431_ clknet_leaf_29_clk _0315_ vssd1 vssd1 vccd1 vccd1 lcdPlayer.nextState\[3\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_122_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3362_ clknet_leaf_23_clk _0251_ net182 vssd1 vssd1 vccd1 vccd1 dispFSM.guesses\[16\]
+ sky130_fd_sc_hd__dfstp_1
X_2313_ _0971_ vssd1 vssd1 vccd1 vccd1 _0972_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_76_Left_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3293_ clknet_leaf_35_clk _0214_ net162 vssd1 vssd1 vccd1 vccd1 gamelogic.rights\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_2244_ net155 net265 _0933_ vssd1 vssd1 vccd1 vccd1 _0045_ sky130_fd_sc_hd__mux2_1
XANTENNA__2639__A2 net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2175_ gamelogic.setWord\[30\] hostdisp.curr_guesses\[30\] net123 vssd1 vssd1 vccd1
+ vccd1 _0890_ sky130_fd_sc_hd__mux2_1
XFILLER_0_164_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_177_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3245__CLK clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_192_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_180_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout231_A net7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2024__B1 net79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1959_ uart_receiver.bit_index\[2\] net149 uart_receiver.bit_index\[0\] vssd1 vssd1
+ vccd1 vccd1 _0799_ sky130_fd_sc_hd__or3b_1
XANTENNA_fanout117_X net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput16 net16 vssd1 vssd1 vccd1 vccd1 gpio_oeb[19] sky130_fd_sc_hd__buf_2
Xoutput38 net38 vssd1 vssd1 vccd1 vccd1 gpio_out[28] sky130_fd_sc_hd__buf_2
Xoutput27 net27 vssd1 vssd1 vccd1 vccd1 gpio_oeb[8] sky130_fd_sc_hd__buf_2
XFILLER_0_3_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_183_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2015__B1 net80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_184 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3118__CLK clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3268__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_186_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_159_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2931_ net460 net89 net65 net444 vssd1 vssd1 vccd1 vccd1 _0298_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_33_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_0_clk clk vssd1 vssd1 vccd1 vccd1 clknet_0_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_84_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2862_ gamelogic.letter\[6\] buffer.temp_guess\[6\] _0918_ vssd1 vssd1 vccd1 vccd1
+ _1388_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_174 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2793_ net153 net151 _0560_ vssd1 vssd1 vccd1 vccd1 _1341_ sky130_fd_sc_hd__or3_1
X_1813_ clock_div.count\[7\] clock_div.count\[8\] _0700_ clock_div.count\[9\] vssd1
+ vssd1 vccd1 vccd1 _0702_ sky130_fd_sc_hd__a31o_1
XFILLER_0_127_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2006__B1 net77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1744_ _0641_ _0650_ _0651_ vssd1 vssd1 vccd1 vccd1 uart_receiver.next_clk_count\[5\]
+ sky130_fd_sc_hd__and3_1
Xhold304 hostdisp.curr_word\[21\] vssd1 vssd1 vccd1 vccd1 net568 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1675_ keypadHostt.scan_col\[0\] _0548_ _0556_ vssd1 vssd1 vccd1 vccd1 _0598_ sky130_fd_sc_hd__or3_1
XFILLER_0_159_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3414_ clknet_leaf_23_clk _0303_ net187 vssd1 vssd1 vccd1 vccd1 dispFSM.guesses\[68\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_110_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_15_Right_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3345_ clknet_leaf_33_clk _0234_ net164 vssd1 vssd1 vccd1 vccd1 gamelogic.letter\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_3276_ clknet_leaf_2_clk hostdisp.nextBottom\[74\] net170 vssd1 vssd1 vccd1 vccd1
+ hostdisp.bottom\[74\] sky130_fd_sc_hd__dfrtp_1
X_2227_ gamelogic.state\[3\] gamelogic.state\[2\] vssd1 vssd1 vccd1 vccd1 _0922_ sky130_fd_sc_hd__or2_1
XFILLER_0_108_70 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout181_A net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2158_ net552 _0881_ net136 vssd1 vssd1 vccd1 vccd1 hostdisp.nextBottom\[61\] sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_127_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_24_Right_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_311 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2089_ _0847_ _0849_ vssd1 vssd1 vccd1 vccd1 _0850_ sky130_fd_sc_hd__nand2_2
XFILLER_0_165_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_165_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_179_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2548__A1 net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_169_Right_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_33_Right_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout94_A _0824_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3410__CLK clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_42_Right_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_168_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_288 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_55_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_183_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_51_Right_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_156_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_136_Right_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1460_ hostdisp.curr_word\[39\] vssd1 vssd1 vccd1 vccd1 _0413_ sky130_fd_sc_hd__inv_2
XANTENNA__3090__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3130_ clknet_leaf_18_clk uart_transmitter.next_clk_count\[10\] net219 vssd1 vssd1
+ vccd1 vccd1 uart_transmitter.clk_count\[10\] sky130_fd_sc_hd__dfrtp_1
X_3061_ clknet_leaf_15_clk _0054_ _0023_ vssd1 vssd1 vccd1 vccd1 keypadFSMPlayer.prev_key\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_60_Right_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_166_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2012_ hostdisp.curr_guesses\[26\] net91 net76 net491 vssd1 vssd1 vccd1 vccd1 hostdisp.next_curr_guesses\[18\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_159_154 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2778__A1 host_message_reg.setLetter\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2914_ dispFSM.guesses\[54\] net85 net60 net508 vssd1 vssd1 vccd1 vccd1 _0281_ sky130_fd_sc_hd__o22a_1
XFILLER_0_57_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2845_ gamelogic.incorrect\[0\] gamelogic.incorrect\[1\] vssd1 vssd1 vccd1 vccd1
+ _1379_ sky130_fd_sc_hd__nand2_1
XFILLER_0_170_330 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold101 keypadFSMHost.prev_key\[3\] vssd1 vssd1 vccd1 vccd1 net365 sky130_fd_sc_hd__dlygate4sd3_1
X_2776_ _1325_ _1326_ vssd1 vssd1 vccd1 vccd1 _1328_ sky130_fd_sc_hd__nor2_1
XFILLER_0_53_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold134 keypadFSMHost.prev_key\[7\] vssd1 vssd1 vccd1 vccd1 net398 sky130_fd_sc_hd__dlygate4sd3_1
Xhold112 keypadFSMHost.prev_key\[2\] vssd1 vssd1 vccd1 vccd1 net376 sky130_fd_sc_hd__dlygate4sd3_1
Xhold123 keypadFSMHost.prev_key\[4\] vssd1 vssd1 vccd1 vccd1 net387 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_103_Right_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1727_ _0619_ net127 _0621_ vssd1 vssd1 vccd1 vccd1 _0640_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_79_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1658_ _0373_ _0490_ _0492_ vssd1 vssd1 vccd1 vccd1 _0588_ sky130_fd_sc_hd__nand3_1
Xhold145 hostdisp.curr_guesses\[13\] vssd1 vssd1 vccd1 vccd1 net409 sky130_fd_sc_hd__dlygate4sd3_1
Xhold167 hostdisp.curr_guesses\[37\] vssd1 vssd1 vccd1 vccd1 net431 sky130_fd_sc_hd__dlygate4sd3_1
Xhold156 hostdisp.curr_guesses\[0\] vssd1 vssd1 vccd1 vccd1 net420 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_186_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold178 uart_transmitter.clk_count\[10\] vssd1 vssd1 vccd1 vccd1 net442 sky130_fd_sc_hd__dlygate4sd3_1
Xhold189 dispFSM.guesses\[61\] vssd1 vssd1 vccd1 vccd1 net453 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_186_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1589_ _0437_ _0532_ _0448_ vssd1 vssd1 vccd1 vccd1 _0533_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_129_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3328_ clknet_leaf_35_clk gamelogic.nextState\[2\] net162 vssd1 vssd1 vccd1 vccd1
+ gamelogic.state\[2\] sky130_fd_sc_hd__dfrtp_4
X_3259_ clknet_leaf_5_clk hostdisp.nextBottom\[57\] net197 vssd1 vssd1 vccd1 vccd1
+ hostdisp.bottom\[57\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout184_X net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2769__A1 host_message_reg.setLetter\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2044__B _0822_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_352 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2941__A1 dispFSM.msg\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout97_X net97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_147_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3306__CLK clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_269 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_280 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2630_ net283 net107 _1202_ net188 vssd1 vssd1 vccd1 vccd1 _0179_ sky130_fd_sc_hd__o211a_1
XANTENNA__3456__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2561_ _1134_ _1135_ _1136_ net226 vssd1 vssd1 vccd1 vccd1 _1137_ sky130_fd_sc_hd__o31a_1
XFILLER_0_50_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1512_ _0460_ _0461_ vssd1 vssd1 vccd1 vccd1 _0462_ sky130_fd_sc_hd__and2_1
X_2492_ net138 _0356_ vssd1 vssd1 vccd1 vccd1 _1070_ sky130_fd_sc_hd__nand2_4
X_1443_ uart_transmitter.state\[2\] vssd1 vssd1 vccd1 vccd1 _0397_ sky130_fd_sc_hd__inv_2
XFILLER_0_120_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3113_ clknet_leaf_28_clk _0103_ vssd1 vssd1 vccd1 vccd1 lcdPlayer.cnt_500hz\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_179_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3044_ clknet_leaf_7_clk clock_div.next_count\[24\] net195 vssd1 vssd1 vccd1 vccd1
+ clock_div.count\[24\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_65_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2129__B net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout144_A gamelogic.letter\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_176_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_12_Left_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2828_ _0815_ _0818_ _1365_ vssd1 vssd1 vccd1 vccd1 _1366_ sky130_fd_sc_hd__a21o_1
X_2759_ _0612_ _1293_ _1307_ vssd1 vssd1 vccd1 vccd1 _1312_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_135_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1990__Y _0823_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_21_Left_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3329__CLK clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_142_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_30_Left_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_153_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout62 net63 vssd1 vssd1 vccd1 vccd1 net62 sky130_fd_sc_hd__buf_2
XANTENNA__2206__A3 net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout51 net52 vssd1 vssd1 vccd1 vccd1 net51 sky130_fd_sc_hd__clkbuf_4
Xfanout73 _1030_ vssd1 vssd1 vccd1 vccd1 net73 sky130_fd_sc_hd__buf_2
XFILLER_0_153_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout84 _0940_ vssd1 vssd1 vccd1 vccd1 net84 sky130_fd_sc_hd__buf_2
Xfanout95 _0823_ vssd1 vssd1 vccd1 vccd1 net95 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_36_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_output38_A net38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_176_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_63_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2850__A0 net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1992_ net104 _0823_ vssd1 vssd1 vccd1 vccd1 _0825_ sky130_fd_sc_hd__nor2_1
XFILLER_0_129_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkload10 clknet_leaf_34_clk vssd1 vssd1 vccd1 vccd1 clkload10/Y sky130_fd_sc_hd__inv_12
XFILLER_0_42_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkload21 clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 clkload21/Y sky130_fd_sc_hd__inv_8
XFILLER_0_152_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkload32 clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 clkload32/X sky130_fd_sc_hd__clkbuf_8
X_2613_ hostdisp.bottom\[61\] dispFSM.guesses\[37\] net227 vssd1 vssd1 vccd1 vccd1
+ _1186_ sky130_fd_sc_hd__mux2_1
XANTENNA__2412__B net92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3593_ net156 vssd1 vssd1 vccd1 vccd1 net18 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2544_ _1117_ _1119_ _1120_ net227 vssd1 vssd1 vccd1 vccd1 _1121_ sky130_fd_sc_hd__o31a_1
XFILLER_0_23_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_171_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2118__C1 net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2475_ hostdisp.curr_word\[38\] net75 net68 net525 _1034_ vssd1 vssd1 vccd1 vccd1
+ _0170_ sky130_fd_sc_hd__a221o_1
X_1426_ gamelogic.letter\[3\] vssd1 vssd1 vccd1 vccd1 _0380_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_3_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_182_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3027_ clknet_leaf_8_clk clock_div.next_count\[7\] net213 vssd1 vssd1 vccd1 vccd1
+ clock_div.count\[7\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_190_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkload4 clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 clkload4/Y sky130_fd_sc_hd__inv_12
XFILLER_0_18_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_250 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout230 net231 vssd1 vssd1 vccd1 vccd1 net230 sky130_fd_sc_hd__clkbuf_2
XANTENNA__2124__A2 net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_144_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_17_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2260_ net305 buffer.temp_guess\[6\] net127 vssd1 vssd1 vccd1 vccd1 _0073_ sky130_fd_sc_hd__mux2_1
XANTENNA__1469__A4 net3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2191_ gamelogic.setWord\[38\] hostdisp.curr_guesses\[38\] net123 vssd1 vssd1 vccd1
+ vccd1 _0898_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_162_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_66 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_222 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1975_ buffer.Rx_byte\[6\] net2 _0809_ vssd1 vssd1 vccd1 vccd1 _0810_ sky130_fd_sc_hd__mux2_1
XFILLER_0_172_266 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_174 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3174__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3576_ net157 vssd1 vssd1 vccd1 vccd1 net28 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout107_A _0759_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2527_ _1089_ _1092_ _1104_ vssd1 vssd1 vccd1 vccd1 _1105_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_93_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2458_ hostdisp.curr_word\[26\] net119 vssd1 vssd1 vccd1 vccd1 _1052_ sky130_fd_sc_hd__or2_1
X_1409_ net151 vssd1 vssd1 vccd1 vccd1 _0363_ sky130_fd_sc_hd__inv_2
Xhold27 uart_transmitter.next_clk_count\[1\] vssd1 vssd1 vccd1 vccd1 net291 sky130_fd_sc_hd__dlygate4sd3_1
Xhold38 message_reg.msg\[2\] vssd1 vssd1 vccd1 vccd1 net302 sky130_fd_sc_hd__dlygate4sd3_1
Xhold16 _0070_ vssd1 vssd1 vccd1 vccd1 net280 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_89_Right_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2389_ lcdPlayer.cnt_20ms\[16\] lcdPlayer.cnt_20ms\[15\] _1014_ vssd1 vssd1 vccd1
+ vccd1 _1018_ sky130_fd_sc_hd__and3_1
Xhold49 hostdisp.top\[77\] vssd1 vssd1 vccd1 vccd1 net313 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2511__C1 _0360_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_98_Right_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_163_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_22_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_191_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2593__A2 _1078_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3517__CLK clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_5_Left_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3047__CLK clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1760_ _0397_ uart_transmitter.state\[1\] vssd1 vssd1 vccd1 vccd1 _0662_ sky130_fd_sc_hd__nand2_1
XFILLER_0_52_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3197__CLK clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1691_ keypadFSMHost.state\[2\] _0565_ _0606_ keypadFSMHost.state\[3\] vssd1 vssd1
+ vccd1 vccd1 _0007_ sky130_fd_sc_hd__a22o_1
XFILLER_0_122_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3430_ clknet_leaf_29_clk _0004_ vssd1 vssd1 vccd1 vccd1 lcdPlayer.nextState\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_3361_ clknet_leaf_21_clk _0250_ net204 vssd1 vssd1 vccd1 vccd1 dispFSM.guesses\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_2312_ lcdPlayer.cnt_500hz\[8\] lcdPlayer.cnt_500hz\[9\] lcdPlayer.cnt_500hz\[10\]
+ _0965_ vssd1 vssd1 vccd1 vccd1 _0971_ sky130_fd_sc_hd__and4_1
XFILLER_0_57_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3292_ clknet_leaf_35_clk _0213_ net162 vssd1 vssd1 vccd1 vccd1 gamelogic.rights\[0\]
+ sky130_fd_sc_hd__dfrtp_2
X_2243_ net155 _0933_ vssd1 vssd1 vccd1 vccd1 _0934_ sky130_fd_sc_hd__or2_2
X_2174_ gamelogic.setWord\[21\] _0889_ net137 vssd1 vssd1 vccd1 vccd1 hostdisp.nextBottom\[69\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2272__A1 dispFSM.msg\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_192_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_185_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2811__A3 _1286_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_288 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout224_A net225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1958_ _0618_ _0798_ vssd1 vssd1 vccd1 vccd1 uart_receiver.temp_byte\[0\] sky130_fd_sc_hd__and2_1
XANTENNA__2575__A2 net105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1889_ uart_transmitter.clk_count\[6\] uart_transmitter.clk_count\[7\] _0740_ uart_transmitter.clk_count\[8\]
+ vssd1 vssd1 vccd1 vccd1 _0745_ sky130_fd_sc_hd__a31o_1
XANTENNA__1992__A net104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput39 net39 vssd1 vssd1 vccd1 vccd1 gpio_out[29] sky130_fd_sc_hd__buf_2
XFILLER_0_113_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput17 net17 vssd1 vssd1 vccd1 vccd1 gpio_oeb[25] sky130_fd_sc_hd__buf_2
Xoutput28 net28 vssd1 vssd1 vccd1 vccd1 gpio_oeb[9] sky130_fd_sc_hd__buf_2
X_3559_ clknet_leaf_7_clk hostdisp.next_curr_guesses\[41\] net196 vssd1 vssd1 vccd1
+ vccd1 hostdisp.curr_guesses\[41\] sky130_fd_sc_hd__dfstp_1
XFILLER_0_11_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_183_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_117_Right_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_151_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2998__A net221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2566__A2 net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkload2_A clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_186_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2930_ dispFSM.guesses\[70\] net85 net61 net485 vssd1 vssd1 vccd1 vccd1 _0297_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_33_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_79 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1796__B _0693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2861_ net66 _1387_ vssd1 vssd1 vccd1 vccd1 _0232_ sky130_fd_sc_hd__and2_1
XFILLER_0_84_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1812_ net372 _0701_ vssd1 vssd1 vccd1 vccd1 clock_div.next_count\[8\] sky130_fd_sc_hd__xnor2_1
X_2792_ _0560_ _1339_ vssd1 vssd1 vccd1 vccd1 _1340_ sky130_fd_sc_hd__nand2_1
XFILLER_0_111_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1743_ uart_receiver.clk_count\[4\] _0646_ uart_receiver.clk_count\[5\] vssd1 vssd1
+ vccd1 vccd1 _0651_ sky130_fd_sc_hd__a21o_1
XANTENNA__2557__A2 net114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1674_ _0596_ vssd1 vssd1 vccd1 vccd1 _0597_ sky130_fd_sc_hd__inv_2
Xhold305 gamelogic.setWord\[13\] vssd1 vssd1 vccd1 vccd1 net569 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3413_ clknet_leaf_23_clk _0302_ net184 vssd1 vssd1 vccd1 vccd1 dispFSM.guesses\[67\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_68_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2190__A0 gamelogic.setWord\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3344_ clknet_leaf_33_clk _0233_ net163 vssd1 vssd1 vccd1 vccd1 gamelogic.letter\[6\]
+ sky130_fd_sc_hd__dfrtp_4
X_3275_ clknet_leaf_14_clk hostdisp.nextBottom\[73\] net199 vssd1 vssd1 vccd1 vccd1
+ hostdisp.bottom\[73\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_175_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2226_ _0364_ _0916_ vssd1 vssd1 vccd1 vccd1 _0921_ sky130_fd_sc_hd__nor2_1
XFILLER_0_177_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2157_ gamelogic.setWord\[21\] hostdisp.curr_guesses\[21\] net125 vssd1 vssd1 vccd1
+ vccd1 _0881_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout174_A net180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3362__CLK clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2088_ hostdisp.curr_word\[24\] net101 net75 _0848_ gamelogic.indexCorrect\[3\] vssd1
+ vssd1 vccd1 vccd1 _0849_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_48_323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_179_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_180_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2650__D1 net226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1993__Y _0826_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout227_X net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_99_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1926__S _0764_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout87_A _0940_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_95_Left_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_183_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_171_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_30_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2539__A2 _1072_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3060_ clknet_leaf_12_clk _0053_ _0022_ vssd1 vssd1 vccd1 vccd1 keypadFSMPlayer.prev_key\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_2011_ hostdisp.curr_guesses\[25\] net93 net79 net487 vssd1 vssd1 vccd1 vccd1 hostdisp.next_curr_guesses\[17\]
+ sky130_fd_sc_hd__o22a_1
XANTENNA__3385__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_234 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2913_ net388 net90 net64 net373 vssd1 vssd1 vccd1 vccd1 _0280_ sky130_fd_sc_hd__a22o_1
XFILLER_0_45_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2844_ _0821_ _1378_ gamelogic.incorrect\[0\] vssd1 vssd1 vccd1 vccd1 _0224_ sky130_fd_sc_hd__mux2_1
XFILLER_0_170_342 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2775_ _1325_ _1326_ vssd1 vssd1 vccd1 vccd1 _1327_ sky130_fd_sc_hd__and2_1
XFILLER_0_13_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold113 keypadFSMPlayer.prev_key\[2\] vssd1 vssd1 vccd1 vccd1 net377 sky130_fd_sc_hd__dlygate4sd3_1
Xhold102 keypadFSMHost.prev_key\[5\] vssd1 vssd1 vccd1 vccd1 net366 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_239 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold124 dispFSM.guesses\[53\] vssd1 vssd1 vccd1 vccd1 net388 sky130_fd_sc_hd__dlygate4sd3_1
X_1726_ _0618_ _0621_ _0623_ _0631_ vssd1 vssd1 vccd1 vccd1 uart_receiver.next_state\[2\]
+ sky130_fd_sc_hd__a31o_1
Xhold135 lcdPlayer.cnt_20ms\[12\] vssd1 vssd1 vccd1 vccd1 net399 sky130_fd_sc_hd__dlygate4sd3_1
X_1657_ _0016_ _0013_ vssd1 vssd1 vccd1 vccd1 keypadFSMPlayer.next_state\[1\] sky130_fd_sc_hd__or2_1
XFILLER_0_110_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold168 dispFSM.guesses\[4\] vssd1 vssd1 vccd1 vccd1 net432 sky130_fd_sc_hd__dlygate4sd3_1
Xhold157 hostdisp.curr_word\[29\] vssd1 vssd1 vccd1 vccd1 net421 sky130_fd_sc_hd__dlygate4sd3_1
Xhold146 hostdisp.curr_guesses\[2\] vssd1 vssd1 vccd1 vccd1 net410 sky130_fd_sc_hd__dlygate4sd3_1
X_1588_ _0508_ _0531_ vssd1 vssd1 vccd1 vccd1 _0532_ sky130_fd_sc_hd__xnor2_1
Xhold179 lcdPlayer.cnt_20ms\[8\] vssd1 vssd1 vccd1 vccd1 net443 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_186_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2702__A2 gamelogic.setWord\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3327_ clknet_leaf_35_clk gamelogic.nextState\[1\] net162 vssd1 vssd1 vccd1 vccd1
+ gamelogic.state\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_95_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_185_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3258_ clknet_leaf_5_clk hostdisp.nextBottom\[56\] net193 vssd1 vssd1 vccd1 vccd1
+ hostdisp.bottom\[56\] sky130_fd_sc_hd__dfrtp_1
X_2209_ net129 gamelogic.setWord\[39\] vssd1 vssd1 vccd1 vccd1 _0907_ sky130_fd_sc_hd__and2_1
XANTENNA__2466__B2 _0828_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3189_ clknet_leaf_29_clk _0165_ net166 vssd1 vssd1 vccd1 vccd1 hostdisp.top\[73\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_180_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_394 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold301_A hostdisp.top\[79\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_364 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3258__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_147_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2457__B2 _0828_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_43_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_2_0__f_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_2_0__leaf_clk sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_158_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_147 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_117_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2560_ dispFSM.guesses\[42\] net111 net109 dispFSM.guesses\[34\] _1133_ vssd1 vssd1
+ vccd1 vccd1 _1136_ sky130_fd_sc_hd__a221o_1
X_1511_ net148 net155 vssd1 vssd1 vccd1 vccd1 _0461_ sky130_fd_sc_hd__nand2_1
X_2491_ net138 _0356_ vssd1 vssd1 vccd1 vccd1 _1069_ sky130_fd_sc_hd__and2_1
X_1442_ uart_receiver.state\[0\] vssd1 vssd1 vccd1 vccd1 _0396_ sky130_fd_sc_hd__inv_2
X_3112_ clknet_leaf_28_clk _0102_ vssd1 vssd1 vccd1 vccd1 lcdPlayer.cnt_500hz\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_65_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_179_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3043_ clknet_leaf_7_clk clock_div.next_count\[23\] net195 vssd1 vssd1 vccd1 vccd1
+ clock_div.count\[23\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_66_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_124_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout137_A hostdisp.Cstate vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2827_ _0910_ _0911_ _0925_ _0927_ vssd1 vssd1 vccd1 vccd1 _1365_ sky130_fd_sc_hd__or4_1
XFILLER_0_83_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2758_ _1311_ _1309_ _1290_ host_message_reg.setLetter\[0\] vssd1 vssd1 vccd1 vccd1
+ _0205_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_135_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1709_ _0538_ _0596_ vssd1 vssd1 vccd1 vccd1 _0625_ sky130_fd_sc_hd__nor2_1
XANTENNA__3550__CLK clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2689_ net142 gamelogic.setWord\[28\] vssd1 vssd1 vccd1 vccd1 _1254_ sky130_fd_sc_hd__xnor2_1
XANTENNA__2687__A1 net144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_169_Left_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_193_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout63 _1391_ vssd1 vssd1 vccd1 vccd1 net63 sky130_fd_sc_hd__clkbuf_2
Xfanout52 _1393_ vssd1 vssd1 vccd1 vccd1 net52 sky130_fd_sc_hd__buf_2
XANTENNA__3080__CLK clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout74 _0957_ vssd1 vssd1 vccd1 vccd1 net74 sky130_fd_sc_hd__buf_2
XFILLER_0_76_292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout85 net87 vssd1 vssd1 vccd1 vccd1 net85 sky130_fd_sc_hd__buf_2
XFILLER_0_24_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout96 _0626_ vssd1 vssd1 vccd1 vccd1 net96 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_36_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_178_Left_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_187_Left_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2517__Y _1095_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3423__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_71_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1991_ net131 _0821_ vssd1 vssd1 vccd1 vccd1 _0824_ sky130_fd_sc_hd__nand2_1
XFILLER_0_144_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2602__A1 _0360_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkload22 clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 clkload22/Y sky130_fd_sc_hd__inv_8
XFILLER_0_140_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkload33 clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 clkload33/X sky130_fd_sc_hd__clkbuf_4
X_2612_ hostdisp.bottom\[45\] _1081_ _1184_ net227 vssd1 vssd1 vccd1 vccd1 _1185_
+ sky130_fd_sc_hd__a211o_1
X_3592_ net157 vssd1 vssd1 vccd1 vccd1 net17 sky130_fd_sc_hd__clkbuf_1
Xclkload11 clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 clkload11/Y sky130_fd_sc_hd__inv_6
X_2543_ dispFSM.guesses\[25\] net114 _1084_ dispFSM.guesses\[1\] vssd1 vssd1 vccd1
+ vccd1 _1120_ sky130_fd_sc_hd__a22o_1
XFILLER_0_23_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_171_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2474_ net313 net68 _1056_ vssd1 vssd1 vccd1 vccd1 _0169_ sky130_fd_sc_hd__a21bo_1
X_1425_ gamelogic.letter\[2\] vssd1 vssd1 vccd1 vccd1 _0379_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_183_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_182_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3026_ clknet_leaf_8_clk clock_div.next_count\[6\] net217 vssd1 vssd1 vccd1 vccd1
+ clock_div.count\[6\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_65_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkload5 clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 clkload5/Y sky130_fd_sc_hd__clkinv_8
XFILLER_0_18_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout220 net221 vssd1 vssd1 vccd1 vccd1 net220 sky130_fd_sc_hd__buf_2
Xfanout231 net7 vssd1 vssd1 vccd1 vccd1 net231 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_144_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3446__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2734__C_N keypadFSMHost.state\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2190_ gamelogic.setWord\[29\] _0897_ net137 vssd1 vssd1 vccd1 vccd1 hostdisp.nextBottom\[77\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2263__X _0940_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1974_ net150 net149 uart_receiver.bit_index\[2\] vssd1 vssd1 vccd1 vccd1 _0809_
+ sky130_fd_sc_hd__and3b_1
XANTENNA__2051__A2 net96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3575_ net156 vssd1 vssd1 vccd1 vccd1 net27 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_178_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_140_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2526_ _1100_ _1101_ _1103_ vssd1 vssd1 vccd1 vccd1 _1104_ sky130_fd_sc_hd__or3_2
XANTENNA__3469__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2457_ net331 net70 _1051_ _0828_ vssd1 vssd1 vccd1 vccd1 _0157_ sky130_fd_sc_hd__a22o_1
X_1408_ keypadHostt.scan_col\[3\] vssd1 vssd1 vccd1 vccd1 _0362_ sky130_fd_sc_hd__inv_2
Xhold17 message_reg.msg\[4\] vssd1 vssd1 vccd1 vccd1 net281 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_46_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold28 net43 vssd1 vssd1 vccd1 vccd1 net292 sky130_fd_sc_hd__dlygate4sd3_1
Xhold39 buffer.Rx_byte\[4\] vssd1 vssd1 vccd1 vccd1 net303 sky130_fd_sc_hd__dlygate4sd3_1
X_2388_ _1017_ net182 _1016_ vssd1 vssd1 vccd1 vccd1 _0122_ sky130_fd_sc_hd__and3b_1
XFILLER_0_127_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3009_ net211 vssd1 vssd1 vccd1 vccd1 _0034_ sky130_fd_sc_hd__inv_2
XFILLER_0_78_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2614__A net226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2578__B1 net226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_191_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_150_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2033__A2 net95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2569__B1 _1095_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1690_ keypadFSMHost.state\[5\] _0565_ _0606_ keypadFSMHost.state\[2\] vssd1 vssd1
+ vccd1 vccd1 _0010_ sky130_fd_sc_hd__a22o_1
XFILLER_0_52_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3360_ clknet_leaf_20_clk _0249_ net204 vssd1 vssd1 vccd1 vccd1 dispFSM.guesses\[14\]
+ sky130_fd_sc_hd__dfstp_1
X_2311_ net493 _0967_ _0970_ vssd1 vssd1 vccd1 vccd1 _0092_ sky130_fd_sc_hd__o21a_1
X_3291_ clknet_leaf_13_clk host_message_reg.next_state net197 vssd1 vssd1 vccd1 vccd1
+ host_message_reg.Cstate sky130_fd_sc_hd__dfrtp_4
XFILLER_0_20_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2242_ _0360_ _0693_ vssd1 vssd1 vccd1 vccd1 _0933_ sky130_fd_sc_hd__or2_1
X_2173_ gamelogic.setWord\[29\] hostdisp.curr_guesses\[29\] net125 vssd1 vssd1 vccd1
+ vccd1 _0889_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3546__SET_B net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2024__A2 net94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1957_ net2 buffer.Rx_byte\[0\] _0797_ vssd1 vssd1 vccd1 vccd1 _0798_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout217_A net218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1888_ net353 _0742_ _0744_ vssd1 vssd1 vccd1 vccd1 uart_transmitter.next_clk_count\[7\]
+ sky130_fd_sc_hd__a21oi_1
XANTENNA__1992__B _0823_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3558_ clknet_leaf_6_clk hostdisp.next_curr_guesses\[40\] net191 vssd1 vssd1 vccd1
+ vccd1 hostdisp.curr_guesses\[40\] sky130_fd_sc_hd__dfstp_1
Xoutput29 net29 vssd1 vssd1 vccd1 vccd1 gpio_out[10] sky130_fd_sc_hd__buf_2
XFILLER_0_101_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput18 net18 vssd1 vssd1 vccd1 vccd1 gpio_oeb[26] sky130_fd_sc_hd__buf_2
XFILLER_0_3_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2509_ _1060_ _1074_ vssd1 vssd1 vccd1 vccd1 _1087_ sky130_fd_sc_hd__nor2_1
X_3489_ clknet_leaf_30_clk hostdisp.next_curr_word\[11\] net174 vssd1 vssd1 vccd1
+ vccd1 hostdisp.curr_word\[11\] sky130_fd_sc_hd__dfstp_1
XFILLER_0_78_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2015__A2 net95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1423__A net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1710__X _0626_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_27_clk clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_27_clk
+ sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_114_Left_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3164__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2860_ net141 buffer.temp_guess\[5\] _0918_ vssd1 vssd1 vccd1 vccd1 _1387_ sky130_fd_sc_hd__mux2_1
X_1811_ _0687_ _0692_ _0700_ clock_div.count\[7\] _0701_ vssd1 vssd1 vccd1 vccd1 clock_div.next_count\[7\]
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_72_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2791_ _0540_ _0543_ _0551_ vssd1 vssd1 vccd1 vccd1 _1339_ sky130_fd_sc_hd__o21ai_1
XANTENNA__2006__A2 net92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1742_ _0649_ vssd1 vssd1 vccd1 vccd1 _0650_ sky130_fd_sc_hd__inv_2
X_1673_ _0549_ _0584_ vssd1 vssd1 vccd1 vccd1 _0596_ sky130_fd_sc_hd__nand2_1
XANTENNA__2962__B1 net50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_150_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_112 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3412_ clknet_leaf_24_clk _0301_ net189 vssd1 vssd1 vccd1 vccd1 dispFSM.guesses\[66\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_7_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_68 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_123_Left_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3343_ clknet_leaf_33_clk _0232_ net163 vssd1 vssd1 vccd1 vccd1 gamelogic.letter\[5\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_68_88 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3274_ clknet_leaf_5_clk hostdisp.nextBottom\[72\] net191 vssd1 vssd1 vccd1 vccd1
+ hostdisp.bottom\[72\] sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_183_Right_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2225_ _0910_ _0919_ _0815_ vssd1 vssd1 vccd1 vccd1 _0920_ sky130_fd_sc_hd__a21o_1
X_2156_ gamelogic.setWord\[12\] _0880_ net132 vssd1 vssd1 vccd1 vccd1 hostdisp.nextBottom\[60\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3507__CLK clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_18_clk clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_18_clk
+ sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_132_Left_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_127_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_5_Right_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout167_A net169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2087_ hostdisp.curr_word\[26\] hostdisp.curr_word\[28\] _0411_ net101 vssd1 vssd1
+ vccd1 vccd1 _0848_ sky130_fd_sc_hd__a31o_1
XFILLER_0_177_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_335 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_179_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2989_ gamelogic.setWord\[28\] net52 net48 gamelogic.setWord\[36\] vssd1 vssd1 vccd1
+ vccd1 _0352_ sky130_fd_sc_hd__o22a_1
XFILLER_0_16_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout122_X net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_141_Left_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_140_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2953__B1 net50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_150_Right_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3187__CLK clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_150_Left_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3231__Q host_message_reg.setLetter\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_183_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_191_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2802__A net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_145_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2010_ hostdisp.curr_guesses\[24\] net93 net78 net538 vssd1 vssd1 vccd1 vccd1 hostdisp.next_curr_guesses\[16\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_159_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2475__A2 net75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_246 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2912_ dispFSM.guesses\[52\] net83 net58 net505 vssd1 vssd1 vccd1 vccd1 _0279_ sky130_fd_sc_hd__o22a_1
XFILLER_0_45_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2843_ _0815_ _0820_ _1365_ vssd1 vssd1 vccd1 vccd1 _1378_ sky130_fd_sc_hd__a21o_1
X_2774_ _1316_ _1319_ _1300_ vssd1 vssd1 vccd1 vccd1 _1326_ sky130_fd_sc_hd__o21a_1
XFILLER_0_170_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1725_ _0633_ _0637_ _0639_ _0624_ vssd1 vssd1 vccd1 vccd1 uart_receiver.next_state\[1\]
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_53_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold103 keypadFSMPlayer.prev_key\[1\] vssd1 vssd1 vccd1 vccd1 net367 sky130_fd_sc_hd__dlygate4sd3_1
Xhold114 keypadFSMPlayer.prev_key\[7\] vssd1 vssd1 vccd1 vccd1 net378 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold125 _0288_ vssd1 vssd1 vccd1 vccd1 net389 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1656_ keypadFSMPlayer.state\[2\] _0452_ _0587_ keypadFSMPlayer.state\[3\] vssd1
+ vssd1 vccd1 vccd1 _0013_ sky130_fd_sc_hd__a22o_1
Xhold147 clock_div.count\[20\] vssd1 vssd1 vccd1 vccd1 net411 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_7_clk clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_7_clk
+ sky130_fd_sc_hd__clkbuf_8
Xhold136 hostdisp.curr_guesses\[21\] vssd1 vssd1 vccd1 vccd1 net400 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold158 lcdPlayer.cnt_20ms\[10\] vssd1 vssd1 vccd1 vccd1 net422 sky130_fd_sc_hd__dlygate4sd3_1
X_1587_ _0495_ _0499_ _0490_ vssd1 vssd1 vccd1 vccd1 _0531_ sky130_fd_sc_hd__or3b_1
Xhold169 hostdisp.curr_guesses\[31\] vssd1 vssd1 vccd1 vccd1 net433 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_186_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3326_ clknet_leaf_33_clk gamelogic.nextState\[0\] net162 vssd1 vssd1 vccd1 vccd1
+ gamelogic.state\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_95_64 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3257_ clknet_leaf_22_clk hostdisp.nextBottom\[55\] net186 vssd1 vssd1 vccd1 vccd1
+ hostdisp.bottom\[55\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_69_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_185_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2208_ net134 hostdisp.curr_guesses\[46\] net123 _0906_ vssd1 vssd1 vccd1 vccd1 hostdisp.nextBottom\[86\]
+ sky130_fd_sc_hd__a31o_1
XANTENNA__2466__A2 net70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3188_ clknet_leaf_31_clk _0164_ net172 vssd1 vssd1 vccd1 vccd1 hostdisp.top\[72\]
+ sky130_fd_sc_hd__dfrtp_1
X_2139_ gamelogic.setWord\[12\] hostdisp.curr_guesses\[12\] net123 vssd1 vssd1 vccd1
+ vccd1 _0872_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_318 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_290 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1977__A1 net2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_161_376 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_147_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2457__A2 net70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_158_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3202__CLK clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_152_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1510_ net147 net155 vssd1 vssd1 vccd1 vccd1 _0460_ sky130_fd_sc_hd__nand2_1
XFILLER_0_105_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2490_ lcdPlayer.nextState\[3\] lcdPlayer.nextState\[2\] vssd1 vssd1 vccd1 vccd1
+ _1068_ sky130_fd_sc_hd__nor2_1
X_1441_ keypadFSMHost.state\[4\] vssd1 vssd1 vccd1 vccd1 _0395_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3111_ clknet_leaf_28_clk _0101_ vssd1 vssd1 vccd1 vccd1 lcdPlayer.cnt_500hz\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_65_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3042_ clknet_leaf_8_clk clock_div.next_count\[22\] net213 vssd1 vssd1 vccd1 vccd1
+ clock_div.count\[22\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__2448__A2 net71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3601__235 vssd1 vssd1 vccd1 vccd1 _3601__235/HI net235 sky130_fd_sc_hd__conb_1
XANTENNA__2707__A net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_147_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_124_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2426__B net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_99 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_155_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2826_ gamelogic.indexCorrect\[1\] _1364_ _1236_ vssd1 vssd1 vccd1 vccd1 _0220_ sky130_fd_sc_hd__o21a_1
XFILLER_0_143_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2757_ host_message_reg.setLetter\[0\] _0601_ _1310_ vssd1 vssd1 vccd1 vccd1 _1311_
+ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_135_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2688_ _0378_ gamelogic.setWord\[25\] gamelogic.setWord\[29\] _0384_ _1250_ vssd1
+ vssd1 vccd1 vccd1 _1253_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_96_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1708_ _0621_ _0623_ _0619_ vssd1 vssd1 vccd1 vccd1 _0624_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_41_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1639_ _0368_ _0543_ _0552_ vssd1 vssd1 vccd1 vccd1 _0574_ sky130_fd_sc_hd__and3_1
XFILLER_0_111_262 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input4_A gpio_in[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3309_ clknet_leaf_34_clk uart_receiver.next_clk_count\[1\] net158 vssd1 vssd1 vccd1
+ vccd1 uart_receiver.clk_count\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_68_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout53 _1393_ vssd1 vssd1 vccd1 vccd1 net53 sky130_fd_sc_hd__clkbuf_4
Xfanout64 _1390_ vssd1 vssd1 vccd1 vccd1 net64 sky130_fd_sc_hd__buf_2
XFILLER_0_36_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout97 _0626_ vssd1 vssd1 vccd1 vccd1 net97 sky130_fd_sc_hd__buf_2
Xfanout86 net87 vssd1 vssd1 vccd1 vccd1 net86 sky130_fd_sc_hd__buf_2
XFILLER_0_134_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2611__A2 net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout75 _0830_ vssd1 vssd1 vccd1 vccd1 net75 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_134_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3375__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_284 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1431__A gamelogic.letter\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2246__B _0693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1990_ net129 _0822_ vssd1 vssd1 vccd1 vccd1 _0823_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_28_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkload23 clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 clkload23/Y sky130_fd_sc_hd__clkinv_4
X_2611_ hostdisp.bottom\[53\] net115 _1182_ _1183_ vssd1 vssd1 vccd1 vccd1 _1184_
+ sky130_fd_sc_hd__a211o_1
Xclkload34 clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 clkload34/Y sky130_fd_sc_hd__inv_4
XTAP_TAPCELL_ROW_11_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3591_ net263 vssd1 vssd1 vccd1 vccd1 gpio_oeb[24] sky130_fd_sc_hd__buf_2
Xclkload12 clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 clkload12/Y sky130_fd_sc_hd__inv_6
X_2542_ dispFSM.guesses\[17\] _1081_ net108 dispFSM.msg\[1\] _1118_ vssd1 vssd1 vccd1
+ vccd1 _1119_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_171_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_167_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2473_ _0412_ net75 net68 _1034_ vssd1 vssd1 vccd1 vccd1 _1056_ sky130_fd_sc_hd__a211o_1
XFILLER_0_167_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1424_ net144 vssd1 vssd1 vccd1 vccd1 _0378_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_3_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3026__RESET_B net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3025_ clknet_leaf_9_clk clock_div.next_count\[5\] net217 vssd1 vssd1 vccd1 vccd1
+ clock_div.count\[5\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__3248__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_182_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3398__CLK clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_118 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkload6 clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 clkload6/Y sky130_fd_sc_hd__clkinv_8
XFILLER_0_143_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2809_ _1347_ _1353_ _1354_ vssd1 vssd1 vccd1 vccd1 _1355_ sky130_fd_sc_hd__and3_1
XFILLER_0_33_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout202_X net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2109__B2 net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout232 net233 vssd1 vssd1 vccd1 vccd1 net232 sky130_fd_sc_hd__buf_2
Xfanout221 net224 vssd1 vssd1 vccd1 vccd1 net221 sky130_fd_sc_hd__buf_4
Xfanout210 net212 vssd1 vssd1 vccd1 vccd1 net210 sky130_fd_sc_hd__clkbuf_4
XANTENNA_input7_X net7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_144_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_103_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_25_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1426__A gamelogic.letter\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2809__X _1355_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2528__Y _1106_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3540__CLK clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1973_ _0618_ _0808_ vssd1 vssd1 vccd1 vccd1 uart_receiver.temp_byte\[5\] sky130_fd_sc_hd__and2_1
XFILLER_0_15_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_140_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_132_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3574_ net156 vssd1 vssd1 vccd1 vccd1 net26 sky130_fd_sc_hd__clkbuf_1
X_2525_ hostdisp.top\[64\] _1096_ _1097_ hostdisp.top\[48\] _1102_ vssd1 vssd1 vccd1
+ vccd1 _1103_ sky130_fd_sc_hd__a221o_1
X_2456_ hostdisp.curr_word\[25\] net119 vssd1 vssd1 vccd1 vccd1 _1051_ sky130_fd_sc_hd__or2_1
X_1407_ net146 vssd1 vssd1 vccd1 vccd1 _0361_ sky130_fd_sc_hd__inv_2
XANTENNA__3070__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold18 net44 vssd1 vssd1 vccd1 vccd1 net282 sky130_fd_sc_hd__dlygate4sd3_1
Xhold29 net46 vssd1 vssd1 vccd1 vccd1 net293 sky130_fd_sc_hd__dlygate4sd3_1
X_3607__241 vssd1 vssd1 vccd1 vccd1 _3607__241/HI net241 sky130_fd_sc_hd__conb_1
XFILLER_0_39_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2387_ lcdPlayer.cnt_20ms\[15\] lcdPlayer.cnt_20ms\[14\] _1013_ vssd1 vssd1 vccd1
+ vccd1 _1017_ sky130_fd_sc_hd__and3_1
XFILLER_0_127_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3008_ net221 vssd1 vssd1 vccd1 vccd1 _0033_ sky130_fd_sc_hd__inv_2
XFILLER_0_78_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_191_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3614__245 vssd1 vssd1 vccd1 vccd1 _3614__245/HI net245 sky130_fd_sc_hd__conb_1
XFILLER_0_131_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_18_Left_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_150_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3413__CLK clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3234__Q host_message_reg.setLetter\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3563__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3621__249 vssd1 vssd1 vccd1 vccd1 _3621__249/HI net249 sky130_fd_sc_hd__conb_1
XPHY_EDGE_ROW_27_Left_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_139_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_139_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2805__A net142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_36_Left_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_164_Right_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2310_ net74 _0969_ vssd1 vssd1 vccd1 vccd1 _0970_ sky130_fd_sc_hd__nor2_1
X_3290_ clknet_leaf_25_clk net250 net182 vssd1 vssd1 vccd1 vccd1 hostdisp.bottom\[101\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_148_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2241_ lcdPlayer.cnt_500hz\[14\] _0754_ _0932_ vssd1 vssd1 vccd1 vccd1 lcdPlayer.lcd_en
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_57_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2172_ gamelogic.setWord\[20\] _0888_ net132 vssd1 vssd1 vccd1 vccd1 hostdisp.nextBottom\[68\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_23 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_177_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2715__A net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2009__B1 net80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1956_ uart_receiver.bit_index\[2\] net149 net150 vssd1 vssd1 vccd1 vccd1 _0797_
+ sky130_fd_sc_hd__or3_1
XFILLER_0_160_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3319__Q keypadFSMHost.state\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_244 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1887_ uart_transmitter.clk_count\[7\] _0742_ net116 vssd1 vssd1 vccd1 vccd1 _0744_
+ sky130_fd_sc_hd__o21ai_1
XPHY_EDGE_ROW_131_Right_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3557_ clknet_leaf_22_clk net394 net201 vssd1 vssd1 vccd1 vccd1 hostdisp.curr_guesses\[39\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_98_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput19 net19 vssd1 vssd1 vccd1 vccd1 gpio_oeb[27] sky130_fd_sc_hd__buf_2
XFILLER_0_3_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2732__A1 net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2508_ _1061_ _1069_ _1082_ vssd1 vssd1 vccd1 vccd1 _1086_ sky130_fd_sc_hd__and3_4
X_3488_ clknet_leaf_30_clk hostdisp.next_curr_word\[10\] net178 vssd1 vssd1 vccd1
+ vccd1 hostdisp.curr_word\[10\] sky130_fd_sc_hd__dfstp_1
X_2439_ net361 _1041_ net67 vssd1 vssd1 vccd1 vccd1 _0149_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2609__B hostdisp.bottom\[101\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_191_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2420__B1 net69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_159_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_33_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1810_ clock_div.count\[7\] _0700_ vssd1 vssd1 vccd1 vccd1 _0701_ sky130_fd_sc_hd__nand2_1
XFILLER_0_150_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2790_ _0565_ _0601_ _1337_ host_message_reg.setLetter\[6\] vssd1 vssd1 vccd1 vccd1
+ _1338_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_41_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1741_ uart_receiver.clk_count\[5\] uart_receiver.clk_count\[4\] _0646_ vssd1 vssd1
+ vccd1 vccd1 _0649_ sky130_fd_sc_hd__and3_1
XFILLER_0_80_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1672_ _0006_ _0009_ vssd1 vssd1 vccd1 vccd1 keypadFSMHost.next_state\[2\] sky130_fd_sc_hd__or2_1
XANTENNA__2962__A1 gamelogic.setWord\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_282 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3411_ clknet_leaf_20_clk _0300_ net205 vssd1 vssd1 vccd1 vccd1 dispFSM.guesses\[65\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_110_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_34 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3342_ clknet_leaf_31_clk _0231_ net163 vssd1 vssd1 vccd1 vccd1 gamelogic.letter\[4\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_68_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3273_ clknet_leaf_22_clk hostdisp.nextBottom\[71\] net186 vssd1 vssd1 vccd1 vccd1
+ hostdisp.bottom\[71\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_175_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2224_ net122 _0918_ vssd1 vssd1 vccd1 vccd1 _0919_ sky130_fd_sc_hd__nand2_1
X_2155_ gamelogic.setWord\[20\] hostdisp.curr_guesses\[20\] net123 vssd1 vssd1 vccd1
+ vccd1 _0880_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_49_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2086_ hostdisp.curr_word\[25\] hostdisp.curr_word\[27\] _0410_ hostdisp.curr_word\[30\]
+ net101 vssd1 vssd1 vccd1 vccd1 _0847_ sky130_fd_sc_hd__a41o_1
XFILLER_0_75_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_347 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2988_ gamelogic.setWord\[27\] net51 net47 gamelogic.setWord\[35\] vssd1 vssd1 vccd1
+ vccd1 _0351_ sky130_fd_sc_hd__o22a_1
XFILLER_0_16_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_138_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1939_ _0017_ _0766_ vssd1 vssd1 vccd1 vccd1 _0182_ sky130_fd_sc_hd__nor2_1
XFILLER_0_140_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2953__A1 host_message_reg.setLetter\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout115_X net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3609_ gamelogic.green vssd1 vssd1 vccd1 vccd1 net34 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2469__B1 net69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_183_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2641__B1 net110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_11_Right_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_183_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1995__A2 net94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_328 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2944__A1 dispFSM.msg\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_20_Right_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_59 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_167_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1440__Y _0394_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_159_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3281__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2911_ dispFSM.guesses\[51\] net82 net57 net555 vssd1 vssd1 vccd1 vccd1 _0278_ sky130_fd_sc_hd__o22a_1
XANTENNA__2632__B1 _1084_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_199 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_114 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2842_ _1377_ gamelogic.correct\[2\] _1366_ vssd1 vssd1 vccd1 vccd1 _0223_ sky130_fd_sc_hd__mux2_1
X_2773_ net153 _1302_ _1324_ _0560_ vssd1 vssd1 vccd1 vccd1 _1325_ sky130_fd_sc_hd__a22o_1
XFILLER_0_60_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2712__B _1275_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1724_ _0628_ _0634_ _0627_ vssd1 vssd1 vccd1 vccd1 _0639_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_53_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold115 clock_div.count\[16\] vssd1 vssd1 vccd1 vccd1 net379 sky130_fd_sc_hd__dlygate4sd3_1
Xhold126 hostdisp.curr_guesses\[6\] vssd1 vssd1 vccd1 vccd1 net390 sky130_fd_sc_hd__dlygate4sd3_1
Xhold104 hostdisp.top\[48\] vssd1 vssd1 vccd1 vccd1 net368 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1655_ keypadFSMPlayer.state\[5\] _0452_ _0587_ keypadFSMPlayer.state\[2\] vssd1
+ vssd1 vccd1 vccd1 _0016_ sky130_fd_sc_hd__a22o_1
Xhold137 hostdisp.curr_guesses\[45\] vssd1 vssd1 vccd1 vccd1 net401 sky130_fd_sc_hd__dlygate4sd3_1
Xhold159 dispFSM.guesses\[1\] vssd1 vssd1 vccd1 vccd1 net423 sky130_fd_sc_hd__dlygate4sd3_1
Xhold148 hostdisp.top\[41\] vssd1 vssd1 vccd1 vccd1 net412 sky130_fd_sc_hd__dlygate4sd3_1
X_1586_ _0519_ _0529_ _0530_ _0454_ dispFSM.msg\[1\] vssd1 vssd1 vccd1 vccd1 _0059_
+ sky130_fd_sc_hd__o32a_1
XFILLER_0_0_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3325_ clknet_leaf_35_clk _0218_ net161 vssd1 vssd1 vccd1 vccd1 gamelogic.green sky130_fd_sc_hd__dfrtp_1
X_3256_ clknet_leaf_4_clk hostdisp.nextBottom\[54\] net193 vssd1 vssd1 vccd1 vccd1
+ hostdisp.bottom\[54\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2207_ net129 gamelogic.setWord\[38\] vssd1 vssd1 vccd1 vccd1 _0906_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_69_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_185_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3187_ clknet_leaf_29_clk net416 net181 vssd1 vssd1 vccd1 vccd1 hostdisp.top\[71\]
+ sky130_fd_sc_hd__dfrtp_1
X_2138_ gamelogic.setWord\[3\] _0871_ net132 vssd1 vssd1 vccd1 vccd1 hostdisp.nextBottom\[51\]
+ sky130_fd_sc_hd__mux2_1
X_2069_ hostdisp.curr_word\[12\] net102 _0840_ net142 vssd1 vssd1 vccd1 vccd1 hostdisp.next_curr_word\[12\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_48_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout92_A _0824_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_147_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2862__A0 gamelogic.letter\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_158_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2075__D1 gamelogic.indexCorrect\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_171_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1429__A gamelogic.setWord\[37\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_180 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1440_ gamelogic.setWord\[13\] vssd1 vssd1 vccd1 vccd1 _0394_ sky130_fd_sc_hd__inv_2
XFILLER_0_156_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3110_ clknet_leaf_28_clk _0100_ vssd1 vssd1 vccd1 vccd1 lcdPlayer.cnt_500hz\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_65_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3041_ clknet_leaf_8_clk clock_div.next_count\[21\] net213 vssd1 vssd1 vccd1 vccd1
+ clock_div.count\[21\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_164_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2605__B1 net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2081__B2 gamelogic.letter\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2442__B _0827_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2825_ _0928_ _1235_ _1355_ vssd1 vssd1 vccd1 vccd1 _1364_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_170_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2756_ _0565_ _1288_ vssd1 vssd1 vccd1 vccd1 _1310_ sky130_fd_sc_hd__nand2b_2
XTAP_TAPCELL_ROW_135_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3177__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2687_ net144 _0387_ gamelogic.setWord\[30\] _0385_ _1251_ vssd1 vssd1 vccd1 vccd1
+ _1252_ sky130_fd_sc_hd__o221a_1
X_1707_ uart_receiver.bit_index\[2\] net149 net150 vssd1 vssd1 vccd1 vccd1 _0623_
+ sky130_fd_sc_hd__and3_1
X_1638_ _0544_ _0552_ _0367_ vssd1 vssd1 vccd1 vccd1 _0573_ sky130_fd_sc_hd__a21oi_1
X_3569__253 vssd1 vssd1 vccd1 vccd1 net253 _3569__253/LO sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_187_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1569_ _0468_ _0516_ vssd1 vssd1 vccd1 vccd1 _0517_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_6_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3308_ clknet_leaf_34_clk uart_receiver.next_clk_count\[0\] net158 vssd1 vssd1 vccd1
+ vccd1 uart_receiver.clk_count\[0\] sky130_fd_sc_hd__dfrtp_2
X_3239_ clknet_leaf_10_clk keypadFSMHost.next_state\[0\] net215 vssd1 vssd1 vccd1
+ vccd1 _1396_ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_193_255 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout54 _1393_ vssd1 vssd1 vccd1 vccd1 net54 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout65 _1390_ vssd1 vssd1 vccd1 vccd1 net65 sky130_fd_sc_hd__buf_2
XFILLER_0_76_272 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2072__B2 gamelogic.letter\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout87 _0940_ vssd1 vssd1 vccd1 vccd1 net87 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_24_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout98 net100 vssd1 vssd1 vccd1 vccd1 net98 sky130_fd_sc_hd__buf_2
Xfanout76 net77 vssd1 vssd1 vccd1 vccd1 net76 sky130_fd_sc_hd__buf_2
XFILLER_0_91_242 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_153_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3237__Q host_message_reg.setLetter\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout95_X net95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2825__B1_N _1355_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_184_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkload24 clknet_leaf_11_clk vssd1 vssd1 vccd1 vccd1 clkload24/Y sky130_fd_sc_hd__inv_8
XFILLER_0_140_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2610_ hostdisp.bottom\[85\] net117 _1106_ hostdisp.top\[61\] vssd1 vssd1 vccd1 vccd1
+ _1183_ sky130_fd_sc_hd__a22o_1
Xclkload13 clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 clkload13/Y sky130_fd_sc_hd__bufinv_16
XTAP_TAPCELL_ROW_11_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3590_ net262 vssd1 vssd1 vccd1 vccd1 gpio_oeb[23] sky130_fd_sc_hd__buf_2
X_2541_ dispFSM.guesses\[9\] _1078_ net112 dispFSM.guesses\[49\] vssd1 vssd1 vccd1
+ vccd1 _1118_ sky130_fd_sc_hd__a22o_1
XFILLER_0_2_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2472_ hostdisp.curr_word\[36\] net73 net68 net558 vssd1 vssd1 vccd1 vccd1 _0168_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__2118__A2 net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1423_ net145 vssd1 vssd1 vccd1 vccd1 _0377_ sky130_fd_sc_hd__inv_2
XANTENNA__2523__C1 net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_183_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3024_ clknet_leaf_9_clk clock_div.next_count\[4\] net217 vssd1 vssd1 vccd1 vccd1
+ clock_div.count\[4\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_182_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_62_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout142_A gamelogic.letter\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_178_Right_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2054__B2 gamelogic.letter\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload7 clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 clkload7/Y sky130_fd_sc_hd__inv_8
XFILLER_0_41_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2808_ gamelogic.letter\[1\] _0393_ gamelogic.setWord\[15\] _0386_ _1343_ vssd1 vssd1
+ vccd1 vccd1 _1354_ sky130_fd_sc_hd__o221a_1
X_2739_ _0613_ _1292_ keypadFSMHost.state\[3\] vssd1 vssd1 vccd1 vccd1 _1293_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_131_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2599__S net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2109__A2 net96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout222 net223 vssd1 vssd1 vccd1 vccd1 net222 sky130_fd_sc_hd__buf_4
Xfanout211 net212 vssd1 vssd1 vccd1 vccd1 net211 sky130_fd_sc_hd__buf_4
Xfanout200 net224 vssd1 vssd1 vccd1 vccd1 net200 sky130_fd_sc_hd__buf_2
Xfanout233 net5 vssd1 vssd1 vccd1 vccd1 net233 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_5_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3342__CLK clknet_leaf_31_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_181_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_145_Right_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2596__A2 _1086_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3492__CLK clknet_leaf_30_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2348__A2 _0017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2036__A1 gamelogic.letter\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1972_ buffer.Rx_byte\[5\] net2 _0807_ vssd1 vssd1 vccd1 vccd1 _0808_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_173_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_112_Right_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_132_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3573_ net156 vssd1 vssd1 vccd1 vccd1 net25 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_49_Right_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2524_ hostdisp.bottom\[48\] net114 net112 hostdisp.bottom\[72\] vssd1 vssd1 vccd1
+ vccd1 _1102_ sky130_fd_sc_hd__a22o_1
XFILLER_0_121_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2455_ net496 net71 _1050_ _0828_ vssd1 vssd1 vccd1 vccd1 _0156_ sky130_fd_sc_hd__a22o_1
X_1406_ net231 vssd1 vssd1 vccd1 vccd1 _0360_ sky130_fd_sc_hd__clkinv_4
Xhold19 net30 vssd1 vssd1 vccd1 vccd1 net283 sky130_fd_sc_hd__dlygate4sd3_1
X_2386_ lcdPlayer.cnt_20ms\[15\] _1014_ vssd1 vssd1 vccd1 vccd1 _1016_ sky130_fd_sc_hd__or2_1
XANTENNA__2511__A2 net105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_58_Right_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3365__CLK clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3007_ net208 vssd1 vssd1 vccd1 vccd1 _0032_ sky130_fd_sc_hd__inv_2
XANTENNA__3340__Q gamelogic.letter\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_255 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout145_X net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_67_Right_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_150_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_76_Right_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2266__A1 dispFSM.msg\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_120_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3512__SET_B net165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2569__A2 net114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_85_Right_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2240_ lcdPlayer.cnt_500hz\[11\] lcdPlayer.cnt_500hz\[12\] _0931_ lcdPlayer.cnt_500hz\[13\]
+ vssd1 vssd1 vccd1 vccd1 _0932_ sky130_fd_sc_hd__o31a_1
XANTENNA__3388__CLK clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_94_Right_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2171_ gamelogic.setWord\[28\] hostdisp.curr_guesses\[28\] net123 vssd1 vssd1 vccd1
+ vccd1 _0888_ sky130_fd_sc_hd__mux2_1
XFILLER_0_189_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_35 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3160__Q hostdisp.top\[44\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1955_ host_message_reg.Cstate net97 _0607_ vssd1 vssd1 vccd1 vccd1 host_message_reg.next_state
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_7_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_1_Left_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1886_ _0742_ _0743_ vssd1 vssd1 vccd1 vccd1 uart_transmitter.next_clk_count\[6\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_113_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_256 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3556_ clknet_leaf_6_clk hostdisp.next_curr_guesses\[38\] net192 vssd1 vssd1 vccd1
+ vccd1 hostdisp.curr_guesses\[38\] sky130_fd_sc_hd__dfstp_1
XFILLER_0_113_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2193__A0 gamelogic.setWord\[39\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout105_A _1081_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2507_ _1060_ _1071_ vssd1 vssd1 vccd1 vccd1 _1085_ sky130_fd_sc_hd__nor2_2
XFILLER_0_51_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3487_ clknet_leaf_30_clk hostdisp.next_curr_word\[9\] net178 vssd1 vssd1 vccd1 vccd1
+ hostdisp.curr_word\[9\] sky130_fd_sc_hd__dfstp_1
X_2438_ net130 host_message_reg.setLetter\[1\] hostdisp.curr_word\[17\] _0830_ _1034_
+ vssd1 vssd1 vccd1 vccd1 _1041_ sky130_fd_sc_hd__a221o_1
X_2369_ net358 _1002_ net167 vssd1 vssd1 vccd1 vccd1 _1005_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_168_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_307 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_280 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2420__B2 hostdisp.top\[46\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3530__CLK clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3169__RESET_B net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2487__B2 net139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_174_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1998__B1 net77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_175 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_318 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_239 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1740_ net338 _0646_ _0648_ vssd1 vssd1 vccd1 vccd1 uart_receiver.next_clk_count\[4\]
+ sky130_fd_sc_hd__a21oi_1
XANTENNA__1438__Y _0392_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1671_ _0537_ _0593_ _0594_ _0592_ keypadFSMHost.state\[4\] vssd1 vssd1 vccd1 vccd1
+ _0009_ sky130_fd_sc_hd__a32o_1
XFILLER_0_7_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3410_ clknet_leaf_23_clk _0299_ net187 vssd1 vssd1 vccd1 vccd1 dispFSM.guesses\[64\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_150_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3341_ clknet_leaf_35_clk _0230_ net162 vssd1 vssd1 vccd1 vccd1 gamelogic.letter\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_68_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_90_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3272_ clknet_leaf_1_clk hostdisp.nextBottom\[70\] net176 vssd1 vssd1 vccd1 vccd1
+ hostdisp.bottom\[70\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_175_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2223_ _0909_ _0912_ _0915_ vssd1 vssd1 vccd1 vccd1 _0918_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_84_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_49_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2154_ gamelogic.setWord\[11\] _0879_ net131 vssd1 vssd1 vccd1 vccd1 hostdisp.nextBottom\[59\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_177_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2085_ hostdisp.curr_word\[23\] net97 _0846_ net140 vssd1 vssd1 vccd1 vccd1 hostdisp.next_curr_word\[23\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_191_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2650__A1 hostdisp.top\[47\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_192_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_99_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2987_ gamelogic.setWord\[26\] net51 net47 gamelogic.setWord\[34\] vssd1 vssd1 vccd1
+ vccd1 _0350_ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout222_A net223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1938_ _0784_ _0785_ _0779_ _0781_ vssd1 vssd1 vccd1 vccd1 _0000_ sky130_fd_sc_hd__a2bb2o_1
X_1869_ uart_transmitter.clk_count\[0\] net116 vssd1 vssd1 vccd1 vccd1 uart_transmitter.next_clk_count\[0\]
+ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_138_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2953__A2 net53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3608_ message_reg.blue vssd1 vssd1 vccd1 vccd1 net33 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3065__Q dispFSM.msg\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout108_X net108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3539_ clknet_leaf_14_clk hostdisp.next_curr_guesses\[21\] net208 vssd1 vssd1 vccd1
+ vccd1 hostdisp.curr_guesses\[21\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__3262__RESET_B net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_55_Left_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_149_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3083__CLK clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_64_Left_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2157__A0 gamelogic.setWord\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_73_Left_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3426__CLK clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload0_A clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_82_Left_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_161_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_159_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2910_ dispFSM.guesses\[50\] net83 net59 net529 vssd1 vssd1 vccd1 vccd1 _0277_ sky130_fd_sc_hd__o22a_1
XFILLER_0_97_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_123 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2841_ _1375_ _1376_ _0815_ vssd1 vssd1 vccd1 vccd1 _1377_ sky130_fd_sc_hd__o21a_1
XFILLER_0_72_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2772_ _0553_ _0558_ _1323_ _1305_ vssd1 vssd1 vccd1 vccd1 _1324_ sky130_fd_sc_hd__a31o_1
XANTENNA__1609__B net3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1723_ _0624_ _0629_ _0632_ _0638_ vssd1 vssd1 vccd1 vccd1 uart_receiver.next_state\[0\]
+ sky130_fd_sc_hd__or4_1
XFILLER_0_53_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold116 keypadFSMPlayer.unlocked vssd1 vssd1 vccd1 vccd1 net380 sky130_fd_sc_hd__dlygate4sd3_1
Xhold105 keypadFSMPlayer.prev_key\[5\] vssd1 vssd1 vccd1 vccd1 net369 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_91_Left_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1654_ _0451_ _0489_ vssd1 vssd1 vccd1 vccd1 _0587_ sky130_fd_sc_hd__and2_1
Xhold138 clock_div.count\[19\] vssd1 vssd1 vccd1 vccd1 net402 sky130_fd_sc_hd__dlygate4sd3_1
Xhold127 hostdisp.curr_guesses\[29\] vssd1 vssd1 vccd1 vccd1 net391 sky130_fd_sc_hd__dlygate4sd3_1
Xhold149 dispFSM.guesses\[6\] vssd1 vssd1 vccd1 vccd1 net413 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1585_ dispFSM.msg\[1\] _0447_ vssd1 vssd1 vccd1 vccd1 _0530_ sky130_fd_sc_hd__and2_1
XFILLER_0_21_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3324_ clknet_leaf_10_clk _0010_ net218 vssd1 vssd1 vccd1 vccd1 keypadFSMHost.state\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3255_ clknet_leaf_15_clk hostdisp.nextBottom\[53\] net207 vssd1 vssd1 vccd1 vccd1
+ hostdisp.bottom\[53\] sky130_fd_sc_hd__dfrtp_1
X_2206_ net129 net401 net120 _0905_ vssd1 vssd1 vccd1 vccd1 hostdisp.nextBottom\[85\]
+ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_185_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3186_ clknet_leaf_4_clk _0162_ net177 vssd1 vssd1 vccd1 vccd1 hostdisp.top\[70\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_178_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2137_ gamelogic.setWord\[11\] hostdisp.curr_guesses\[11\] net121 vssd1 vssd1 vccd1
+ vccd1 _0871_ sky130_fd_sc_hd__mux2_1
X_2068_ hostdisp.curr_word\[11\] net102 _0840_ gamelogic.letter\[3\] vssd1 vssd1 vccd1
+ vccd1 hostdisp.next_curr_word\[11\] sky130_fd_sc_hd__o22a_1
XFILLER_0_138_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2623__A1 net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1831__C1 _0693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_173_172 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout225_X net225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_9_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3449__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_0_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_158_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_164_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_156_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2550__B1 net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3040_ clknet_leaf_8_clk clock_div.next_count\[20\] net213 vssd1 vssd1 vccd1 vccd1
+ clock_div.count\[20\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_65_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_172_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_159_Right_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_157_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2824_ net311 _1362_ _1363_ vssd1 vssd1 vccd1 vccd1 _0219_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_14_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_164 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2755_ _0597_ _1308_ _0603_ vssd1 vssd1 vccd1 vccd1 _1309_ sky130_fd_sc_hd__o21bai_1
XTAP_TAPCELL_ROW_135_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2686_ net143 gamelogic.setWord\[27\] vssd1 vssd1 vccd1 vccd1 _1251_ sky130_fd_sc_hd__xnor2_1
X_1706_ net149 net150 _0621_ vssd1 vssd1 vccd1 vccd1 _0622_ sky130_fd_sc_hd__and3_1
X_1637_ keypadFSMHost.prev_key\[0\] _0554_ vssd1 vssd1 vccd1 vccd1 _0572_ sky130_fd_sc_hd__xor2_1
X_1568_ _0499_ _0515_ _0512_ vssd1 vssd1 vccd1 vccd1 _0516_ sky130_fd_sc_hd__or3b_1
XANTENNA__2541__B1 net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3307_ clknet_leaf_33_clk uart_receiver.temp_byte\[7\] net158 vssd1 vssd1 vccd1 vccd1
+ buffer.Rx_byte\[7\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__3343__Q gamelogic.letter\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1499_ _0434_ _0450_ vssd1 vssd1 vccd1 vccd1 _0451_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_129_Left_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3238_ clknet_leaf_13_clk _0212_ net208 vssd1 vssd1 vccd1 vccd1 host_message_reg.setLetter\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_3169_ clknet_leaf_30_clk _0145_ net184 vssd1 vssd1 vccd1 vccd1 hostdisp.top\[53\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_126_Right_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_65_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_193_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_267 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_138_Left_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout55 _1392_ vssd1 vssd1 vccd1 vccd1 net55 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_119_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2072__A2 net96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2125__S net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout88 net89 vssd1 vssd1 vccd1 vccd1 net88 sky130_fd_sc_hd__buf_2
Xfanout77 _0826_ vssd1 vssd1 vccd1 vccd1 net77 sky130_fd_sc_hd__clkbuf_4
Xfanout66 _1235_ vssd1 vssd1 vccd1 vccd1 net66 sky130_fd_sc_hd__clkbuf_2
Xfanout99 net100 vssd1 vssd1 vccd1 vccd1 net99 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_91_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_153_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_147_Left_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_169_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_156_Left_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_123_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_184_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_184_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload25 clknet_leaf_12_clk vssd1 vssd1 vccd1 vccd1 clkload25/Y sky130_fd_sc_hd__clkinv_8
XFILLER_0_125_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_11_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload14 clknet_leaf_25_clk vssd1 vssd1 vccd1 vccd1 clkload14/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_152_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2540_ dispFSM.guesses\[73\] _1086_ net110 dispFSM.guesses\[33\] _1116_ vssd1 vssd1
+ vccd1 vccd1 _1117_ sky130_fd_sc_hd__a221o_1
X_2471_ hostdisp.curr_word\[35\] net75 net68 net490 _1034_ vssd1 vssd1 vccd1 vccd1
+ _0167_ sky130_fd_sc_hd__a221o_1
XFILLER_0_167_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1422_ gamelogic.setWord\[32\] vssd1 vssd1 vccd1 vccd1 _0376_ sky130_fd_sc_hd__inv_2
XFILLER_0_50_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2523__B1 _1085_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3163__Q hostdisp.top\[47\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3023_ clknet_leaf_9_clk clock_div.next_count\[3\] net217 vssd1 vssd1 vccd1 vccd1
+ clock_div.count\[3\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__2826__A1 gamelogic.indexCorrect\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_183_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_182_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_175_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_62_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_141_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout135_A net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload8 clknet_leaf_32_clk vssd1 vssd1 vccd1 vccd1 clkload8/Y sky130_fd_sc_hd__inv_16
X_2807_ _1348_ _1349_ _1352_ vssd1 vssd1 vccd1 vccd1 _1353_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_14_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3338__Q gamelogic.letter\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3294__CLK clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2738_ _0369_ _1291_ keypadFSMHost.state\[2\] vssd1 vssd1 vccd1 vccd1 _1292_ sky130_fd_sc_hd__a21o_1
XFILLER_0_14_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1565__A1 net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2669_ net96 _0909_ vssd1 vssd1 vccd1 vccd1 _1235_ sky130_fd_sc_hd__or2_1
Xfanout223 net224 vssd1 vssd1 vccd1 vccd1 net223 sky130_fd_sc_hd__buf_4
Xfanout212 net224 vssd1 vssd1 vccd1 vccd1 net212 sky130_fd_sc_hd__clkbuf_2
Xfanout201 net202 vssd1 vssd1 vccd1 vccd1 net201 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_1_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout48_A net50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_346 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2450__C1 net71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3535__SET_B net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2808__A1 gamelogic.letter\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3167__CLK clknet_leaf_30_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1971_ uart_receiver.bit_index\[1\] net150 uart_receiver.bit_index\[2\] vssd1 vssd1
+ vccd1 vccd1 _0807_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_173_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_54 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3572_ net256 vssd1 vssd1 vccd1 vccd1 gpio_oeb[5] sky130_fd_sc_hd__buf_2
X_2523_ hostdisp.bottom\[40\] _1081_ _1085_ hostdisp.bottom\[64\] net227 vssd1 vssd1
+ vccd1 vccd1 _1101_ sky130_fd_sc_hd__a221o_1
XFILLER_0_11_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2454_ hostdisp.curr_word\[24\] net119 vssd1 vssd1 vccd1 vccd1 _1050_ sky130_fd_sc_hd__or2_1
X_1405_ keypadFSMPlayer.prev_key\[6\] vssd1 vssd1 vccd1 vccd1 _0359_ sky130_fd_sc_hd__inv_2
X_2385_ _1014_ _1015_ vssd1 vssd1 vccd1 vccd1 _0121_ sky130_fd_sc_hd__nor2_1
XFILLER_0_127_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput1 en vssd1 vssd1 vccd1 vccd1 net1 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_143_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3270__D hostdisp.nextBottom\[68\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3006_ net208 vssd1 vssd1 vccd1 vccd1 _0031_ sky130_fd_sc_hd__inv_2
XFILLER_0_78_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_148_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_267 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_163_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3068__Q dispFSM.msg\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2983__B1 net49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_150_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_161_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_204 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2423__C1 _1034_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2170_ gamelogic.setWord\[19\] _0887_ net131 vssd1 vssd1 vccd1 vccd1 hostdisp.nextBottom\[67\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_164_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_177_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1465__B1 net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_180_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2009__A2 _0823_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1954_ _0770_ _0777_ _0789_ _0795_ _0778_ vssd1 vssd1 vccd1 vccd1 _0004_ sky130_fd_sc_hd__a32o_1
XFILLER_0_113_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_189_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1885_ uart_transmitter.clk_count\[6\] _0740_ net116 vssd1 vssd1 vccd1 vccd1 _0743_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_43_268 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3555_ clknet_leaf_14_clk hostdisp.next_curr_guesses\[37\] net207 vssd1 vssd1 vccd1
+ vccd1 hostdisp.curr_guesses\[37\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_113_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2506_ _1069_ _1083_ vssd1 vssd1 vccd1 vccd1 _1084_ sky130_fd_sc_hd__and2_4
X_3486_ clknet_leaf_4_clk hostdisp.next_curr_word\[8\] net178 vssd1 vssd1 vccd1 vccd1
+ hostdisp.curr_word\[8\] sky130_fd_sc_hd__dfstp_1
X_2437_ net314 _1033_ _1040_ vssd1 vssd1 vccd1 vccd1 _0148_ sky130_fd_sc_hd__o21a_1
XANTENNA__3332__CLK clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_102_Left_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2368_ lcdPlayer.cnt_20ms\[9\] lcdPlayer.cnt_20ms\[8\] _1000_ vssd1 vssd1 vccd1 vccd1
+ _1004_ sky130_fd_sc_hd__and3_1
X_2299_ _0957_ _0962_ vssd1 vssd1 vccd1 vccd1 _0088_ sky130_fd_sc_hd__nor2_1
XFILLER_0_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3050__RESET_B net221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_24_clk_X clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2956__B1 net48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2133__S net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout70_X net70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2287__A_N net106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_187 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3205__CLK clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_182_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1670_ _0537_ _0594_ vssd1 vssd1 vccd1 vccd1 _0595_ sky130_fd_sc_hd__nand2_1
XFILLER_0_135_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3355__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3340_ clknet_leaf_33_clk _0229_ net162 vssd1 vssd1 vccd1 vccd1 gamelogic.letter\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_0_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_90_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3271_ clknet_leaf_15_clk hostdisp.nextBottom\[69\] net209 vssd1 vssd1 vccd1 vccd1
+ hostdisp.bottom\[69\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_187_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2222_ net100 _0909_ _0917_ vssd1 vssd1 vccd1 vccd1 gamelogic.nextState\[0\] sky130_fd_sc_hd__o21ai_1
XFILLER_0_108_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2153_ gamelogic.setWord\[19\] hostdisp.curr_guesses\[19\] net121 vssd1 vssd1 vccd1
+ vccd1 _0879_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2084_ hostdisp.curr_word\[22\] net103 _0845_ gamelogic.letter\[6\] vssd1 vssd1 vccd1
+ vccd1 hostdisp.next_curr_word\[22\] sky130_fd_sc_hd__o22a_1
XFILLER_0_191_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_158_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2650__A2 _1098_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_185_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2986_ gamelogic.setWord\[25\] net54 net49 gamelogic.setWord\[33\] vssd1 vssd1 vccd1
+ vccd1 _0349_ sky130_fd_sc_hd__o22a_1
XFILLER_0_133_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1937_ _0771_ _0780_ _0783_ _0187_ vssd1 vssd1 vccd1 vccd1 _0785_ sky130_fd_sc_hd__a31o_1
XFILLER_0_71_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2461__B _0827_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout215_A net218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1868_ _0662_ _0671_ _0664_ vssd1 vssd1 vccd1 vccd1 _0732_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_138_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3607_ net241 vssd1 vssd1 vccd1 vccd1 gpio_out[15] sky130_fd_sc_hd__buf_2
XFILLER_0_101_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1799_ clock_div.count\[1\] clock_div.count\[0\] net448 vssd1 vssd1 vccd1 vccd1 _0695_
+ sky130_fd_sc_hd__a21oi_1
X_3538_ clknet_leaf_1_clk hostdisp.next_curr_guesses\[20\] net176 vssd1 vssd1 vccd1
+ vccd1 hostdisp.curr_guesses\[20\] sky130_fd_sc_hd__dfstp_1
X_3469_ clknet_leaf_14_clk _0347_ net194 vssd1 vssd1 vccd1 vccd1 gamelogic.setWord\[31\]
+ sky130_fd_sc_hd__dfrtp_4
XPHY_EDGE_ROW_110_Left_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2641__A2 net105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3378__CLK clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_156_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_19_clk_A clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_135 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2632__A2 net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2840_ _1370_ _1371_ _1374_ vssd1 vssd1 vccd1 vccd1 _1376_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_72_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2771_ net152 net151 _0546_ _0362_ vssd1 vssd1 vccd1 vccd1 _1323_ sky130_fd_sc_hd__o211a_1
XFILLER_0_155_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1722_ _0634_ _0637_ vssd1 vssd1 vccd1 vccd1 _0638_ sky130_fd_sc_hd__nor2_1
XFILLER_0_53_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1653_ message_reg.state\[0\] message_reg.state\[1\] vssd1 vssd1 vccd1 vccd1 message_reg.blue
+ sky130_fd_sc_hd__and2_1
Xhold117 hostdisp.curr_guesses\[15\] vssd1 vssd1 vccd1 vccd1 net381 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold106 lcdPlayer.cnt_20ms\[6\] vssd1 vssd1 vccd1 vccd1 net370 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold128 hostdisp.next_curr_guesses\[29\] vssd1 vssd1 vccd1 vccd1 net392 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_9_Right_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1906__A _0752_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold139 hostdisp.curr_word\[37\] vssd1 vssd1 vccd1 vccd1 net403 sky130_fd_sc_hd__dlygate4sd3_1
X_1584_ _0450_ _0528_ vssd1 vssd1 vccd1 vccd1 _0529_ sky130_fd_sc_hd__and2b_1
X_3323_ clknet_leaf_10_clk _0009_ net215 vssd1 vssd1 vccd1 vccd1 keypadFSMHost.state\[4\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_119_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_107_Right_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3254_ clknet_leaf_3_clk hostdisp.nextBottom\[52\] net177 vssd1 vssd1 vccd1 vccd1
+ hostdisp.bottom\[52\] sky130_fd_sc_hd__dfrtp_1
X_2205_ net137 gamelogic.setWord\[37\] vssd1 vssd1 vccd1 vccd1 _0905_ sky130_fd_sc_hd__or2_1
XFILLER_0_28_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_185_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3185_ clknet_leaf_30_clk _0161_ net184 vssd1 vssd1 vccd1 vccd1 hostdisp.top\[69\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__2456__B net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2136_ gamelogic.setWord\[2\] _0870_ net132 vssd1 vssd1 vccd1 vccd1 hostdisp.nextBottom\[50\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout165_A net225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2067_ hostdisp.curr_word\[10\] net102 _0840_ gamelogic.letter\[2\] vssd1 vssd1 vccd1
+ vccd1 hostdisp.next_curr_word\[10\] sky130_fd_sc_hd__o22a_1
XFILLER_0_193_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3520__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_151_83 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2969_ gamelogic.setWord\[8\] net53 net49 gamelogic.setWord\[16\] vssd1 vssd1 vccd1
+ vccd1 _0332_ sky130_fd_sc_hd__o22a_1
XFILLER_0_8_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_330 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout218_X net218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout120_X net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1816__A _0693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3290__250 vssd1 vssd1 vccd1 vccd1 net250 _3290__250/LO sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_9_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_90 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout78_A net79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2075__B1 net75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_0_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_158_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3543__CLK clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2605__A2 _1072_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_176_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2823_ net100 _0827_ net122 _0909_ vssd1 vssd1 vccd1 vccd1 _1363_ sky130_fd_sc_hd__or4_1
XFILLER_0_170_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2754_ _1301_ _1307_ vssd1 vssd1 vccd1 vccd1 _1308_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_143_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_300 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_176 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1705_ uart_receiver.clk_count\[9\] uart_receiver.clk_count\[8\] _0620_ uart_receiver.clk_count\[10\]
+ vssd1 vssd1 vccd1 vccd1 _0621_ sky130_fd_sc_hd__o31a_2
XTAP_TAPCELL_ROW_135_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2685_ _0385_ gamelogic.setWord\[30\] vssd1 vssd1 vccd1 vccd1 _1250_ sky130_fd_sc_hd__nand2_1
X_1636_ keypadFSMHost.prev_key\[1\] _0546_ net152 vssd1 vssd1 vccd1 vccd1 _0571_ sky130_fd_sc_hd__and3b_1
X_1567_ _0499_ _0514_ vssd1 vssd1 vccd1 vccd1 _0515_ sky130_fd_sc_hd__xnor2_1
X_3306_ clknet_leaf_33_clk uart_receiver.temp_byte\[6\] net160 vssd1 vssd1 vccd1 vccd1
+ buffer.Rx_byte\[6\] sky130_fd_sc_hd__dfrtp_1
X_1498_ _0442_ _0449_ vssd1 vssd1 vccd1 vccd1 _0450_ sky130_fd_sc_hd__or2_1
X_3237_ clknet_leaf_12_clk _0211_ net215 vssd1 vssd1 vccd1 vccd1 host_message_reg.setLetter\[6\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_146_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3168_ clknet_leaf_30_clk _0144_ net178 vssd1 vssd1 vccd1 vccd1 hostdisp.top\[52\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_65_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2119_ gamelogic.setWord\[2\] net121 vssd1 vssd1 vccd1 vccd1 _0862_ sky130_fd_sc_hd__or2_1
XFILLER_0_166_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3099_ clknet_leaf_27_clk _0089_ vssd1 vssd1 vccd1 vccd1 lcdPlayer.cnt_500hz\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout56 net59 vssd1 vssd1 vccd1 vccd1 net56 sky130_fd_sc_hd__buf_2
XFILLER_0_193_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout78 net79 vssd1 vssd1 vccd1 vccd1 net78 sky130_fd_sc_hd__clkbuf_4
Xfanout89 _0939_ vssd1 vssd1 vccd1 vccd1 net89 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout67 _1033_ vssd1 vssd1 vccd1 vccd1 net67 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_91_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_153_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2141__S net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3566__CLK clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_123_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2048__B1 net75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3001__A net221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_152_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload26 clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 clkload26/Y sky130_fd_sc_hd__inv_4
Xclkload15 clknet_leaf_26_clk vssd1 vssd1 vccd1 vccd1 clkload15/Y sky130_fd_sc_hd__clkinv_8
XTAP_TAPCELL_ROW_11_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2470_ hostdisp.curr_word\[34\] net75 net68 net470 _1034_ vssd1 vssd1 vccd1 vccd1
+ _0166_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_192_Right_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_167_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1421_ net137 vssd1 vssd1 vccd1 vccd1 _0375_ sky130_fd_sc_hd__inv_2
XFILLER_0_183_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3022_ clknet_leaf_10_clk clock_div.next_count\[2\] net217 vssd1 vssd1 vccd1 vccd1
+ clock_div.count\[2\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_87_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_182_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_175_202 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2039__B1 net80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_141_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_173 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload9 clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 clkload9/Y sky130_fd_sc_hd__bufinv_16
X_2806_ gamelogic.letter\[5\] _0394_ _1350_ _1351_ gamelogic.indexCorrect\[1\] vssd1
+ vssd1 vccd1 vccd1 _1352_ sky130_fd_sc_hd__a221o_1
X_2737_ _0395_ _1396_ keypadFSMHost.state\[1\] vssd1 vssd1 vccd1 vccd1 _1291_ sky130_fd_sc_hd__a21o_1
XANTENNA__2211__A0 _0607_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2668_ net339 _0665_ _1234_ vssd1 vssd1 vccd1 vccd1 _0192_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_14_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1619_ _0542_ _0545_ keypadHostt.scan_col\[0\] vssd1 vssd1 vccd1 vccd1 _0554_ sky130_fd_sc_hd__o21a_1
Xfanout213 net218 vssd1 vssd1 vccd1 vccd1 net213 sky130_fd_sc_hd__clkbuf_4
Xfanout202 net206 vssd1 vssd1 vccd1 vccd1 net202 sky130_fd_sc_hd__clkbuf_4
X_2599_ hostdisp.bottom\[68\] dispFSM.guesses\[44\] net228 vssd1 vssd1 vccd1 vccd1
+ _1173_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout224 net225 vssd1 vssd1 vccd1 vccd1 net224 sky130_fd_sc_hd__clkbuf_4
XANTENNA__2197__A net130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input2_A gpio_in[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_166_202 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_166_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2136__S net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_181_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2450__B1 _0828_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_170_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_16_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1970_ _0618_ _0806_ vssd1 vssd1 vccd1 vccd1 uart_receiver.temp_byte\[4\] sky130_fd_sc_hd__and2_1
XFILLER_0_55_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_173_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3439__Q gamelogic.setWord\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3515__RESET_B net169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_154 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2992__B2 gamelogic.setWord\[39\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2992__A1 gamelogic.setWord\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_176 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_66 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3571_ net255 vssd1 vssd1 vccd1 vccd1 gpio_oeb[4] sky130_fd_sc_hd__buf_2
XFILLER_0_178_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2522_ hostdisp.bottom\[80\] net118 net109 hostdisp.bottom\[56\] _1099_ vssd1 vssd1
+ vccd1 vccd1 _1100_ sky130_fd_sc_hd__a221o_1
XFILLER_0_113_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_93_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2453_ net349 net67 _1049_ vssd1 vssd1 vccd1 vccd1 _0155_ sky130_fd_sc_hd__o21a_1
X_1404_ net269 vssd1 vssd1 vccd1 vccd1 _0358_ sky130_fd_sc_hd__inv_2
X_2384_ net427 _1013_ net182 vssd1 vssd1 vccd1 vccd1 _1015_ sky130_fd_sc_hd__o21ai_1
Xinput2 gpio_in[20] vssd1 vssd1 vccd1 vccd1 net2 sky130_fd_sc_hd__buf_2
X_3005_ net219 vssd1 vssd1 vccd1 vccd1 _0030_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_143_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2680__B1 gamelogic.setWord\[39\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3261__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_148_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_163_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_175_Left_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout200_X net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_150_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_179 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2499__B1 net114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_184_Left_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_161_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_358 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_193_Left_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2423__B1 net70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2974__B2 gamelogic.setWord\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_148_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3284__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_180_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_227 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2414__B1 net69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1953_ _0778_ _0795_ _0796_ _0773_ vssd1 vssd1 vccd1 vccd1 _0003_ sky130_fd_sc_hd__a22o_1
XFILLER_0_90_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1884_ uart_transmitter.clk_count\[6\] _0740_ vssd1 vssd1 vccd1 vccd1 _0742_ sky130_fd_sc_hd__and2_1
XFILLER_0_138_290 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_190_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_189_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3554_ clknet_leaf_1_clk hostdisp.next_curr_guesses\[36\] net179 vssd1 vssd1 vccd1
+ vccd1 hostdisp.curr_guesses\[36\] sky130_fd_sc_hd__dfstp_1
XFILLER_0_11_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3485_ clknet_leaf_28_clk hostdisp.next_curr_word\[7\] net166 vssd1 vssd1 vccd1 vccd1
+ hostdisp.curr_word\[7\] sky130_fd_sc_hd__dfrtp_1
X_2505_ lcdPlayer.nextState\[5\] lcdPlayer.nextState\[4\] _1082_ vssd1 vssd1 vccd1
+ vccd1 _1083_ sky130_fd_sc_hd__and3_1
X_2436_ net129 host_message_reg.setLetter\[0\] _0828_ _1039_ net70 vssd1 vssd1 vccd1
+ vccd1 _1040_ sky130_fd_sc_hd__a221o_1
XFILLER_0_138_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2367_ _1002_ _1003_ vssd1 vssd1 vccd1 vccd1 _0115_ sky130_fd_sc_hd__nor2_1
X_2298_ lcdPlayer.cnt_500hz\[5\] _0752_ vssd1 vssd1 vccd1 vccd1 _0962_ sky130_fd_sc_hd__xor2_1
XFILLER_0_154_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2653__B1 net110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2956__A1 host_message_reg.setLetter\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_109_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1998__A2 net92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_182_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_159_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3270_ clknet_leaf_22_clk hostdisp.nextBottom\[68\] net186 vssd1 vssd1 vccd1 vccd1
+ hostdisp.bottom\[68\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_90_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2221_ _0912_ _0915_ _0916_ gamelogic.state\[0\] _0814_ vssd1 vssd1 vccd1 vccd1 _0917_
+ sky130_fd_sc_hd__o221a_1
X_2152_ gamelogic.setWord\[10\] _0878_ net131 vssd1 vssd1 vccd1 vccd1 hostdisp.nextBottom\[58\]
+ sky130_fd_sc_hd__mux2_1
X_2083_ net568 net97 _0846_ net141 vssd1 vssd1 vccd1 vccd1 hostdisp.next_curr_word\[21\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__1911__B _0752_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_191_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2635__B1 net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_158_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2985_ gamelogic.setWord\[24\] net53 net49 gamelogic.setWord\[32\] vssd1 vssd1 vccd1
+ vccd1 _0348_ sky130_fd_sc_hd__o22a_1
XFILLER_0_90_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1936_ _0771_ _0780_ _0783_ vssd1 vssd1 vccd1 vccd1 _0784_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_83_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1867_ keypadHostt.scan_col\[3\] net146 net230 vssd1 vssd1 vccd1 vccd1 net42 sky130_fd_sc_hd__mux2_1
XANTENNA__1610__A1 net4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3606_ net240 vssd1 vssd1 vccd1 vccd1 gpio_out[14] sky130_fd_sc_hd__buf_2
X_1798_ clock_div.count\[1\] clock_div.count\[0\] clock_div.count\[2\] vssd1 vssd1
+ vccd1 vccd1 _0694_ sky130_fd_sc_hd__and3_1
X_3537_ clknet_leaf_0_clk hostdisp.next_curr_guesses\[19\] net170 vssd1 vssd1 vccd1
+ vccd1 hostdisp.curr_guesses\[19\] sky130_fd_sc_hd__dfstp_1
X_3468_ clknet_leaf_6_clk _0346_ net191 vssd1 vssd1 vccd1 vccd1 gamelogic.setWord\[30\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_58_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_149_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3399_ clknet_leaf_22_clk net389 net201 vssd1 vssd1 vccd1 vccd1 dispFSM.guesses\[53\]
+ sky130_fd_sc_hd__dfrtp_1
X_2419_ hostdisp.curr_word\[5\] _1031_ net67 net277 vssd1 vssd1 vccd1 vccd1 _0137_
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_98_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_181_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2144__S net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_156_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_126_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2617__B1 _1095_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2093__B2 gamelogic.letter\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_147 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2770_ host_message_reg.setLetter\[1\] _1290_ _1322_ vssd1 vssd1 vccd1 vccd1 _0206_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_115_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1721_ uart_receiver.clk_count\[8\] _0620_ _0635_ _0636_ vssd1 vssd1 vccd1 vccd1
+ _0637_ sky130_fd_sc_hd__or4_1
X_1652_ keypadFSMHost.state\[1\] _0565_ _0586_ vssd1 vssd1 vccd1 vccd1 _0006_ sky130_fd_sc_hd__a21o_1
XFILLER_0_13_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold107 hostdisp.top\[67\] vssd1 vssd1 vccd1 vccd1 net371 sky130_fd_sc_hd__dlygate4sd3_1
Xhold118 hostdisp.next_curr_guesses\[15\] vssd1 vssd1 vccd1 vccd1 net382 sky130_fd_sc_hd__dlygate4sd3_1
Xhold129 hostdisp.curr_guesses\[39\] vssd1 vssd1 vccd1 vccd1 net393 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1906__B _0758_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_186_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1583_ _0527_ _0502_ _0499_ vssd1 vssd1 vccd1 vccd1 _0528_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3322_ clknet_leaf_10_clk _0008_ net215 vssd1 vssd1 vccd1 vccd1 keypadFSMHost.state\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_3253_ clknet_leaf_3_clk hostdisp.nextBottom\[51\] net174 vssd1 vssd1 vccd1 vccd1
+ hostdisp.bottom\[51\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_23_clk_X clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2204_ net132 hostdisp.curr_guesses\[44\] net121 _0904_ vssd1 vssd1 vccd1 vccd1 hostdisp.nextBottom\[84\]
+ sky130_fd_sc_hd__a31o_1
X_3184_ clknet_leaf_4_clk _0160_ net178 vssd1 vssd1 vccd1 vccd1 hostdisp.top\[68\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__2856__A0 net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_185_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2135_ gamelogic.setWord\[10\] hostdisp.curr_guesses\[10\] net122 vssd1 vssd1 vccd1
+ vccd1 _0870_ sky130_fd_sc_hd__mux2_1
X_2066_ hostdisp.curr_word\[9\] net101 _0840_ net144 vssd1 vssd1 vccd1 vccd1 hostdisp.next_curr_word\[9\]
+ sky130_fd_sc_hd__o22a_1
XANTENNA__2084__B2 gamelogic.letter\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_171 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2968_ gamelogic.setWord\[7\] net55 _1394_ gamelogic.setWord\[15\] vssd1 vssd1 vccd1
+ vccd1 _0331_ sky130_fd_sc_hd__a22o_1
XFILLER_0_8_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_342 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_139 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1919_ _0770_ vssd1 vssd1 vccd1 vccd1 _0184_ sky130_fd_sc_hd__inv_2
X_2899_ dispFSM.guesses\[39\] net88 net65 net450 vssd1 vssd1 vccd1 vccd1 _0266_ sky130_fd_sc_hd__a22o_1
XFILLER_0_114_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout113_X net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2139__S net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3345__CLK clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_0_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_158_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_173_Right_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2950__X _1393_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3495__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2550__A2 net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3122__RESET_B net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2066__B2 net144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_176_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2822_ _0827_ _0910_ _1362_ net364 vssd1 vssd1 vccd1 vccd1 _0218_ sky130_fd_sc_hd__a22o_1
X_2753_ _0560_ _1304_ _1306_ _1302_ vssd1 vssd1 vccd1 vccd1 _1307_ sky130_fd_sc_hd__a31oi_2
XPHY_EDGE_ROW_140_Right_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_14_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_312 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1704_ uart_receiver.clk_count\[6\] uart_receiver.clk_count\[7\] uart_receiver.clk_count\[5\]
+ uart_receiver.clk_count\[4\] vssd1 vssd1 vccd1 vccd1 _0620_ sky130_fd_sc_hd__or4_1
XFILLER_0_170_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2684_ gamelogic.indexCorrect\[4\] _1249_ _1236_ vssd1 vssd1 vccd1 vccd1 _0193_ sky130_fd_sc_hd__o21a_1
X_1635_ net151 _0546_ keypadFSMHost.prev_key\[2\] vssd1 vssd1 vccd1 vccd1 _0570_ sky130_fd_sc_hd__a21oi_1
XANTENNA__3218__CLK clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1566_ _0505_ _0513_ _0429_ vssd1 vssd1 vccd1 vccd1 _0514_ sky130_fd_sc_hd__mux2_1
XANTENNA__2541__A2 _1078_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3305_ clknet_leaf_33_clk uart_receiver.temp_byte\[5\] net160 vssd1 vssd1 vccd1 vccd1
+ buffer.Rx_byte\[5\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkload12_A clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1497_ _0437_ _0439_ _0444_ vssd1 vssd1 vccd1 vccd1 _0449_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_146_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3236_ clknet_leaf_13_clk _0210_ net198 vssd1 vssd1 vccd1 vccd1 host_message_reg.setLetter\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_6_Left_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3167_ clknet_leaf_30_clk _0143_ net184 vssd1 vssd1 vccd1 vccd1 hostdisp.top\[51\]
+ sky130_fd_sc_hd__dfrtp_1
X_2118_ hostdisp.curr_guesses\[1\] net120 _0861_ net136 vssd1 vssd1 vccd1 vccd1 hostdisp.nextBottom\[41\]
+ sky130_fd_sc_hd__o211a_1
X_3098_ clknet_leaf_27_clk _0088_ vssd1 vssd1 vccd1 vccd1 lcdPlayer.cnt_500hz\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_2049_ _0833_ vssd1 vssd1 vccd1 vccd1 _0834_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_65_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_178_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2057__B2 net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_18_clk_A clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout79 _0826_ vssd1 vssd1 vccd1 vccd1 net79 sky130_fd_sc_hd__buf_2
Xfanout68 net69 vssd1 vssd1 vccd1 vccd1 net68 sky130_fd_sc_hd__buf_2
Xfanout57 net59 vssd1 vssd1 vccd1 vccd1 net57 sky130_fd_sc_hd__buf_2
XFILLER_0_134_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_161_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_161_199 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_153_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2532__A2 net106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_164_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_169_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_169_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_157_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_123_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkload16 clknet_leaf_27_clk vssd1 vssd1 vccd1 vccd1 clkload16/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_82_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload27 clknet_leaf_15_clk vssd1 vssd1 vccd1 vccd1 clkload27/Y sky130_fd_sc_hd__inv_6
XTAP_TAPCELL_ROW_11_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1420_ keypadFSMPlayer.state\[0\] vssd1 vssd1 vccd1 vccd1 _0374_ sky130_fd_sc_hd__inv_2
XFILLER_0_50_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2523__A2 _1081_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3510__CLK clknet_leaf_31_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_79_Left_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_183_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3021_ clknet_leaf_9_clk net438 net217 vssd1 vssd1 vccd1 vccd1 clock_div.count\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_162_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2039__A1 net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_175_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_62_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_141_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_88_Left_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2805_ net142 gamelogic.setWord\[12\] vssd1 vssd1 vccd1 vccd1 _1351_ sky130_fd_sc_hd__nand2_1
XFILLER_0_73_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_193_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2736_ _0537_ _1288_ _0565_ vssd1 vssd1 vccd1 vccd1 _1290_ sky130_fd_sc_hd__o21ai_2
XANTENNA__2211__A1 net97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2667_ uart_transmitter.bit_index\[2\] _0665_ _0669_ vssd1 vssd1 vccd1 vccd1 _1234_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_14_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1618_ _0543_ _0552_ vssd1 vssd1 vccd1 vccd1 _0553_ sky130_fd_sc_hd__and2_1
XFILLER_0_1_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout214 net218 vssd1 vssd1 vccd1 vccd1 net214 sky130_fd_sc_hd__clkbuf_2
Xfanout203 net205 vssd1 vssd1 vccd1 vccd1 net203 sky130_fd_sc_hd__clkbuf_4
X_2598_ _1169_ _1170_ _1171_ net226 vssd1 vssd1 vccd1 vccd1 _1172_ sky130_fd_sc_hd__o31a_1
XPHY_EDGE_ROW_97_Left_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3190__CLK clknet_leaf_31_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2514__A2 net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1549_ _0372_ _0373_ _1401_ vssd1 vssd1 vccd1 vccd1 _0497_ sky130_fd_sc_hd__and3_1
XFILLER_0_5_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout225 net8 vssd1 vssd1 vccd1 vccd1 net225 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_2_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout180_X net180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3219_ clknet_leaf_2_clk _0195_ net172 vssd1 vssd1 vccd1 vccd1 gamelogic.indexCorrect\[2\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_166_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_166_269 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2450__A1 net130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_122 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2202__A1 net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3533__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_380 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_170_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold290 dispFSM.guesses\[20\] vssd1 vssd1 vccd1 vccd1 net554 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_46_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_189_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2269__A1 dispFSM.msg\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_16_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_258 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_173_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1467__A net4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3570_ net254 vssd1 vssd1 vccd1 vccd1 gpio_oeb[3] sky130_fd_sc_hd__buf_2
XFILLER_0_178_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2521_ hostdisp.top\[72\] _1095_ _1098_ hostdisp.top\[40\] vssd1 vssd1 vccd1 vccd1
+ _1099_ sky130_fd_sc_hd__a22o_1
XFILLER_0_11_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2452_ net130 host_message_reg.setLetter\[7\] hostdisp.curr_word\[23\] net73 net71
+ vssd1 vssd1 vccd1 vccd1 _1049_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_18_Right_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1403_ net273 vssd1 vssd1 vccd1 vccd1 _0357_ sky130_fd_sc_hd__inv_2
X_2383_ lcdPlayer.cnt_20ms\[14\] lcdPlayer.cnt_20ms\[13\] _1010_ vssd1 vssd1 vccd1
+ vccd1 _1014_ sky130_fd_sc_hd__and3_1
Xinput3 gpio_in[21] vssd1 vssd1 vccd1 vccd1 net3 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_143_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3004_ net211 vssd1 vssd1 vccd1 vccd1 _0029_ sky130_fd_sc_hd__inv_2
XFILLER_0_36_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3406__CLK clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_27_Right_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_22_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout140_A gamelogic.letter\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2983__A2 net53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3556__CLK clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2719_ net140 _0391_ _1279_ _1281_ vssd1 vssd1 vccd1 vccd1 _1282_ sky130_fd_sc_hd__a211o_1
XFILLER_0_14_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_36_Right_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_186_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_161_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout53_A _1393_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_45_Right_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_54_Right_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_189_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3429__CLK clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_63_Right_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_189_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1465__A2 net6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_307 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_145_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1952_ _0770_ _0185_ _0789_ _0186_ vssd1 vssd1 vccd1 vccd1 _0796_ sky130_fd_sc_hd__a31o_1
X_1883_ _0740_ _0741_ vssd1 vssd1 vccd1 vccd1 uart_transmitter.next_clk_count\[5\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_125_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_190_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_72_Right_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3553_ clknet_leaf_0_clk hostdisp.next_curr_guesses\[35\] net170 vssd1 vssd1 vccd1
+ vccd1 hostdisp.curr_guesses\[35\] sky130_fd_sc_hd__dfstp_1
X_3484_ clknet_leaf_31_clk hostdisp.next_curr_word\[6\] net164 vssd1 vssd1 vccd1 vccd1
+ hostdisp.curr_word\[6\] sky130_fd_sc_hd__dfstp_1
X_2504_ lcdPlayer.nextState\[3\] lcdPlayer.nextState\[2\] vssd1 vssd1 vccd1 vccd1
+ _1082_ sky130_fd_sc_hd__and2b_1
X_2435_ hostdisp.curr_word\[16\] net119 vssd1 vssd1 vccd1 vccd1 _1039_ sky130_fd_sc_hd__or2_1
XFILLER_0_11_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2366_ net443 _1000_ net167 vssd1 vssd1 vccd1 vccd1 _1003_ sky130_fd_sc_hd__o21ai_1
X_2297_ _0752_ _0955_ _0961_ vssd1 vssd1 vccd1 vccd1 _0087_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_81_Right_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_71 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_191_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout143_X net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_356 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2956__A2 net52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_90_Right_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_179_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2644__A1 net108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_186_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_182_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3101__CLK clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_90_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2220_ gamelogic.state\[1\] _0812_ vssd1 vssd1 vccd1 vccd1 _0916_ sky130_fd_sc_hd__or2_2
XFILLER_0_175_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2151_ gamelogic.setWord\[18\] hostdisp.curr_guesses\[18\] net122 vssd1 vssd1 vccd1
+ vccd1 _0878_ sky130_fd_sc_hd__mux2_1
X_2082_ hostdisp.curr_word\[20\] net103 _0845_ gamelogic.letter\[4\] vssd1 vssd1 vccd1
+ vccd1 hostdisp.next_curr_word\[20\] sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_49_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_191_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_187_Right_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_179_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2984_ gamelogic.setWord\[23\] net55 _1394_ gamelogic.setWord\[31\] vssd1 vssd1 vccd1
+ vccd1 _0347_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_32_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_239 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1935_ _0777_ _0782_ vssd1 vssd1 vccd1 vccd1 _0783_ sky130_fd_sc_hd__or2_1
XANTENNA__3405__SET_B net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1866_ keypadHostt.scan_col\[2\] net147 net230 vssd1 vssd1 vccd1 vccd1 net41 sky130_fd_sc_hd__mux2_1
XANTENNA__1610__A2 net3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_15_Left_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3605_ net239 vssd1 vssd1 vccd1 vccd1 gpio_out[5] sky130_fd_sc_hd__buf_2
X_1797_ net437 clock_div.count\[0\] vssd1 vssd1 vccd1 vccd1 clock_div.next_count\[1\]
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_140_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout103_A net104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3536_ clknet_leaf_2_clk hostdisp.next_curr_guesses\[18\] net176 vssd1 vssd1 vccd1
+ vccd1 hostdisp.curr_guesses\[18\] sky130_fd_sc_hd__dfstp_1
X_3467_ clknet_leaf_13_clk _0345_ net198 vssd1 vssd1 vccd1 vccd1 gamelogic.setWord\[29\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_149_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3398_ clknet_leaf_24_clk _0287_ net188 vssd1 vssd1 vccd1 vccd1 dispFSM.guesses\[52\]
+ sky130_fd_sc_hd__dfstp_1
X_2418_ hostdisp.curr_word\[4\] net72 net69 hostdisp.top\[44\] vssd1 vssd1 vccd1 vccd1
+ _0136_ sky130_fd_sc_hd__a22o_1
XANTENNA__2486__A net106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_24_Left_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2349_ lcdPlayer.cnt_20ms\[1\] lcdPlayer.cnt_20ms\[0\] vssd1 vssd1 vccd1 vccd1 _0993_
+ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_154_Right_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2626__A1 net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_0_Right_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_181_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_33_Left_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_156_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3274__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_42_Left_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2396__A _0017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_121_Right_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_262 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2617__A1 net226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_126_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_51_Left_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_182_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1720_ uart_receiver.clk_count\[10\] uart_receiver.clk_count\[2\] uart_receiver.clk_count\[3\]
+ uart_receiver.clk_count\[9\] vssd1 vssd1 vccd1 vccd1 _0636_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_79_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1651_ _0537_ _0564_ _0582_ _0585_ vssd1 vssd1 vccd1 vccd1 _0586_ sky130_fd_sc_hd__and4_1
Xhold108 clock_div.count\[8\] vssd1 vssd1 vccd1 vccd1 net372 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold119 hostdisp.top\[49\] vssd1 vssd1 vccd1 vccd1 net383 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_186_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1582_ _0509_ _0511_ vssd1 vssd1 vccd1 vccd1 _0527_ sky130_fd_sc_hd__xnor2_1
X_3321_ clknet_leaf_9_clk _0007_ net215 vssd1 vssd1 vccd1 vccd1 keypadFSMHost.state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2553__B1 _1097_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_192_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_60_Left_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3252_ clknet_leaf_3_clk hostdisp.nextBottom\[50\] net178 vssd1 vssd1 vccd1 vccd1
+ hostdisp.bottom\[50\] sky130_fd_sc_hd__dfrtp_1
X_2203_ net132 _0381_ vssd1 vssd1 vccd1 vccd1 _0904_ sky130_fd_sc_hd__nor2_1
X_3183_ clknet_leaf_30_clk _0159_ net181 vssd1 vssd1 vccd1 vccd1 hostdisp.top\[67\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_185_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2134_ gamelogic.setWord\[1\] _0869_ net136 vssd1 vssd1 vccd1 vccd1 hostdisp.nextBottom\[49\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2065_ hostdisp.curr_word\[8\] net102 _0840_ gamelogic.letter\[0\] vssd1 vssd1 vccd1
+ vccd1 hostdisp.next_curr_word\[8\] sky130_fd_sc_hd__o22a_1
XFILLER_0_146_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_158_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2967_ gamelogic.setWord\[6\] net53 net49 gamelogic.setWord\[14\] vssd1 vssd1 vccd1
+ vccd1 _0330_ sky130_fd_sc_hd__o22a_1
XFILLER_0_60_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout220_A net221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2898_ dispFSM.guesses\[38\] net85 net63 net556 vssd1 vssd1 vccd1 vccd1 _0265_ sky130_fd_sc_hd__o22a_1
XFILLER_0_97_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1918_ net166 _0769_ vssd1 vssd1 vccd1 vccd1 _0770_ sky130_fd_sc_hd__nand2_2
X_1849_ net355 _0723_ vssd1 vssd1 vccd1 vccd1 clock_div.next_count\[23\] sky130_fd_sc_hd__xor2_1
XFILLER_0_114_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2544__B1 net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout106_X net106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3519_ clknet_leaf_13_clk hostdisp.next_curr_guesses\[1\] net197 vssd1 vssd1 vccd1
+ vccd1 hostdisp.curr_guesses\[1\] sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_68_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2155__S net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_158_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_310 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_20_clk clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_20_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__1586__B2 dispFSM.msg\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2535__B1 _1106_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2471__C1 _1034_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_176_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2821_ net122 _0910_ _0929_ _0909_ vssd1 vssd1 vccd1 vccd1 _1362_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_11_clk clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_11_clk
+ sky130_fd_sc_hd__clkbuf_8
X_2752_ _0557_ _0547_ _0543_ net153 vssd1 vssd1 vccd1 vccd1 _1306_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_143_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1577__B2 dispFSM.msg\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1703_ _0396_ _0617_ vssd1 vssd1 vccd1 vccd1 _0619_ sky130_fd_sc_hd__or2_1
XFILLER_0_41_324 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2683_ _0923_ net66 _1248_ vssd1 vssd1 vccd1 vccd1 _1249_ sky130_fd_sc_hd__a21oi_1
X_1634_ net151 keypadFSMHost.prev_key\[2\] _0546_ vssd1 vssd1 vccd1 vccd1 _0569_ sky130_fd_sc_hd__and3_1
XFILLER_0_111_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1565_ net233 _0435_ _0467_ _0506_ vssd1 vssd1 vccd1 vccd1 _0513_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_111_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3304_ clknet_leaf_33_clk uart_receiver.temp_byte\[4\] net160 vssd1 vssd1 vccd1 vccd1
+ buffer.Rx_byte\[4\] sky130_fd_sc_hd__dfrtp_1
X_3235_ clknet_leaf_15_clk _0209_ net215 vssd1 vssd1 vccd1 vccd1 host_message_reg.setLetter\[4\]
+ sky130_fd_sc_hd__dfstp_2
X_1496_ _0439_ _0447_ vssd1 vssd1 vccd1 vccd1 _0448_ sky130_fd_sc_hd__nor2_1
XFILLER_0_39_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_146_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3166_ clknet_leaf_3_clk _0142_ net178 vssd1 vssd1 vccd1 vccd1 hostdisp.top\[50\]
+ sky130_fd_sc_hd__dfrtp_1
X_2117_ gamelogic.setWord\[1\] net125 vssd1 vssd1 vccd1 vccd1 _0861_ sky130_fd_sc_hd__or2_1
X_3097_ clknet_leaf_27_clk _0087_ vssd1 vssd1 vccd1 vccd1 lcdPlayer.cnt_500hz\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_105_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2057__A2 net96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2048_ _0405_ net98 net75 _0832_ gamelogic.indexCorrect\[0\] vssd1 vssd1 vccd1 vccd1
+ _0833_ sky130_fd_sc_hd__o2111a_1
XTAP_TAPCELL_ROW_65_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout47 net48 vssd1 vssd1 vccd1 vccd1 net47 sky130_fd_sc_hd__clkbuf_4
Xfanout58 net59 vssd1 vssd1 vccd1 vccd1 net58 sky130_fd_sc_hd__buf_2
XFILLER_0_29_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout69 net71 vssd1 vssd1 vccd1 vccd1 net69 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout223_X net223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_134 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_107_Left_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3312__CLK clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_164_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_116_Left_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3462__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_192_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2613__S net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_22_clk_X clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload17 clknet_leaf_28_clk vssd1 vssd1 vccd1 vccd1 clkload17/Y sky130_fd_sc_hd__inv_6
Xclkload28 clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 clkload28/Y sky130_fd_sc_hd__clkinv_8
XFILLER_0_140_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3020_ clknet_leaf_9_clk clock_div.next_count\[0\] net217 vssd1 vssd1 vccd1 vccd1
+ clock_div.count\[0\] sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_0_clk clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_0_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_155_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2039__A2 net95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_141_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_183_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2804_ net142 gamelogic.setWord\[12\] vssd1 vssd1 vccd1 vccd1 _1350_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_193_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2735_ _0537_ _1288_ vssd1 vssd1 vccd1 vccd1 _1289_ sky130_fd_sc_hd__nor2_1
XFILLER_0_26_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2666_ uart_transmitter.bit_index\[1\] _1232_ _0669_ _0666_ vssd1 vssd1 vccd1 vccd1
+ _0191_ sky130_fd_sc_hd__o211a_1
X_1617_ keypadHostt.scan_col\[0\] net153 keypadHostt.scan_col\[3\] net151 vssd1 vssd1
+ vccd1 vccd1 _0552_ sky130_fd_sc_hd__or4_4
Xfanout204 net205 vssd1 vssd1 vccd1 vccd1 net204 sky130_fd_sc_hd__clkbuf_4
X_2597_ dispFSM.guesses\[68\] _1072_ net113 dispFSM.guesses\[52\] _1167_ vssd1 vssd1
+ vccd1 vccd1 _1171_ sky130_fd_sc_hd__a221o_1
XFILLER_0_1_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1548_ _0471_ _0495_ _0490_ vssd1 vssd1 vccd1 vccd1 _0496_ sky130_fd_sc_hd__nor3b_2
XFILLER_0_157_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout215 net218 vssd1 vssd1 vccd1 vccd1 net215 sky130_fd_sc_hd__clkbuf_4
Xfanout226 net228 vssd1 vssd1 vccd1 vccd1 net226 sky130_fd_sc_hd__clkbuf_4
X_1479_ _0429_ _0430_ _0422_ vssd1 vssd1 vccd1 vccd1 _0431_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_2_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3218_ clknet_leaf_3_clk _0194_ net172 vssd1 vssd1 vccd1 vccd1 gamelogic.indexCorrect\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_3149_ clknet_leaf_26_clk _0125_ vssd1 vssd1 vccd1 vccd1 lcdPlayer.cnt_20ms\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2986__B1 net49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2450__A2 host_message_reg.setLetter\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2669__A net96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold280 hostdisp.curr_guesses\[19\] vssd1 vssd1 vccd1 vccd1 net544 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold291 dispFSM.guesses\[43\] vssd1 vssd1 vccd1 vccd1 net555 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_189_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_86_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3208__CLK clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2977__B1 net49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_165_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2441__A2 net67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1467__B net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3358__CLK clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2520_ lcdPlayer.nextState\[2\] _1060_ _1062_ vssd1 vssd1 vccd1 vccd1 _1098_ sky130_fd_sc_hd__nor3_4
X_2451_ net341 net67 _1048_ vssd1 vssd1 vccd1 vccd1 _0154_ sky130_fd_sc_hd__o21a_1
XFILLER_0_11_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1507__A_N dispFSM.msg\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1402_ net139 vssd1 vssd1 vccd1 vccd1 _0356_ sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_17_clk_A clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2298__B _0752_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2382_ _1013_ net168 _1012_ vssd1 vssd1 vccd1 vccd1 _0120_ sky130_fd_sc_hd__and3b_1
XFILLER_0_46_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput4 gpio_in[22] vssd1 vssd1 vccd1 vccd1 net4 sky130_fd_sc_hd__clkbuf_2
X_3003_ net211 vssd1 vssd1 vccd1 vccd1 _0028_ sky130_fd_sc_hd__inv_2
Xclkbuf_2_1__f_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_2_1__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_148_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_143_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_102_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout133_A hostdisp.Cstate vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2718_ _0378_ gamelogic.setWord\[1\] gamelogic.setWord\[2\] _0379_ _1280_ vssd1 vssd1
+ vccd1 vccd1 _1281_ sky130_fd_sc_hd__a221o_1
XFILLER_0_14_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2649_ hostdisp.bottom\[79\] net112 net109 hostdisp.bottom\[63\] _1218_ vssd1 vssd1
+ vccd1 vccd1 _1220_ sky130_fd_sc_hd__a221o_1
XANTENNA__2499__A2 _1072_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_161_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2952__A net97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2959__B1 net49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2163__S net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2671__B net144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3500__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2423__A2 _0830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_352 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_168_Right_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3291__Q host_message_reg.Cstate vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkload9_A clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2111__B2 net140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3180__CLK clknet_leaf_31_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_207 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1951_ _0185_ _0794_ vssd1 vssd1 vccd1 vccd1 _0795_ sky130_fd_sc_hd__nor2_1
X_1882_ net523 _0739_ _0732_ vssd1 vssd1 vccd1 vccd1 _0741_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_22_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3621_ net249 vssd1 vssd1 vccd1 vccd1 gpio_out[33] sky130_fd_sc_hd__buf_2
XFILLER_0_189_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_58 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3552_ clknet_leaf_0_clk hostdisp.next_curr_guesses\[34\] net175 vssd1 vssd1 vccd1
+ vccd1 hostdisp.curr_guesses\[34\] sky130_fd_sc_hd__dfstp_1
XFILLER_0_11_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_260 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2503_ net138 net139 _1075_ vssd1 vssd1 vccd1 vccd1 _1081_ sky130_fd_sc_hd__and3_2
XFILLER_0_51_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3483_ clknet_leaf_28_clk hostdisp.next_curr_word\[5\] net166 vssd1 vssd1 vccd1 vccd1
+ hostdisp.curr_word\[5\] sky130_fd_sc_hd__dfrtp_1
X_2434_ hostdisp.curr_word\[15\] net73 net70 net347 vssd1 vssd1 vccd1 vccd1 _0147_
+ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_135_Right_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2365_ lcdPlayer.cnt_20ms\[8\] lcdPlayer.cnt_20ms\[7\] _0998_ vssd1 vssd1 vccd1 vccd1
+ _1002_ sky130_fd_sc_hd__and3_1
X_2296_ lcdPlayer.cnt_500hz\[4\] _0751_ vssd1 vssd1 vccd1 vccd1 _0961_ sky130_fd_sc_hd__or2_1
XFILLER_0_2_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2653__A2 net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_176_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_138 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout136_X net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_368 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_179_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3588__260 vssd1 vssd1 vccd1 vccd1 net260 _3588__260/LO sky130_fd_sc_hd__conb_1
XFILLER_0_2_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_102_Right_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2158__S net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout49_X net49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_190 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2621__S net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2150_ gamelogic.setWord\[9\] _0877_ net135 vssd1 vssd1 vccd1 vccd1 hostdisp.nextBottom\[57\]
+ sky130_fd_sc_hd__mux2_1
X_3604__238 vssd1 vssd1 vccd1 vccd1 _3604__238/HI net238 sky130_fd_sc_hd__conb_1
X_2081_ hostdisp.curr_word\[19\] net103 _0845_ gamelogic.letter\[3\] vssd1 vssd1 vccd1
+ vccd1 hostdisp.next_curr_word\[19\] sky130_fd_sc_hd__o22a_1
XFILLER_0_191_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2635__A2 net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_179_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2983_ gamelogic.setWord\[22\] net53 net49 gamelogic.setWord\[30\] vssd1 vssd1 vccd1
+ vccd1 _0346_ sky130_fd_sc_hd__o22a_1
XFILLER_0_118_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_32_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_173_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1934_ _0185_ _0776_ vssd1 vssd1 vccd1 vccd1 _0782_ sky130_fd_sc_hd__and2_1
X_1865_ net152 keypadplayer.scan_col\[1\] net230 vssd1 vssd1 vccd1 vccd1 net40 sky130_fd_sc_hd__mux2_1
XFILLER_0_140_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3604_ net238 vssd1 vssd1 vccd1 vccd1 gpio_out[4] sky130_fd_sc_hd__buf_2
X_1796_ clock_div.count\[0\] _0693_ vssd1 vssd1 vccd1 vccd1 clock_div.next_count\[0\]
+ sky130_fd_sc_hd__and2b_1
X_3535_ clknet_leaf_5_clk hostdisp.next_curr_guesses\[17\] net200 vssd1 vssd1 vccd1
+ vccd1 hostdisp.curr_guesses\[17\] sky130_fd_sc_hd__dfstp_1
XFILLER_0_141_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3466_ clknet_leaf_6_clk _0344_ net192 vssd1 vssd1 vccd1 vccd1 gamelogic.setWord\[28\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_58_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2417_ hostdisp.curr_word\[3\] net72 net69 net447 vssd1 vssd1 vccd1 vccd1 _0135_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3397_ clknet_leaf_25_clk _0286_ net184 vssd1 vssd1 vccd1 vccd1 dispFSM.guesses\[51\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_149_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2348_ net520 _0017_ _0955_ vssd1 vssd1 vccd1 vccd1 _0107_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_165_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2279_ _0358_ _0947_ vssd1 vssd1 vccd1 vccd1 _0948_ sky130_fd_sc_hd__nor2_1
XFILLER_0_168_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_207 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2011__B1 net79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2562__A1 dispFSM.msg\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_167_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_187_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_126_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_155_313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_240 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1650_ keypadFSMHost.state\[5\] _0583_ _0584_ vssd1 vssd1 vccd1 vccd1 _0585_ sky130_fd_sc_hd__and3_1
X_1581_ _0519_ _0524_ _0526_ _0454_ dispFSM.msg\[2\] vssd1 vssd1 vccd1 vccd1 _0060_
+ sky130_fd_sc_hd__o32a_1
XFILLER_0_123_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold109 dispFSM.guesses\[45\] vssd1 vssd1 vccd1 vccd1 net373 sky130_fd_sc_hd__dlygate4sd3_1
X_3320_ clknet_leaf_10_clk _0006_ net215 vssd1 vssd1 vccd1 vccd1 keypadFSMHost.state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3251_ clknet_leaf_13_clk hostdisp.nextBottom\[49\] net198 vssd1 vssd1 vccd1 vccd1
+ hostdisp.bottom\[49\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_185_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3182_ clknet_leaf_31_clk _0158_ net174 vssd1 vssd1 vccd1 vccd1 hostdisp.top\[66\]
+ sky130_fd_sc_hd__dfrtp_1
X_2202_ net129 gamelogic.setWord\[35\] _0903_ vssd1 vssd1 vccd1 vccd1 hostdisp.nextBottom\[83\]
+ sky130_fd_sc_hd__a21o_1
X_2133_ gamelogic.setWord\[9\] hostdisp.curr_guesses\[9\] net125 vssd1 vssd1 vccd1
+ vccd1 _0869_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2608__A2 _1086_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2064_ _0840_ vssd1 vssd1 vccd1 vccd1 _0841_ sky130_fd_sc_hd__inv_2
XFILLER_0_48_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2966_ net566 net55 _1394_ net552 vssd1 vssd1 vccd1 vccd1 _0329_ sky130_fd_sc_hd__a22o_1
XFILLER_0_29_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2897_ dispFSM.guesses\[37\] net90 net64 net434 vssd1 vssd1 vccd1 vccd1 _0264_ sky130_fd_sc_hd__a22o_1
X_1917_ lcdPlayer.nextState\[2\] lcdPlayer.currentState\[2\] _0764_ vssd1 vssd1 vccd1
+ vccd1 _0769_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_390 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout213_A net218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1848_ _0722_ _0723_ vssd1 vssd1 vccd1 vccd1 clock_div.next_count\[22\] sky130_fd_sc_hd__nor2_1
XFILLER_0_8_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1779_ message_reg.msg\[6\] message_reg.msg\[7\] uart_transmitter.bit_index\[0\]
+ vssd1 vssd1 vccd1 vccd1 _0678_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3518_ clknet_leaf_5_clk hostdisp.next_curr_guesses\[0\] net199 vssd1 vssd1 vccd1
+ vccd1 hostdisp.curr_guesses\[0\] sky130_fd_sc_hd__dfstp_1
X_3449_ clknet_leaf_4_clk _0327_ net177 vssd1 vssd1 vccd1 vccd1 gamelogic.setWord\[11\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_176_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_169_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_68_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_211 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_322 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_176 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2783__A1 host_message_reg.setLetter\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2171__S net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3391__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2694__X _1259_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_155_143 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2820_ _0670_ _0672_ message_reg.state\[0\] _0370_ vssd1 vssd1 vccd1 vccd1 _0217_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_85_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2751_ _1304_ vssd1 vssd1 vccd1 vccd1 _1305_ sky130_fd_sc_hd__inv_2
XFILLER_0_143_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1702_ _0396_ _0617_ vssd1 vssd1 vccd1 vccd1 _0618_ sky130_fd_sc_hd__nor2_2
X_2682_ _1242_ _1247_ _0924_ vssd1 vssd1 vccd1 vccd1 _1248_ sky130_fd_sc_hd__a21oi_1
X_1633_ net152 _0546_ keypadFSMHost.prev_key\[1\] vssd1 vssd1 vccd1 vccd1 _0568_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_151_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_187_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1564_ _0509_ _0510_ _0504_ vssd1 vssd1 vccd1 vccd1 _0512_ sky130_fd_sc_hd__a21o_1
XFILLER_0_111_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1495_ _0442_ _0444_ vssd1 vssd1 vccd1 vccd1 _0447_ sky130_fd_sc_hd__or2_1
XFILLER_0_39_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3303_ clknet_leaf_34_clk uart_receiver.temp_byte\[3\] net159 vssd1 vssd1 vccd1 vccd1
+ buffer.Rx_byte\[3\] sky130_fd_sc_hd__dfrtp_1
X_3234_ clknet_leaf_12_clk _0208_ net221 vssd1 vssd1 vccd1 vccd1 host_message_reg.setLetter\[3\]
+ sky130_fd_sc_hd__dfstp_2
XTAP_TAPCELL_ROW_146_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3165_ clknet_leaf_30_clk _0141_ net185 vssd1 vssd1 vccd1 vccd1 hostdisp.top\[49\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_146_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2116_ hostdisp.curr_guesses\[0\] net120 _0860_ net135 vssd1 vssd1 vccd1 vccd1 hostdisp.nextBottom\[40\]
+ sky130_fd_sc_hd__o211a_1
X_3096_ clknet_leaf_27_clk _0086_ vssd1 vssd1 vccd1 vccd1 lcdPlayer.cnt_500hz\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__3264__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout163_A net164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2047_ hostdisp.curr_word\[1\] hostdisp.curr_word\[2\] hostdisp.curr_word\[3\] _0404_
+ net98 vssd1 vssd1 vccd1 vccd1 _0832_ sky130_fd_sc_hd__a41o_1
XTAP_TAPCELL_ROW_65_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_105_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_162_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout48 net50 vssd1 vssd1 vccd1 vccd1 net48 sky130_fd_sc_hd__buf_2
Xfanout59 _1391_ vssd1 vssd1 vccd1 vccd1 net59 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_161_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2949_ host_message_reg.Cstate keypadFSMHost.state\[4\] keypadFSMHost.state\[0\]
+ _0595_ vssd1 vssd1 vccd1 vccd1 _1392_ sky130_fd_sc_hd__nor4_1
XFILLER_0_29_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_146 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2498__Y _1076_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_187_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout76_A net77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_164_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_169_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2690__A gamelogic.letter\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload29 clknet_leaf_17_clk vssd1 vssd1 vccd1 vccd1 clkload29/Y sky130_fd_sc_hd__inv_12
XFILLER_0_152_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload18 clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 clkload18/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_133_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3287__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2692__B1 gamelogic.setWord\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3383__RESET_B net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_141_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3469__Q gamelogic.setWord\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3530__SET_B net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2803_ gamelogic.letter\[3\] gamelogic.setWord\[11\] vssd1 vssd1 vccd1 vccd1 _1349_
+ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_70_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_193_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_183_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2734_ _0602_ keypadFSMHost.state\[4\] keypadFSMHost.state\[0\] vssd1 vssd1 vccd1
+ vccd1 _1288_ sky130_fd_sc_hd__or3b_2
X_2665_ _1232_ _1233_ vssd1 vssd1 vccd1 vccd1 _0190_ sky130_fd_sc_hd__nor2_1
X_1616_ net153 _0547_ vssd1 vssd1 vccd1 vccd1 _0551_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_152_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2596_ dispFSM.guesses\[76\] _1086_ _1142_ vssd1 vssd1 vccd1 vccd1 _1170_ sky130_fd_sc_hd__a21o_1
Xfanout205 net206 vssd1 vssd1 vccd1 vccd1 net205 sky130_fd_sc_hd__buf_2
Xfanout216 net217 vssd1 vssd1 vccd1 vccd1 net216 sky130_fd_sc_hd__clkbuf_4
X_1547_ _0371_ _0492_ _0494_ keypadFSMPlayer.state\[3\] vssd1 vssd1 vccd1 vccd1 _0495_
+ sky130_fd_sc_hd__a31oi_2
Xfanout227 net228 vssd1 vssd1 vccd1 vccd1 net227 sky130_fd_sc_hd__clkbuf_4
X_1478_ keypadplayer.scan_col\[1\] keypadplayer.scan_col\[0\] net147 vssd1 vssd1 vccd1
+ vccd1 _0430_ sky130_fd_sc_hd__or3_4
XTAP_TAPCELL_ROW_2_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3217_ clknet_leaf_31_clk _0193_ net164 vssd1 vssd1 vccd1 vccd1 gamelogic.indexCorrect\[4\]
+ sky130_fd_sc_hd__dfrtp_2
X_3148_ clknet_leaf_25_clk _0124_ vssd1 vssd1 vccd1 vccd1 lcdPlayer.cnt_20ms\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_173_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_173_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3079_ clknet_leaf_33_clk net301 net161 vssd1 vssd1 vccd1 vccd1 buffer.temp_guess\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_280 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_149_Right_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold270 gamelogic.setWord\[5\] vssd1 vssd1 vccd1 vccd1 net534 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold292 dispFSM.guesses\[30\] vssd1 vssd1 vccd1 vccd1 net556 sky130_fd_sc_hd__dlygate4sd3_1
Xhold281 hostdisp.curr_guesses\[44\] vssd1 vssd1 vccd1 vccd1 net545 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout79_X net79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_116_Right_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_132_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2450_ net130 host_message_reg.setLetter\[6\] _0828_ _1047_ net71 vssd1 vssd1 vccd1
+ vccd1 _1048_ sky130_fd_sc_hd__a221o_1
XFILLER_0_11_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2381_ lcdPlayer.cnt_20ms\[13\] _1009_ vssd1 vssd1 vccd1 vccd1 _1013_ sky130_fd_sc_hd__and2_1
Xinput5 gpio_in[23] vssd1 vssd1 vccd1 vccd1 net5 sky130_fd_sc_hd__clkbuf_1
X_3002_ net208 vssd1 vssd1 vccd1 vccd1 _0027_ sky130_fd_sc_hd__inv_2
XFILLER_0_127_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_135_Left_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_102_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2417__B1 net69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1939__A _0017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3302__CLK clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2717_ _0382_ gamelogic.setWord\[4\] gamelogic.setWord\[7\] _0386_ vssd1 vssd1 vccd1
+ vccd1 _1280_ sky130_fd_sc_hd__a22o_1
XFILLER_0_14_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3452__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_144_Left_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2648_ hostdisp.bottom\[71\] _1085_ net108 hostdisp.top\[63\] vssd1 vssd1 vccd1 vccd1
+ _1219_ sky130_fd_sc_hd__a22o_1
XFILLER_0_168_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2579_ hostdisp.top\[59\] dispFSM.msg\[3\] net226 vssd1 vssd1 vccd1 vccd1 _1154_
+ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_21_clk_X clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_184_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_161_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2656__B1 _1084_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2120__A2 net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_153_Left_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_114 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2959__A1 host_message_reg.setLetter\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_172_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_162_Left_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2619__S net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_189_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_171_Left_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2647__B1 _1095_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2111__A2 net96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_136 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3325__CLK clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_350 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_145_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1950_ _0771_ _0182_ vssd1 vssd1 vccd1 vccd1 _0794_ sky130_fd_sc_hd__nor2_1
XFILLER_0_83_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1881_ uart_transmitter.clk_count\[4\] uart_transmitter.clk_count\[5\] _0736_ vssd1
+ vssd1 vccd1 vccd1 _0740_ sky130_fd_sc_hd__and3_1
XFILLER_0_113_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_189_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3475__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3620_ lcdPlayer.lcd_en vssd1 vssd1 vccd1 vccd1 net38 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_180_Left_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3551_ clknet_leaf_7_clk hostdisp.next_curr_guesses\[33\] net196 vssd1 vssd1 vccd1
+ vccd1 hostdisp.curr_guesses\[33\] sky130_fd_sc_hd__dfstp_1
XFILLER_0_113_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1925__A2 _0764_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2502_ _1071_ _1073_ vssd1 vssd1 vccd1 vccd1 _1080_ sky130_fd_sc_hd__nor2_1
XFILLER_0_11_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3482_ clknet_leaf_32_clk hostdisp.next_curr_word\[4\] net164 vssd1 vssd1 vccd1 vccd1
+ hostdisp.curr_word\[4\] sky130_fd_sc_hd__dfstp_1
XFILLER_0_11_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2433_ net329 net68 _1038_ _0828_ vssd1 vssd1 vccd1 vccd1 _0146_ sky130_fd_sc_hd__a22o_1
XANTENNA__1689__A1 keypadFSMHost.state\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2364_ _1000_ _1001_ vssd1 vssd1 vccd1 vccd1 _0114_ sky130_fd_sc_hd__nor2_1
XANTENNA__2529__S net226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2295_ _0751_ _0955_ _0960_ vssd1 vssd1 vccd1 vccd1 _0086_ sky130_fd_sc_hd__and3b_1
XANTENNA__2638__B1 _1098_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_40 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_176_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout129_X net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input3_X net3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2439__S net67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3415__RESET_B net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3348__CLK clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2174__S net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3498__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_2_0__f_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_16_clk_A clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2203__A net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3497__SET_B net179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2080_ hostdisp.curr_word\[18\] net103 _0845_ gamelogic.letter\[2\] vssd1 vssd1 vccd1
+ vccd1 hostdisp.next_curr_word\[18\] sky130_fd_sc_hd__o22a_1
XFILLER_0_17_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2096__B2 net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2982_ gamelogic.setWord\[21\] net55 _1394_ gamelogic.setWord\[29\] vssd1 vssd1 vccd1
+ vccd1 _0345_ sky130_fd_sc_hd__a22o_1
XFILLER_0_130_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3477__Q gamelogic.setWord\[39\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1933_ _0766_ _0771_ _0780_ vssd1 vssd1 vccd1 vccd1 _0781_ sky130_fd_sc_hd__o21a_1
XFILLER_0_140_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3603_ net237 vssd1 vssd1 vccd1 vccd1 gpio_out[3] sky130_fd_sc_hd__buf_2
X_1864_ keypadHostt.scan_col\[0\] keypadplayer.scan_col\[0\] net230 vssd1 vssd1 vccd1
+ vccd1 net39 sky130_fd_sc_hd__mux2_1
XFILLER_0_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1795_ _0687_ _0692_ vssd1 vssd1 vccd1 vccd1 _0693_ sky130_fd_sc_hd__or2_4
XTAP_TAPCELL_ROW_99_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3534_ clknet_leaf_6_clk hostdisp.next_curr_guesses\[16\] net196 vssd1 vssd1 vccd1
+ vccd1 hostdisp.curr_guesses\[16\] sky130_fd_sc_hd__dfstp_1
XANTENNA__2113__A _0827_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3465_ clknet_leaf_1_clk _0343_ net176 vssd1 vssd1 vccd1 vccd1 gamelogic.setWord\[27\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__2571__A2 net105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2416_ hostdisp.curr_word\[2\] net72 net69 net559 vssd1 vssd1 vccd1 vccd1 _0134_
+ sky130_fd_sc_hd__a22o_1
X_3396_ clknet_leaf_24_clk _0285_ net189 vssd1 vssd1 vccd1 vccd1 dispFSM.guesses\[50\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_149_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2347_ uart_receiver.bit_index\[2\] _0992_ _0624_ vssd1 vssd1 vccd1 vccd1 _0106_
+ sky130_fd_sc_hd__o21a_1
X_2278_ lcdPlayer.cnt_20ms\[4\] _0945_ vssd1 vssd1 vccd1 vccd1 _0947_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_50 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_181_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_176_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_191_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2547__C1 _0752_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3170__CLK clknet_leaf_30_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_167_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2078__B2 net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_182_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_155_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_170_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1580_ _0437_ _0525_ _0448_ vssd1 vssd1 vccd1 vccd1 _0526_ sky130_fd_sc_hd__o21a_1
XFILLER_0_111_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3513__CLK clknet_leaf_31_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2553__A2 net105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_186_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3250_ clknet_leaf_5_clk hostdisp.nextBottom\[48\] net199 vssd1 vssd1 vccd1 vccd1
+ hostdisp.bottom\[48\] sky130_fd_sc_hd__dfrtp_1
X_3181_ clknet_leaf_30_clk _0157_ net177 vssd1 vssd1 vccd1 vccd1 hostdisp.top\[65\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_28_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2201_ net131 hostdisp.curr_guesses\[43\] net121 vssd1 vssd1 vccd1 vccd1 _0903_ sky130_fd_sc_hd__and3_1
XFILLER_0_178_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2132_ gamelogic.setWord\[0\] _0868_ net135 vssd1 vssd1 vccd1 vccd1 hostdisp.nextBottom\[48\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2069__B2 net142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2063_ _0837_ _0839_ vssd1 vssd1 vccd1 vccd1 _0840_ sky130_fd_sc_hd__nand2_2
XFILLER_0_135_88 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_158_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_173_100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3043__CLK clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2965_ gamelogic.setWord\[4\] net51 net47 gamelogic.setWord\[12\] vssd1 vssd1 vccd1
+ vccd1 _0328_ sky130_fd_sc_hd__o22a_1
XFILLER_0_60_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_200 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2896_ dispFSM.guesses\[36\] net85 net60 net507 vssd1 vssd1 vccd1 vccd1 _0263_ sky130_fd_sc_hd__o22a_1
X_1916_ _0768_ vssd1 vssd1 vccd1 vccd1 _0183_ sky130_fd_sc_hd__inv_2
X_1847_ clock_div.count\[21\] clock_div.count\[20\] clock_div.count\[22\] _0719_ vssd1
+ vssd1 vccd1 vccd1 _0723_ sky130_fd_sc_hd__and4_1
XFILLER_0_44_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_155_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_255 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout206_A net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1778_ message_reg.msg\[4\] message_reg.msg\[5\] uart_transmitter.bit_index\[0\]
+ vssd1 vssd1 vccd1 vccd1 _0677_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3517_ clknet_leaf_29_clk hostdisp.next_curr_word\[39\] net169 vssd1 vssd1 vccd1
+ vccd1 hostdisp.curr_word\[39\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3193__CLK clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3448_ clknet_leaf_3_clk _0326_ net175 vssd1 vssd1 vccd1 vccd1 gamelogic.setWord\[10\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__3480__SET_B net164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3379_ clknet_leaf_21_clk _0268_ net210 vssd1 vssd1 vccd1 vccd1 dispFSM.guesses\[33\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_68_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_192_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_223 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_51_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3536__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2535__A2 net105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_236 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_155 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2750_ _0557_ _1303_ vssd1 vssd1 vccd1 vccd1 _1304_ sky130_fd_sc_hd__nand2_1
XFILLER_0_26_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2681_ _1243_ _1244_ _1246_ vssd1 vssd1 vccd1 vccd1 _1247_ sky130_fd_sc_hd__and3b_1
XFILLER_0_26_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1701_ uart_receiver.state\[2\] uart_receiver.state\[1\] vssd1 vssd1 vccd1 vccd1
+ _0617_ sky130_fd_sc_hd__nand2b_1
X_1632_ keypadFSMHost.prev_key\[6\] _0557_ vssd1 vssd1 vccd1 vccd1 _0567_ sky130_fd_sc_hd__xor2_1
XFILLER_0_30_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_187_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1563_ _0504_ _0510_ vssd1 vssd1 vccd1 vccd1 _0511_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_39_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1494_ _0426_ _0430_ vssd1 vssd1 vccd1 vccd1 _0446_ sky130_fd_sc_hd__or2_1
X_3302_ clknet_leaf_33_clk uart_receiver.temp_byte\[2\] net159 vssd1 vssd1 vccd1 vccd1
+ buffer.Rx_byte\[2\] sky130_fd_sc_hd__dfrtp_1
X_3233_ clknet_leaf_12_clk _0207_ net197 vssd1 vssd1 vccd1 vccd1 host_message_reg.setLetter\[2\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_146_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3164_ clknet_leaf_4_clk _0140_ net177 vssd1 vssd1 vccd1 vccd1 hostdisp.top\[48\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__3409__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2115_ _0390_ net120 vssd1 vssd1 vccd1 vccd1 _0860_ sky130_fd_sc_hd__nand2_1
X_3095_ clknet_leaf_27_clk _0085_ vssd1 vssd1 vccd1 vccd1 lcdPlayer.cnt_500hz\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_2046_ hostdisp.curr_word\[4\] hostdisp.curr_word\[6\] net98 vssd1 vssd1 vccd1 vccd1
+ _0831_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_65_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3559__CLK clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout49 net50 vssd1 vssd1 vccd1 vccd1 net49 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_29_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2948_ _0186_ _0794_ _0795_ _0187_ vssd1 vssd1 vccd1 vccd1 _0315_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_161_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_199 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_161_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout111_X net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2879_ dispFSM.guesses\[19\] net82 net57 net509 vssd1 vssd1 vccd1 vccd1 _0246_ sky130_fd_sc_hd__o22a_1
XFILLER_0_142_372 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout69_A net71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_164_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_192_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_192_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_180_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_175_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_158 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload19 clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 clkload19/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_23_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_39_Left_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_48_Left_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_141_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_183_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2802_ net143 gamelogic.setWord\[11\] vssd1 vssd1 vccd1 vccd1 _1348_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_70_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_193_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2733_ net398 net6 _1287_ vssd1 vssd1 vccd1 vccd1 _0204_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1955__B1 _0607_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_57_Left_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2664_ _0664_ _0669_ uart_transmitter.bit_index\[0\] vssd1 vssd1 vccd1 vccd1 _1233_
+ sky130_fd_sc_hd__a21oi_1
X_1615_ net152 _0547_ vssd1 vssd1 vccd1 vccd1 _0550_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_152_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2595_ dispFSM.guesses\[60\] net117 net108 dispFSM.msg\[4\] _1168_ vssd1 vssd1 vccd1
+ vccd1 _1169_ sky130_fd_sc_hd__a221o_1
X_1546_ keypadFSMPlayer.state\[5\] _0493_ vssd1 vssd1 vccd1 vccd1 _0494_ sky130_fd_sc_hd__or2_1
Xfanout217 net218 vssd1 vssd1 vccd1 vccd1 net217 sky130_fd_sc_hd__clkbuf_4
Xfanout206 net224 vssd1 vssd1 vccd1 vccd1 net206 sky130_fd_sc_hd__clkbuf_2
Xfanout228 net7 vssd1 vssd1 vccd1 vccd1 net228 sky130_fd_sc_hd__clkbuf_4
X_1477_ net231 net6 net155 net128 vssd1 vssd1 vccd1 vccd1 _0429_ sky130_fd_sc_hd__nand4_4
X_3216_ clknet_leaf_18_clk _0192_ net219 vssd1 vssd1 vccd1 vccd1 uart_transmitter.bit_index\[2\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_2_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_66_Left_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3147_ clknet_leaf_25_clk _0123_ vssd1 vssd1 vccd1 vccd1 lcdPlayer.cnt_20ms\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_82_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3078_ clknet_leaf_35_clk net327 net161 vssd1 vssd1 vccd1 vccd1 buffer.temp_guess\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_166_217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2029_ hostdisp.curr_guesses\[43\] net91 net76 net542 vssd1 vssd1 vccd1 vccd1 hostdisp.next_curr_guesses\[35\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_49_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3022__RESET_B net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold260 dispFSM.guesses\[68\] vssd1 vssd1 vccd1 vccd1 net524 sky130_fd_sc_hd__dlygate4sd3_1
Xhold271 uart_receiver.clk_count\[10\] vssd1 vssd1 vccd1 vccd1 net535 sky130_fd_sc_hd__dlygate4sd3_1
Xhold293 dispFSM.guesses\[35\] vssd1 vssd1 vccd1 vccd1 net557 sky130_fd_sc_hd__dlygate4sd3_1
Xhold282 dispFSM.guesses\[24\] vssd1 vssd1 vccd1 vccd1 net546 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2177__S net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_178 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_84_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2977__A2 net53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_180_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3254__CLK clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2380_ lcdPlayer.cnt_20ms\[13\] _1009_ vssd1 vssd1 vccd1 vccd1 _1012_ sky130_fd_sc_hd__or2_1
Xinput6 gpio_in[24] vssd1 vssd1 vccd1 vccd1 net6 sky130_fd_sc_hd__clkbuf_4
X_3001_ net221 vssd1 vssd1 vccd1 vccd1 _0026_ sky130_fd_sc_hd__inv_2
XFILLER_0_160_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_148_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3533__RESET_B net206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2716_ gamelogic.letter\[0\] _0390_ gamelogic.setWord\[6\] _0385_ vssd1 vssd1 vccd1
+ vccd1 _1279_ sky130_fd_sc_hd__a22o_1
XFILLER_0_6_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2647_ hostdisp.bottom\[55\] net114 _1095_ hostdisp.top\[79\] vssd1 vssd1 vccd1 vccd1
+ _1218_ sky130_fd_sc_hd__a22o_1
XFILLER_0_14_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_168_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2578_ _1150_ _1151_ _1152_ net226 vssd1 vssd1 vccd1 vccd1 _1153_ sky130_fd_sc_hd__o31a_1
X_1529_ _0473_ _0474_ _0475_ _0476_ vssd1 vssd1 vccd1 vccd1 _0477_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_161_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_38_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_182_Right_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2959__A2 net53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_14_Right_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_172_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2592__B1 net108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_23_Right_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2647__B2 hostdisp.top\[79\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_148 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3457__SET_B net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_32_Right_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1880_ _0739_ net116 _0738_ vssd1 vssd1 vccd1 vccd1 uart_transmitter.next_clk_count\[4\]
+ sky130_fd_sc_hd__and3b_1
XFILLER_0_113_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3550_ clknet_leaf_6_clk hostdisp.next_curr_guesses\[32\] net191 vssd1 vssd1 vccd1
+ vccd1 hostdisp.curr_guesses\[32\] sky130_fd_sc_hd__dfstp_1
XFILLER_0_98_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2501_ net138 net139 _1061_ _1068_ vssd1 vssd1 vccd1 vccd1 _1079_ sky130_fd_sc_hd__and4_1
XFILLER_0_11_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3481_ clknet_leaf_32_clk hostdisp.next_curr_word\[3\] net164 vssd1 vssd1 vccd1 vccd1
+ hostdisp.curr_word\[3\] sky130_fd_sc_hd__dfstp_1
XPHY_EDGE_ROW_41_Right_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2432_ hostdisp.curr_word\[14\] net119 vssd1 vssd1 vccd1 vccd1 _1038_ sky130_fd_sc_hd__or2_1
X_2363_ net456 _0998_ net167 vssd1 vssd1 vccd1 vccd1 _1001_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_47_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2294_ lcdPlayer.cnt_500hz\[3\] _0750_ vssd1 vssd1 vccd1 vccd1 _0960_ sky130_fd_sc_hd__or2_1
XANTENNA__2638__B2 hostdisp.top\[46\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2545__S net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_50_Right_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_176_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_170_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2574__B1 _1078_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_186_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout51_A net52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2190__S net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_150_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2096__A2 net96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3442__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2981_ gamelogic.setWord\[20\] net52 net48 gamelogic.setWord\[28\] vssd1 vssd1 vccd1
+ vccd1 _0344_ sky130_fd_sc_hd__o22a_1
XFILLER_0_33_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_173_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1932_ _0183_ _0770_ vssd1 vssd1 vccd1 vccd1 _0780_ sky130_fd_sc_hd__nand2_1
X_1863_ net271 _0731_ vssd1 vssd1 vccd1 vccd1 clock_div.next_count\[29\] sky130_fd_sc_hd__xnor2_1
XFILLER_0_126_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3602_ net236 vssd1 vssd1 vccd1 vccd1 gpio_out[2] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_40_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1794_ clock_div.count\[6\] clock_div.count\[8\] _0688_ _0691_ vssd1 vssd1 vccd1
+ vccd1 _0692_ sky130_fd_sc_hd__or4_1
XANTENNA__2556__B1 net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3533_ clknet_leaf_14_clk net382 net206 vssd1 vssd1 vccd1 vccd1 hostdisp.curr_guesses\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3464_ clknet_leaf_2_clk _0342_ net175 vssd1 vssd1 vccd1 vccd1 gamelogic.setWord\[26\]
+ sky130_fd_sc_hd__dfstp_1
X_2415_ hostdisp.curr_word\[1\] net72 net69 net412 vssd1 vssd1 vccd1 vccd1 _0133_
+ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_35_clk_X clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3395_ clknet_leaf_20_clk _0284_ net212 vssd1 vssd1 vccd1 vccd1 dispFSM.guesses\[49\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_149_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2346_ _0619_ _0621_ net149 net150 vssd1 vssd1 vccd1 vccd1 _0992_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout186_A net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2277_ _0945_ vssd1 vssd1 vccd1 vccd1 _0946_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_62 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_164_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_32_clk clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_32_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout141_X net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2547__B1 _0758_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3315__CLK clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout99_A net100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_167_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_11_Left_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_46_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_155_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_23_clk clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_23_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_53_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2538__B1 _0360_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_20_Left_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2214__A net100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2200_ net131 hostdisp.curr_guesses\[42\] net122 _0902_ vssd1 vssd1 vccd1 vccd1 hostdisp.nextBottom\[82\]
+ sky130_fd_sc_hd__a31o_1
XANTENNA__3377__RESET_B net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3180_ clknet_leaf_31_clk _0156_ net174 vssd1 vssd1 vccd1 vccd1 hostdisp.top\[64\]
+ sky130_fd_sc_hd__dfrtp_1
X_2131_ gamelogic.setWord\[8\] hostdisp.curr_guesses\[8\] net124 vssd1 vssd1 vccd1
+ vccd1 _0868_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2062_ hostdisp.curr_word\[8\] net102 net75 _0838_ gamelogic.indexCorrect\[1\] vssd1
+ vssd1 vccd1 vccd1 _0839_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_146_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_87 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2964_ gamelogic.setWord\[3\] net51 net47 gamelogic.setWord\[11\] vssd1 vssd1 vccd1
+ vccd1 _0327_ sky130_fd_sc_hd__o22a_1
XANTENNA__3513__SET_B net165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_14_clk clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_14_clk
+ sky130_fd_sc_hd__clkbuf_8
X_1915_ net166 _0767_ vssd1 vssd1 vccd1 vccd1 _0768_ sky130_fd_sc_hd__nand2_1
XFILLER_0_173_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2895_ dispFSM.guesses\[35\] net81 net57 net528 vssd1 vssd1 vccd1 vccd1 _0262_ sky130_fd_sc_hd__o22a_1
X_1846_ net467 _0721_ vssd1 vssd1 vccd1 vccd1 _0722_ sky130_fd_sc_hd__nor2_1
XFILLER_0_114_212 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3338__CLK clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_155_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1777_ uart_transmitter.bit_index\[1\] _0402_ message_reg.msg\[2\] _0675_ vssd1 vssd1
+ vccd1 vccd1 _0676_ sky130_fd_sc_hd__a31o_1
XFILLER_0_114_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3516_ clknet_leaf_31_clk hostdisp.next_curr_word\[38\] net165 vssd1 vssd1 vccd1
+ vccd1 hostdisp.curr_word\[38\] sky130_fd_sc_hd__dfstp_1
XFILLER_0_69_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout101_A net104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_4_Right_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_176_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3447_ clknet_leaf_13_clk _0325_ net197 vssd1 vssd1 vccd1 vccd1 gamelogic.setWord\[9\]
+ sky130_fd_sc_hd__dfstp_2
XANTENNA__3488__CLK clknet_leaf_30_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_15_clk_A clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3378_ clknet_leaf_23_clk _0267_ net182 vssd1 vssd1 vccd1 vccd1 dispFSM.guesses\[32\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_176_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2329_ lcdPlayer.cnt_500hz\[16\] _0980_ vssd1 vssd1 vccd1 vccd1 _0982_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_68_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_149_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_268 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_117_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_8_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2209__A net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2643__S net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2471__A2 net75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1700_ keypadFSMPlayer.state\[0\] _0453_ _0587_ keypadFSMPlayer.state\[4\] _0616_
+ vssd1 vssd1 vccd1 vccd1 _0011_ sky130_fd_sc_hd__a221o_1
X_2680_ gamelogic.setWord\[35\] _0380_ gamelogic.setWord\[39\] _0386_ _1245_ vssd1
+ vssd1 vccd1 vccd1 _1246_ sky130_fd_sc_hd__o221a_1
XFILLER_0_26_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_14_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1631_ keypadHostt.scan_col\[3\] _0546_ _0366_ vssd1 vssd1 vccd1 vccd1 _0566_ sky130_fd_sc_hd__a21o_1
XFILLER_0_41_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1562_ _0496_ _0502_ _0503_ vssd1 vssd1 vccd1 vccd1 _0510_ sky130_fd_sc_hd__or3_1
X_3301_ clknet_leaf_34_clk uart_receiver.temp_byte\[1\] net159 vssd1 vssd1 vccd1 vccd1
+ buffer.Rx_byte\[1\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_187_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1493_ _0426_ _0430_ vssd1 vssd1 vccd1 vccd1 _0445_ sky130_fd_sc_hd__nor2_1
XFILLER_0_190_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3232_ clknet_leaf_13_clk _0206_ net197 vssd1 vssd1 vccd1 vccd1 host_message_reg.setLetter\[1\]
+ sky130_fd_sc_hd__dfstp_1
Xclkbuf_leaf_3_clk clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_3_clk
+ sky130_fd_sc_hd__clkbuf_8
X_3163_ clknet_leaf_29_clk _0139_ net166 vssd1 vssd1 vccd1 vccd1 hostdisp.top\[47\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_2_2__f_clk_X clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2114_ _0827_ _0857_ vssd1 vssd1 vccd1 vccd1 _0859_ sky130_fd_sc_hd__or2_1
XFILLER_0_146_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3094_ clknet_leaf_27_clk _0084_ vssd1 vssd1 vccd1 vccd1 lcdPlayer.cnt_500hz\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__2447__C1 net67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_65_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2045_ _0827_ _0829_ vssd1 vssd1 vccd1 vccd1 _0830_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_105_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2462__A2 net70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_146_156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2947_ dispFSM.msg\[7\] net88 net65 net482 vssd1 vssd1 vccd1 vccd1 _0314_ sky130_fd_sc_hd__a22o_1
XFILLER_0_17_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2878_ dispFSM.guesses\[18\] net84 net58 net469 vssd1 vssd1 vccd1 vccd1 _0245_ sky130_fd_sc_hd__o22a_1
XFILLER_0_4_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1693__A keypadFSMHost.state\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1829_ clock_div.count\[15\] _0711_ vssd1 vssd1 vccd1 vccd1 _0712_ sky130_fd_sc_hd__and2_1
XFILLER_0_142_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout104_X net104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_5_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_164_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_79_Right_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2438__C1 _1034_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2989__B1 net48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3503__CLK clknet_leaf_30_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_177_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2453__A2 net67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_175_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1964__A1 net2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_88_Right_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2699__A net140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_97_Right_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_182_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2692__A2 gamelogic.setWord\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3183__CLK clknet_leaf_30_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2444__A2 net67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_141_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_183_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2801_ _0385_ gamelogic.setWord\[14\] _1344_ _1346_ vssd1 vssd1 vccd1 vccd1 _1347_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_26_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_193_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2732_ net404 net233 _1287_ vssd1 vssd1 vccd1 vccd1 _0203_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1955__A1 host_message_reg.Cstate vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_4_Left_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2663_ _0398_ _0662_ _0664_ uart_transmitter.bit_index\[0\] vssd1 vssd1 vccd1 vccd1
+ _1232_ sky130_fd_sc_hd__o31a_1
X_1614_ net153 _0548_ vssd1 vssd1 vccd1 vccd1 _0549_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_152_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2594_ dispFSM.guesses\[28\] net115 _1084_ dispFSM.guesses\[4\] vssd1 vssd1 vccd1
+ vccd1 _1168_ sky130_fd_sc_hd__a22o_1
X_1545_ _0372_ _1399_ keypadFSMPlayer.state\[1\] vssd1 vssd1 vccd1 vccd1 _0493_ sky130_fd_sc_hd__a21oi_1
Xfanout229 net231 vssd1 vssd1 vccd1 vccd1 net229 sky130_fd_sc_hd__buf_2
Xfanout218 net224 vssd1 vssd1 vccd1 vccd1 net218 sky130_fd_sc_hd__clkbuf_2
Xfanout207 net209 vssd1 vssd1 vccd1 vccd1 net207 sky130_fd_sc_hd__clkbuf_4
X_1476_ net229 net6 _0427_ vssd1 vssd1 vccd1 vccd1 _0428_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_163_Right_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3215_ clknet_leaf_19_clk _0191_ net212 vssd1 vssd1 vccd1 vccd1 uart_transmitter.bit_index\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3526__CLK clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3146_ clknet_leaf_25_clk _0122_ vssd1 vssd1 vccd1 vccd1 lcdPlayer.cnt_20ms\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_3077_ clknet_leaf_33_clk net318 net161 vssd1 vssd1 vccd1 vccd1 buffer.temp_guess\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2028_ hostdisp.curr_guesses\[42\] net91 net76 net504 vssd1 vssd1 vccd1 vccd1 hostdisp.next_curr_guesses\[34\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_166_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1688__A _0607_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_174_273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout221_X net221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold250 hostdisp.curr_word\[7\] vssd1 vssd1 vccd1 vccd1 net514 sky130_fd_sc_hd__dlygate4sd3_1
Xhold261 hostdisp.top\[78\] vssd1 vssd1 vccd1 vccd1 net525 sky130_fd_sc_hd__dlygate4sd3_1
Xhold272 dispFSM.guesses\[65\] vssd1 vssd1 vccd1 vccd1 net536 sky130_fd_sc_hd__dlygate4sd3_1
Xhold294 hostdisp.top\[76\] vssd1 vssd1 vccd1 vccd1 net558 sky130_fd_sc_hd__dlygate4sd3_1
Xhold283 dispFSM.guesses\[16\] vssd1 vssd1 vccd1 vccd1 net547 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_130_Right_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_76_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2193__S net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_180_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_310 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3549__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3000_ net221 vssd1 vssd1 vccd1 vccd1 _0025_ sky130_fd_sc_hd__inv_2
XFILLER_0_127_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput7 gpio_in[33] vssd1 vssd1 vccd1 vccd1 net7 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_188_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_102_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1711__C_N host_message_reg.Cstate vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1795__X _0693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2715_ net143 gamelogic.setWord\[3\] vssd1 vssd1 vccd1 vccd1 _1278_ sky130_fd_sc_hd__xnor2_1
XANTENNA__3079__CLK clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2646_ hostdisp.bottom\[87\] net117 _1096_ hostdisp.top\[71\] vssd1 vssd1 vccd1 vccd1
+ _1217_ sky130_fd_sc_hd__a22o_1
XFILLER_0_168_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2577_ dispFSM.guesses\[59\] net117 net113 dispFSM.guesses\[51\] _1148_ vssd1 vssd1
+ vccd1 vccd1 _1152_ sky130_fd_sc_hd__a221o_1
XFILLER_0_168_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1528_ keypadFSMPlayer.prev_key\[6\] _0416_ _0424_ vssd1 vssd1 vccd1 vccd1 _0476_
+ sky130_fd_sc_hd__or3b_1
X_1459_ hostdisp.curr_word\[37\] vssd1 vssd1 vccd1 vccd1 _0412_ sky130_fd_sc_hd__inv_2
XFILLER_0_184_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2105__B2 net144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_184_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2656__A2 _1072_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_161_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3129_ clknet_leaf_18_clk uart_transmitter.next_clk_count\[9\] net219 vssd1 vssd1
+ vccd1 vccd1 uart_transmitter.clk_count\[9\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_38_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_162_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_172_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2041__B1 net80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2592__A1 hostdisp.top\[44\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_92_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2188__S net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2647__A2 net114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_185_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_85_Left_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_153_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3572__256 vssd1 vssd1 vccd1 vccd1 net256 _3572__256/LO sky130_fd_sc_hd__conb_1
XFILLER_0_153_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2032__B1 net79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3480_ clknet_leaf_31_clk hostdisp.next_curr_word\[2\] net164 vssd1 vssd1 vccd1 vccd1
+ hostdisp.curr_word\[2\] sky130_fd_sc_hd__dfstp_1
X_2500_ _1070_ _1074_ vssd1 vssd1 vccd1 vccd1 _1078_ sky130_fd_sc_hd__nor2_4
X_2431_ hostdisp.curr_word\[13\] _1031_ net67 net272 vssd1 vssd1 vccd1 vccd1 _0145_
+ sky130_fd_sc_hd__o22a_1
XPHY_EDGE_ROW_94_Left_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2362_ lcdPlayer.cnt_20ms\[7\] _0998_ vssd1 vssd1 vccd1 vccd1 _1000_ sky130_fd_sc_hd__and2_1
X_2293_ _0750_ _0955_ _0959_ vssd1 vssd1 vccd1 vccd1 _0085_ sky130_fd_sc_hd__and3b_1
XANTENNA__2638__A2 net114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_188_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_191_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_176_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_240 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout229_A net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout131_A net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2629_ _1181_ _1185_ _1201_ vssd1 vssd1 vccd1 vccd1 _1202_ sky130_fd_sc_hd__a21o_1
XANTENNA__2797__A gamelogic.letter\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_167_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3244__CLK clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_243 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2014__B1 net77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3394__CLK clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2043__Y _0828_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkload7_A clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2980_ gamelogic.setWord\[19\] net51 net47 gamelogic.setWord\[27\] vssd1 vssd1 vccd1
+ vccd1 _0343_ sky130_fd_sc_hd__o22a_1
XFILLER_0_56_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1931_ _0187_ _0777_ vssd1 vssd1 vccd1 vccd1 _0779_ sky130_fd_sc_hd__and2_1
XFILLER_0_173_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1862_ _0730_ _0731_ vssd1 vssd1 vccd1 vccd1 clock_div.next_count\[28\] sky130_fd_sc_hd__and2b_1
X_3601_ net235 vssd1 vssd1 vccd1 vccd1 gpio_out[1] sky130_fd_sc_hd__buf_2
XFILLER_0_126_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_40_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2005__B1 net77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_181_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1793_ clock_div.count\[2\] clock_div.count\[4\] _0689_ _0690_ vssd1 vssd1 vccd1
+ vccd1 _0691_ sky130_fd_sc_hd__or4_1
XFILLER_0_3_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3532_ clknet_leaf_6_clk hostdisp.next_curr_guesses\[14\] net191 vssd1 vssd1 vccd1
+ vccd1 hostdisp.curr_guesses\[14\] sky130_fd_sc_hd__dfstp_1
X_3463_ clknet_leaf_7_clk _0341_ net195 vssd1 vssd1 vccd1 vccd1 gamelogic.setWord\[25\]
+ sky130_fd_sc_hd__dfstp_2
X_2414_ hostdisp.curr_word\[0\] net72 net69 net397 vssd1 vssd1 vccd1 vccd1 _0132_
+ sky130_fd_sc_hd__a22o_1
X_3394_ clknet_leaf_23_clk _0283_ net183 vssd1 vssd1 vccd1 vccd1 dispFSM.guesses\[48\]
+ sky130_fd_sc_hd__dfstp_1
X_2345_ _0622_ _0991_ _0618_ vssd1 vssd1 vccd1 vccd1 _0105_ sky130_fd_sc_hd__and3b_1
XANTENNA__3536__SET_B net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2276_ lcdPlayer.cnt_20ms\[3\] lcdPlayer.cnt_20ms\[2\] lcdPlayer.cnt_20ms\[1\] lcdPlayer.cnt_20ms\[0\]
+ vssd1 vssd1 vccd1 vccd1 _0945_ sky130_fd_sc_hd__and4_1
XFILLER_0_74_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_108_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout179_A net180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_176_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_191_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_174 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_167_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_54_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_178_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_159_Left_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2786__A1 host_message_reg.setLetter\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_168_Left_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2130_ net345 net120 _0867_ net136 vssd1 vssd1 vccd1 vccd1 hostdisp.nextBottom\[47\]
+ sky130_fd_sc_hd__o211a_1
X_2061_ hostdisp.curr_word\[9\] hostdisp.curr_word\[10\] _0406_ hostdisp.curr_word\[14\]
+ net102 vssd1 vssd1 vccd1 vccd1 _0838_ sky130_fd_sc_hd__a41o_1
XFILLER_0_135_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_266 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_177_Left_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_173_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2963_ gamelogic.setWord\[2\] net51 net47 gamelogic.setWord\[10\] vssd1 vssd1 vccd1
+ vccd1 _0326_ sky130_fd_sc_hd__o22a_1
XFILLER_0_56_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1914_ lcdPlayer.nextState\[1\] lcdPlayer.currentState\[1\] _0764_ vssd1 vssd1 vccd1
+ vccd1 _0767_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2894_ dispFSM.guesses\[34\] net84 net59 net511 vssd1 vssd1 vccd1 vccd1 _0261_ sky130_fd_sc_hd__o22a_1
X_1845_ _0720_ _0721_ vssd1 vssd1 vccd1 vccd1 clock_div.next_count\[21\] sky130_fd_sc_hd__nor2_1
XFILLER_0_114_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2529__A1 dispFSM.msg\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_155_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1776_ _0401_ _0673_ _0674_ vssd1 vssd1 vccd1 vccd1 _0675_ sky130_fd_sc_hd__a21o_1
XFILLER_0_71_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkload33_A clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2411__Y _1031_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3515_ clknet_leaf_29_clk hostdisp.next_curr_word\[37\] net169 vssd1 vssd1 vccd1
+ vccd1 hostdisp.curr_word\[37\] sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_186_Left_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3446_ clknet_leaf_5_clk _0324_ net196 vssd1 vssd1 vccd1 vccd1 gamelogic.setWord\[8\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_176_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3377_ clknet_leaf_21_clk net451 net202 vssd1 vssd1 vccd1 vccd1 dispFSM.guesses\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_176_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2328_ net287 _0978_ _0981_ vssd1 vssd1 vccd1 vccd1 _0098_ sky130_fd_sc_hd__o21a_1
XFILLER_0_192_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2259_ net297 buffer.temp_guess\[5\] _0630_ vssd1 vssd1 vccd1 vccd1 _0072_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_68_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_51_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_177_Right_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_268 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2940__A1 dispFSM.msg\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2209__B gamelogic.setWord\[39\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_170_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1630_ _0537_ _0564_ vssd1 vssd1 vccd1 vccd1 _0565_ sky130_fd_sc_hd__nand2_2
XPHY_EDGE_ROW_144_Right_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1561_ _0495_ _0508_ _0490_ vssd1 vssd1 vccd1 vccd1 _0509_ sky130_fd_sc_hd__and3b_1
X_3300_ clknet_leaf_33_clk uart_receiver.temp_byte\[0\] net158 vssd1 vssd1 vccd1 vccd1
+ buffer.Rx_byte\[0\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_187_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1492_ keypadFSMPlayer.strobe_edge1 keypadFSMPlayer.strobe_edge vssd1 vssd1 vccd1
+ vccd1 _0444_ sky130_fd_sc_hd__nand2b_1
X_3231_ clknet_leaf_13_clk _0205_ net197 vssd1 vssd1 vccd1 vccd1 host_message_reg.setLetter\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_39_77 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3162_ clknet_leaf_31_clk _0138_ net163 vssd1 vssd1 vccd1 vccd1 hostdisp.top\[46\]
+ sky130_fd_sc_hd__dfrtp_1
X_2113_ _0827_ _0857_ vssd1 vssd1 vccd1 vccd1 _0858_ sky130_fd_sc_hd__nor2_1
XFILLER_0_178_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3093_ clknet_leaf_27_clk _0083_ vssd1 vssd1 vccd1 vccd1 lcdPlayer.cnt_500hz\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_178_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2044_ net133 _0822_ vssd1 vssd1 vccd1 vccd1 _0829_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_105_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3305__CLK clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_157_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_146_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2946_ dispFSM.msg\[6\] net85 net62 net495 vssd1 vssd1 vccd1 vccd1 _0313_ sky130_fd_sc_hd__o22a_1
XFILLER_0_127_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2877_ dispFSM.guesses\[17\] net86 net62 net532 vssd1 vssd1 vccd1 vccd1 _0244_ sky130_fd_sc_hd__o22a_1
XFILLER_0_154_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1828_ _0710_ _0711_ vssd1 vssd1 vccd1 vccd1 clock_div.next_count\[14\] sky130_fd_sc_hd__nor2_1
XANTENNA__3455__CLK clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_330 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2422__X _1034_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_111_Right_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1759_ message_reg.state\[0\] uart_transmitter.state\[0\] vssd1 vssd1 vccd1 vccd1
+ _0661_ sky130_fd_sc_hd__nand2_1
XFILLER_0_102_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3429_ clknet_leaf_29_clk _0003_ vssd1 vssd1 vccd1 vccd1 lcdPlayer.nextState\[4\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_5_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_164_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_177_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_123_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_175_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2045__A _0827_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2610__B1 _1106_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3328__CLK clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2800_ _0378_ gamelogic.setWord\[9\] _0394_ gamelogic.letter\[5\] _1345_ vssd1 vssd1
+ vccd1 vccd1 _1346_ sky130_fd_sc_hd__o221a_1
XFILLER_0_41_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3478__CLK clknet_leaf_31_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_193_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2731_ net366 _0553_ _1287_ vssd1 vssd1 vccd1 vccd1 _0202_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_14_clk_A clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2062__D1 gamelogic.indexCorrect\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1955__A2 net97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2662_ net266 _0936_ _0937_ vssd1 vssd1 vccd1 vccd1 _0188_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_10_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_136 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1613_ _0542_ _0545_ _0547_ vssd1 vssd1 vccd1 vccd1 _0548_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_152_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2593_ dispFSM.guesses\[12\] _1078_ net110 dispFSM.guesses\[36\] vssd1 vssd1 vccd1
+ vccd1 _1167_ sky130_fd_sc_hd__a22o_1
XFILLER_0_41_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_29_clk_A clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1544_ _0491_ keypadFSMPlayer.state\[5\] vssd1 vssd1 vccd1 vccd1 _0492_ sky130_fd_sc_hd__nand2b_1
Xfanout219 net221 vssd1 vssd1 vccd1 vccd1 net219 sky130_fd_sc_hd__clkbuf_4
Xfanout208 net209 vssd1 vssd1 vccd1 vccd1 net208 sky130_fd_sc_hd__clkbuf_4
X_1475_ net155 net128 vssd1 vssd1 vccd1 vccd1 _0427_ sky130_fd_sc_hd__and2_1
XFILLER_0_157_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3214_ clknet_leaf_19_clk _0190_ net211 vssd1 vssd1 vccd1 vccd1 uart_transmitter.bit_index\[0\]
+ sky130_fd_sc_hd__dfrtp_4
X_3582__258 vssd1 vssd1 vccd1 vccd1 net258 _3582__258/LO sky130_fd_sc_hd__conb_1
XPHY_EDGE_ROW_105_Left_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3145_ clknet_leaf_25_clk _0121_ vssd1 vssd1 vccd1 vccd1 lcdPlayer.cnt_20ms\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_3076_ clknet_leaf_11_clk _0066_ net216 vssd1 vssd1 vccd1 vccd1 keypadFSMHost.unlocked
+ sky130_fd_sc_hd__dfrtp_1
X_2027_ hostdisp.curr_guesses\[41\] net93 net78 net462 vssd1 vssd1 vccd1 vccd1 hostdisp.next_curr_guesses\[33\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_89_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2929_ net430 net90 net64 net453 vssd1 vssd1 vccd1 vccd1 _0296_ sky130_fd_sc_hd__a22o_1
XFILLER_0_142_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_170_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold262 dispFSM.guesses\[41\] vssd1 vssd1 vccd1 vccd1 net526 sky130_fd_sc_hd__dlygate4sd3_1
Xhold251 dispFSM.guesses\[73\] vssd1 vssd1 vccd1 vccd1 net515 sky130_fd_sc_hd__dlygate4sd3_1
Xhold240 hostdisp.curr_guesses\[34\] vssd1 vssd1 vccd1 vccd1 net504 sky130_fd_sc_hd__dlygate4sd3_1
Xhold295 hostdisp.top\[42\] vssd1 vssd1 vccd1 vccd1 net559 sky130_fd_sc_hd__dlygate4sd3_1
Xhold273 dispFSM.guesses\[40\] vssd1 vssd1 vccd1 vccd1 net537 sky130_fd_sc_hd__dlygate4sd3_1
Xhold284 hostdisp.curr_guesses\[26\] vssd1 vssd1 vccd1 vccd1 net548 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_16_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_180_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_180_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_322 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput8 nrst vssd1 vssd1 vccd1 vccd1 net8 sky130_fd_sc_hd__buf_1
XFILLER_0_127_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_188_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_188_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_102_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2714_ net141 gamelogic.setWord\[5\] vssd1 vssd1 vccd1 vccd1 _1277_ sky130_fd_sc_hd__xnor2_1
XANTENNA__2413__A net97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2050__A1 net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2645_ net296 net107 _1216_ net203 vssd1 vssd1 vccd1 vccd1 _0180_ sky130_fd_sc_hd__o211a_1
X_2576_ dispFSM.guesses\[3\] _1084_ _1086_ dispFSM.guesses\[75\] vssd1 vssd1 vccd1
+ vccd1 _1151_ sky130_fd_sc_hd__a22o_1
X_1527_ net229 net232 net154 _0424_ _0359_ vssd1 vssd1 vccd1 vccd1 _0475_ sky130_fd_sc_hd__a41o_1
XPHY_EDGE_ROW_113_Left_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1458_ hostdisp.curr_word\[31\] vssd1 vssd1 vccd1 vccd1 _0411_ sky130_fd_sc_hd__inv_2
XFILLER_0_184_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3128_ clknet_leaf_18_clk uart_transmitter.next_clk_count\[8\] net219 vssd1 vssd1
+ vccd1 vccd1 uart_transmitter.clk_count\[8\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3059_ clknet_leaf_16_clk _0052_ _0021_ vssd1 vssd1 vccd1 vccd1 keypadFSMPlayer.prev_key\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_38_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout164_X net164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_122_Left_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_120_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_147_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_172_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_21_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2041__A1 net140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_300 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_220 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2592__A2 _1098_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_163 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3173__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_131_Left_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout77_X net77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1402__A net139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1607__A1 net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_140_Left_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_190_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3516__CLK clknet_leaf_31_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2430_ hostdisp.curr_word\[12\] net73 net70 net309 vssd1 vssd1 vccd1 vccd1 _0144_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_121_196 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2361_ _0998_ _0999_ vssd1 vssd1 vccd1 vccd1 _0113_ sky130_fd_sc_hd__nor2_1
X_2292_ lcdPlayer.cnt_500hz\[0\] lcdPlayer.cnt_500hz\[1\] lcdPlayer.cnt_500hz\[2\]
+ vssd1 vssd1 vccd1 vccd1 _0959_ sky130_fd_sc_hd__a21o_1
XFILLER_0_188_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3046__CLK clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_252 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2810__A3 _1355_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout124_A net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3196__CLK clknet_leaf_30_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2574__A2 _1072_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2628_ _1159_ _1197_ _1199_ _1200_ vssd1 vssd1 vccd1 vccd1 _1201_ sky130_fd_sc_hd__or4_1
XFILLER_0_2_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2559_ dispFSM.guesses\[50\] net112 _1084_ dispFSM.guesses\[2\] _1132_ vssd1 vssd1
+ vccd1 vccd1 _1135_ sky130_fd_sc_hd__a221o_1
XANTENNA__1921__S _0764_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_175_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3539__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1930_ _0773_ _0776_ vssd1 vssd1 vccd1 vccd1 _0778_ sky130_fd_sc_hd__nor2_1
X_1861_ clock_div.count\[28\] _0729_ vssd1 vssd1 vccd1 vccd1 _0731_ sky130_fd_sc_hd__nand2_1
XFILLER_0_16_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3600_ net234 vssd1 vssd1 vccd1 vccd1 gpio_out[0] sky130_fd_sc_hd__buf_2
XFILLER_0_181_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1792_ clock_div.count\[7\] clock_div.count\[9\] vssd1 vssd1 vccd1 vccd1 _0690_ sky130_fd_sc_hd__nand2_1
X_3531_ clknet_leaf_15_clk hostdisp.next_curr_guesses\[13\] net208 vssd1 vssd1 vccd1
+ vccd1 hostdisp.curr_guesses\[13\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_141_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2556__A2 _1072_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3462_ clknet_leaf_5_clk _0340_ net196 vssd1 vssd1 vccd1 vccd1 gamelogic.setWord\[24\]
+ sky130_fd_sc_hd__dfstp_1
X_3393_ clknet_leaf_15_clk _0282_ net207 vssd1 vssd1 vccd1 vccd1 dispFSM.guesses\[47\]
+ sky130_fd_sc_hd__dfrtp_1
X_2413_ net97 net95 vssd1 vssd1 vccd1 vccd1 _1033_ sky130_fd_sc_hd__nand2_1
XANTENNA__2410__B net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2344_ net150 _0621_ net149 vssd1 vssd1 vccd1 vccd1 _0991_ sky130_fd_sc_hd__a21o_1
XFILLER_0_165_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2275_ lcdPlayer.cnt_20ms\[2\] lcdPlayer.cnt_20ms\[1\] lcdPlayer.cnt_20ms\[0\] vssd1
+ vssd1 vccd1 vccd1 _0944_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_108_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_164_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_158_Right_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_191_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_191_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_94 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_167_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3211__CLK clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3361__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_178_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_125_Right_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_163_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2060_ hostdisp.curr_word\[11\] hostdisp.curr_word\[12\] _0407_ net102 vssd1 vssd1
+ vccd1 vccd1 _0837_ sky130_fd_sc_hd__a31o_1
XFILLER_0_88_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_278 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2962_ gamelogic.setWord\[1\] net54 net50 gamelogic.setWord\[9\] vssd1 vssd1 vccd1
+ vccd1 _0325_ sky130_fd_sc_hd__o22a_1
XFILLER_0_173_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1913_ _0765_ vssd1 vssd1 vccd1 vccd1 _0766_ sky130_fd_sc_hd__inv_2
X_2893_ dispFSM.guesses\[33\] net86 net63 net549 vssd1 vssd1 vccd1 vccd1 _0260_ sky130_fd_sc_hd__o22a_1
X_1844_ clock_div.count\[21\] clock_div.count\[20\] _0719_ vssd1 vssd1 vccd1 vccd1
+ _0721_ sky130_fd_sc_hd__and3_1
XFILLER_0_4_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1775_ uart_transmitter.bit_index\[1\] uart_transmitter.bit_index\[0\] message_reg.msg\[3\]
+ uart_transmitter.bit_index\[2\] vssd1 vssd1 vccd1 vccd1 _0674_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_155_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3514_ clknet_leaf_31_clk hostdisp.next_curr_word\[36\] net165 vssd1 vssd1 vccd1
+ vccd1 hostdisp.curr_word\[36\] sky130_fd_sc_hd__dfstp_1
X_3445_ clknet_leaf_14_clk _0323_ net193 vssd1 vssd1 vccd1 vccd1 gamelogic.setWord\[7\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_100_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3376_ clknet_leaf_20_clk _0265_ net204 vssd1 vssd1 vccd1 vccd1 dispFSM.guesses\[30\]
+ sky130_fd_sc_hd__dfstp_1
X_2327_ net74 _0980_ vssd1 vssd1 vccd1 vccd1 _0981_ sky130_fd_sc_hd__nor2_1
XFILLER_0_33_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2258_ net303 buffer.temp_guess\[4\] net127 vssd1 vssd1 vccd1 vccd1 _0071_ sky130_fd_sc_hd__mux2_1
XFILLER_0_192_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2189_ gamelogic.setWord\[37\] hostdisp.curr_guesses\[37\] net125 vssd1 vssd1 vccd1
+ vccd1 _0897_ sky130_fd_sc_hd__mux2_1
XFILLER_0_192_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_0_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_0_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1560_ net147 _0507_ _0429_ vssd1 vssd1 vccd1 vccd1 _0508_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3257__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_187_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1491_ keypadFSMPlayer.strobe_edge1 keypadFSMPlayer.strobe_edge vssd1 vssd1 vccd1
+ vccd1 _0443_ sky130_fd_sc_hd__and2b_2
X_3230_ clknet_leaf_11_clk _0204_ net217 vssd1 vssd1 vccd1 vccd1 keypadFSMHost.prev_key\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2695__A1 _1252_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3161_ clknet_leaf_30_clk _0137_ net181 vssd1 vssd1 vccd1 vccd1 hostdisp.top\[45\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_176_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2112_ gamelogic.incorrect\[0\] gamelogic.incorrect\[1\] gamelogic.incorrect\[2\]
+ vssd1 vssd1 vccd1 vccd1 _0857_ sky130_fd_sc_hd__and3b_1
X_3092_ clknet_leaf_21_clk _0082_ net210 vssd1 vssd1 vccd1 vccd1 message_reg.msg\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__2447__B2 _1031_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2447__A1 net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2043_ net129 _0821_ vssd1 vssd1 vccd1 vccd1 _0828_ sky130_fd_sc_hd__nor2_4
XTAP_TAPCELL_ROW_105_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2945_ dispFSM.msg\[5\] net90 net64 net426 vssd1 vssd1 vccd1 vccd1 _0312_ sky130_fd_sc_hd__a22o_1
XFILLER_0_17_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2876_ dispFSM.guesses\[16\] net81 net56 net512 vssd1 vssd1 vccd1 vccd1 _0243_ sky130_fd_sc_hd__o22a_1
X_1827_ clock_div.count\[13\] clock_div.count\[14\] _0709_ vssd1 vssd1 vccd1 vccd1
+ _0711_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_13_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1758_ net535 _0658_ _0660_ vssd1 vssd1 vccd1 vccd1 uart_receiver.next_clk_count\[10\]
+ sky130_fd_sc_hd__o21a_1
X_1689_ keypadFSMHost.state\[0\] _0592_ _0606_ keypadFSMHost.state\[4\] _0611_ vssd1
+ vssd1 vccd1 vccd1 _0005_ sky130_fd_sc_hd__a221o_1
XANTENNA__1990__A net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3428_ clknet_leaf_29_clk _0002_ vssd1 vssd1 vccd1 vccd1 lcdPlayer.nextState\[2\]
+ sky130_fd_sc_hd__dfxtp_2
X_3359_ clknet_leaf_20_clk _0248_ net203 vssd1 vssd1 vccd1 vccd1 dispFSM.guesses\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_5_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_164_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1989__X _0822_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2438__A1 net130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2438__B2 _0830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3600__234 vssd1 vssd1 vccd1 vccd1 _3600__234/HI net234 sky130_fd_sc_hd__conb_1
XANTENNA__2989__A2 net52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_184_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_123_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_192_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_175_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_192_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_160_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_95_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2507__Y _1085_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_17_Left_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2730_ net387 net3 _1287_ vssd1 vssd1 vccd1 vccd1 _0201_ sky130_fd_sc_hd__mux2_1
XFILLER_0_143_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2601__B2 net105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2601__A1 net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_193_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2661_ net299 net107 _1231_ net187 vssd1 vssd1 vccd1 vccd1 _0181_ sky130_fd_sc_hd__o211a_1
X_1612_ keypadHostt.scan_col\[3\] keypadHostt.scan_col\[2\] vssd1 vssd1 vccd1 vccd1
+ _0547_ sky130_fd_sc_hd__or2_2
XFILLER_0_41_148 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_295 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2592_ hostdisp.top\[44\] _1098_ net108 hostdisp.top\[60\] _1165_ vssd1 vssd1 vccd1
+ vccd1 _1166_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_10_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1543_ _0430_ _0438_ _0436_ vssd1 vssd1 vccd1 vccd1 _0491_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_152_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_26_Left_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1474_ net4 _0417_ _0425_ vssd1 vssd1 vccd1 vccd1 _0426_ sky130_fd_sc_hd__or3_2
Xfanout209 net212 vssd1 vssd1 vccd1 vccd1 net209 sky130_fd_sc_hd__clkbuf_2
X_3213_ clknet_leaf_17_clk _0189_ _0038_ vssd1 vssd1 vccd1 vccd1 keypadFSMPlayer.unlocked
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_157_67 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3144_ clknet_leaf_25_clk _0120_ vssd1 vssd1 vccd1 vccd1 lcdPlayer.cnt_20ms\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_3075_ clknet_leaf_17_clk keypadFSMPlayer.next_state\[2\] _0037_ vssd1 vssd1 vccd1
+ vccd1 _1401_ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_173_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2026_ hostdisp.curr_guesses\[40\] net93 net78 net476 vssd1 vssd1 vccd1 vccd1 hostdisp.next_curr_guesses\[32\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_106_71 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3422__CLK clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_174_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_106 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2928_ dispFSM.guesses\[68\] net83 net58 net478 vssd1 vssd1 vccd1 vccd1 _0295_ sky130_fd_sc_hd__o22a_1
XFILLER_0_134_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2859_ net66 _1386_ vssd1 vssd1 vccd1 vccd1 _0231_ sky130_fd_sc_hd__and2_1
XANTENNA__1991__Y _0824_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_170_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold241 dispFSM.guesses\[44\] vssd1 vssd1 vccd1 vccd1 net505 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold252 hostdisp.curr_guesses\[11\] vssd1 vssd1 vccd1 vccd1 net516 sky130_fd_sc_hd__dlygate4sd3_1
Xhold230 hostdisp.curr_guesses\[10\] vssd1 vssd1 vccd1 vccd1 net494 sky130_fd_sc_hd__dlygate4sd3_1
Xhold274 hostdisp.curr_guesses\[16\] vssd1 vssd1 vccd1 vccd1 net538 sky130_fd_sc_hd__dlygate4sd3_1
Xhold285 dispFSM.guesses\[25\] vssd1 vssd1 vccd1 vccd1 net549 sky130_fd_sc_hd__dlygate4sd3_1
Xhold263 hostdisp.curr_guesses\[42\] vssd1 vssd1 vccd1 vccd1 net527 sky130_fd_sc_hd__dlygate4sd3_1
Xhold296 hostdisp.curr_word\[15\] vssd1 vssd1 vccd1 vccd1 net560 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_33_clk_X clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2659__A1 net105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_2_3__f_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2595__B1 net108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_150 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2503__B net139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1406__Y _0360_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3445__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2518__X _1096_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2822__A1 _0827_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_256 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2413__B net95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2713_ gamelogic.indexCorrect\[2\] _1276_ _1236_ vssd1 vssd1 vccd1 vccd1 _0195_ sky130_fd_sc_hd__o21a_1
X_2644_ net108 _1215_ _1208_ _1065_ _1214_ vssd1 vssd1 vccd1 vccd1 _1216_ sky130_fd_sc_hd__a2111o_1
X_2575_ dispFSM.guesses\[19\] net105 net111 dispFSM.guesses\[43\] _1149_ vssd1 vssd1
+ vccd1 vccd1 _1150_ sky130_fd_sc_hd__a221o_1
X_1526_ net148 net154 keypadFSMPlayer.prev_key\[1\] vssd1 vssd1 vccd1 vccd1 _0474_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_10_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1457_ hostdisp.curr_word\[29\] vssd1 vssd1 vccd1 vccd1 _0410_ sky130_fd_sc_hd__inv_2
XFILLER_0_184_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3127_ clknet_leaf_18_clk uart_transmitter.next_clk_count\[7\] net219 vssd1 vssd1
+ vccd1 vccd1 uart_transmitter.clk_count\[7\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__2510__B1 net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3058_ clknet_leaf_16_clk _0051_ _0020_ vssd1 vssd1 vccd1 vccd1 keypadFSMPlayer.prev_key\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_117_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_38_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2009_ hostdisp.curr_guesses\[23\] _0823_ net80 net381 vssd1 vssd1 vccd1 vccd1 hostdisp.next_curr_guesses\[15\]
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_120_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_172_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2577__B1 net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_267 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2041__A2 net95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_312 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3318__CLK clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3468__CLK clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3606__240 vssd1 vssd1 vccd1 vccd1 _3606__240/HI net240 sky130_fd_sc_hd__conb_1
XANTENNA_clkbuf_leaf_13_clk_A clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1607__A2 net6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_28_clk_A clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2568__B1 _1097_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3613__244 vssd1 vssd1 vccd1 vccd1 _3613__244/HI net244 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_190_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2032__A2 net94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2520__Y _1098_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2360_ net370 _0997_ net167 vssd1 vssd1 vccd1 vccd1 _0999_ sky130_fd_sc_hd__o21ai_1
X_2291_ _0749_ _0956_ _0958_ vssd1 vssd1 vccd1 vccd1 _0084_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_10_Right_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_139_Right_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_188_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_188_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2559__B1 _1084_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2023__A2 _0823_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2711__X _1275_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout117_A net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2627_ _1096_ _1187_ _1191_ _1097_ _1189_ vssd1 vssd1 vccd1 vccd1 _1200_ sky130_fd_sc_hd__a221o_1
XFILLER_0_88_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2558_ dispFSM.guesses\[10\] _1078_ net105 dispFSM.guesses\[18\] vssd1 vssd1 vccd1
+ vccd1 _1134_ sky130_fd_sc_hd__a22o_1
X_1509_ _0416_ _0435_ _0458_ vssd1 vssd1 vccd1 vccd1 _0459_ sky130_fd_sc_hd__a21o_1
XFILLER_0_10_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2489_ net181 _1067_ vssd1 vssd1 vccd1 vccd1 _0173_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_106_Right_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_167_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_35_clk clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_35_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_182_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2014__A2 net92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2970__B1 net50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_26_clk clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_26_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_68_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1860_ clock_div.count\[28\] _0729_ vssd1 vssd1 vccd1 vccd1 _0730_ sky130_fd_sc_hd__nor2_1
XFILLER_0_140_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1791_ clock_div.count\[1\] clock_div.count\[0\] clock_div.count\[3\] clock_div.count\[5\]
+ vssd1 vssd1 vccd1 vccd1 _0689_ sky130_fd_sc_hd__or4b_1
XFILLER_0_24_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2005__A2 net92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_181_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3530_ clknet_leaf_6_clk hostdisp.next_curr_guesses\[12\] net176 vssd1 vssd1 vccd1
+ vccd1 hostdisp.curr_guesses\[12\] sky130_fd_sc_hd__dfstp_1
XANTENNA__2961__B1 net49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3461_ clknet_leaf_14_clk _0339_ net193 vssd1 vssd1 vccd1 vccd1 gamelogic.setWord\[23\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_149_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3392_ clknet_leaf_20_clk _0281_ net203 vssd1 vssd1 vccd1 vccd1 dispFSM.guesses\[46\]
+ sky130_fd_sc_hd__dfstp_1
X_2412_ net102 net92 vssd1 vssd1 vccd1 vccd1 _1032_ sky130_fd_sc_hd__nor2_1
XFILLER_0_58_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2343_ net150 _0621_ _0990_ vssd1 vssd1 vccd1 vccd1 _0104_ sky130_fd_sc_hd__o21a_1
X_2274_ lcdPlayer.cnt_20ms\[1\] lcdPlayer.cnt_20ms\[0\] vssd1 vssd1 vccd1 vccd1 _0943_
+ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_108_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_9_Left_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_304 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_17_clk clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_17_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__3163__CLK clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1993__A net97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1989_ _0816_ _0820_ vssd1 vssd1 vccd1 vccd1 _0822_ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_167_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3506__CLK clknet_leaf_31_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_167_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_54_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_178_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2999__A net221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3186__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_158_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2526__X _1104_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2961_ gamelogic.setWord\[0\] net53 net49 gamelogic.setWord\[8\] vssd1 vssd1 vccd1
+ vccd1 _0324_ sky130_fd_sc_hd__o22a_1
XFILLER_0_29_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1912_ lcdPlayer.currentState\[0\] net139 net106 vssd1 vssd1 vccd1 vccd1 _0765_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_89 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2892_ dispFSM.guesses\[32\] net81 net56 net546 vssd1 vssd1 vccd1 vccd1 _0259_ sky130_fd_sc_hd__o22a_1
X_1843_ clock_div.count\[20\] _0719_ net488 vssd1 vssd1 vccd1 vccd1 _0720_ sky130_fd_sc_hd__a21oi_1
X_1774_ message_reg.msg\[0\] message_reg.msg\[1\] uart_transmitter.bit_index\[0\]
+ vssd1 vssd1 vccd1 vccd1 _0673_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_155_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3513_ clknet_leaf_31_clk hostdisp.next_curr_word\[35\] net165 vssd1 vssd1 vccd1
+ vccd1 hostdisp.curr_word\[35\] sky130_fd_sc_hd__dfstp_1
X_3444_ clknet_leaf_14_clk _0322_ net193 vssd1 vssd1 vccd1 vccd1 gamelogic.setWord\[6\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_122_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_6_clk clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_6_clk
+ sky130_fd_sc_hd__clkbuf_8
X_3375_ clknet_leaf_21_clk net435 net204 vssd1 vssd1 vccd1 vccd1 dispFSM.guesses\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkload19_A clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_191_Right_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_176_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2326_ lcdPlayer.cnt_500hz\[15\] lcdPlayer.cnt_500hz\[14\] _0977_ vssd1 vssd1 vccd1
+ vccd1 _0980_ sky130_fd_sc_hd__and3_1
XANTENNA__3529__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2257_ net279 buffer.temp_guess\[3\] net127 vssd1 vssd1 vccd1 vccd1 _0070_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout184_A net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_192_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2188_ gamelogic.setWord\[28\] _0896_ net132 vssd1 vssd1 vccd1 vccd1 hostdisp.nextBottom\[76\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_189_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_104 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_51_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_168 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3025__RESET_B net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout97_A _0626_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout52_X net52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_187_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1490_ _0430_ _0440_ _0426_ vssd1 vssd1 vccd1 vccd1 _0442_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_39_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3160_ clknet_leaf_32_clk _0136_ net163 vssd1 vssd1 vccd1 vccd1 hostdisp.top\[44\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1 keypadFSMPlayer.strobe vssd1 vssd1 vccd1 vccd1 net265 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_146_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3091_ clknet_leaf_19_clk _0081_ net211 vssd1 vssd1 vccd1 vccd1 message_reg.msg\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_2111_ hostdisp.curr_word\[39\] net96 _0856_ net140 vssd1 vssd1 vccd1 vccd1 hostdisp.next_curr_word\[39\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__2695__A2 _1259_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_78 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2042_ gamelogic.correct\[1\] gamelogic.correct\[2\] gamelogic.correct\[0\] vssd1
+ vssd1 vccd1 vccd1 _0827_ sky130_fd_sc_hd__and3b_4
XTAP_TAPCELL_ROW_105_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_8_Right_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_115 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2944_ dispFSM.msg\[4\] net84 net58 net473 vssd1 vssd1 vccd1 vccd1 _0311_ sky130_fd_sc_hd__o22a_1
XFILLER_0_17_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2875_ dispFSM.guesses\[15\] net89 net65 net315 vssd1 vssd1 vccd1 vccd1 _0242_ sky130_fd_sc_hd__a22o_1
XFILLER_0_17_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1826_ clock_div.count\[13\] _0709_ net564 vssd1 vssd1 vccd1 vccd1 _0710_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_13_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1757_ uart_receiver.clk_count\[10\] _0658_ _0641_ vssd1 vssd1 vccd1 vccd1 _0660_
+ sky130_fd_sc_hd__a21boi_1
X_1688_ _0607_ _0610_ vssd1 vssd1 vccd1 vccd1 _0611_ sky130_fd_sc_hd__or2_1
XANTENNA__3351__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1990__B _0822_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_39_Right_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3427_ clknet_leaf_29_clk _0001_ vssd1 vssd1 vccd1 vccd1 lcdPlayer.nextState\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_3358_ clknet_leaf_24_clk _0247_ net188 vssd1 vssd1 vccd1 vccd1 dispFSM.guesses\[12\]
+ sky130_fd_sc_hd__dfstp_1
X_2309_ lcdPlayer.cnt_500hz\[9\] _0967_ vssd1 vssd1 vccd1 vccd1 _0969_ sky130_fd_sc_hd__and2_1
X_3289_ clknet_leaf_30_clk hostdisp.nextBottom\[87\] net185 vssd1 vssd1 vccd1 vccd1
+ hostdisp.bottom\[87\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__2438__A2 host_message_reg.setLetter\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_48_Right_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_175_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_7_clk_X clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2610__A2 net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_160_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_95_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_57_Right_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3568__252 vssd1 vssd1 vccd1 vccd1 net252 _3568__252/LO sky130_fd_sc_hd__conb_1
XANTENNA__2488__S _0764_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1899__Y _0752_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1421__A net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_62_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_66_Right_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_168_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_193_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2062__B1 net75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_193_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_100_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2660_ _0760_ _1065_ _1222_ _1228_ _1230_ vssd1 vssd1 vccd1 vccd1 _1231_ sky130_fd_sc_hd__a221o_1
X_1611_ _0542_ _0545_ vssd1 vssd1 vccd1 vccd1 _0546_ sky130_fd_sc_hd__or2_2
XFILLER_0_124_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3374__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2591_ hostdisp.top\[52\] _1097_ _1162_ _1164_ vssd1 vssd1 vccd1 vccd1 _1165_ sky130_fd_sc_hd__a211o_1
XPHY_EDGE_ROW_75_Right_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1542_ _0374_ _0483_ _0488_ vssd1 vssd1 vccd1 vccd1 _0490_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_152_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1473_ _0418_ net128 vssd1 vssd1 vccd1 vccd1 _0425_ sky130_fd_sc_hd__nand2_1
XFILLER_0_1_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3212_ clknet_leaf_11_clk _0188_ net216 vssd1 vssd1 vccd1 vccd1 keypadFSMHost.strobe
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_157_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_111_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3143_ clknet_leaf_26_clk _0119_ vssd1 vssd1 vccd1 vccd1 lcdPlayer.cnt_20ms\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_3074_ clknet_leaf_17_clk keypadFSMPlayer.next_state\[1\] _0036_ vssd1 vssd1 vccd1
+ vccd1 _1400_ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_84_Right_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2025_ net393 net95 net80 net433 vssd1 vssd1 vccd1 vccd1 hostdisp.next_curr_guesses\[31\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_49_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2927_ dispFSM.guesses\[67\] net82 net56 net479 vssd1 vssd1 vccd1 vccd1 _0294_ sky130_fd_sc_hd__o22a_1
XFILLER_0_93_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2858_ net142 buffer.temp_guess\[4\] _0918_ vssd1 vssd1 vccd1 vccd1 _1386_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_93_Right_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1809_ net288 _0698_ vssd1 vssd1 vccd1 vccd1 clock_div.next_count\[6\] sky130_fd_sc_hd__xnor2_1
X_2789_ _0565_ _1288_ vssd1 vssd1 vccd1 vccd1 _1337_ sky130_fd_sc_hd__nor2_1
Xhold220 hostdisp.curr_guesses\[24\] vssd1 vssd1 vccd1 vccd1 net484 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_170_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold231 dispFSM.guesses\[78\] vssd1 vssd1 vccd1 vccd1 net495 sky130_fd_sc_hd__dlygate4sd3_1
Xhold253 hostdisp.curr_guesses\[46\] vssd1 vssd1 vccd1 vccd1 net517 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold242 dispFSM.guesses\[51\] vssd1 vssd1 vccd1 vccd1 net506 sky130_fd_sc_hd__dlygate4sd3_1
Xhold286 dispFSM.guesses\[50\] vssd1 vssd1 vccd1 vccd1 net550 sky130_fd_sc_hd__dlygate4sd3_1
Xhold264 dispFSM.guesses\[27\] vssd1 vssd1 vccd1 vccd1 net528 sky130_fd_sc_hd__dlygate4sd3_1
Xhold275 dispFSM.guesses\[32\] vssd1 vssd1 vccd1 vccd1 net539 sky130_fd_sc_hd__dlygate4sd3_1
Xhold297 lcdPlayer.cnt_500hz\[14\] vssd1 vssd1 vccd1 vccd1 net561 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2108__B2 net142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_0_Left_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3247__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_16_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_140_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_24_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2595__B2 dispFSM.msg\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_376 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_171_202 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2712_ _0926_ _1275_ vssd1 vssd1 vccd1 vccd1 _1276_ sky130_fd_sc_hd__and2b_1
XANTENNA__2586__A1 _0360_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2643_ hostdisp.top\[62\] dispFSM.msg\[6\] net227 vssd1 vssd1 vccd1 vccd1 _1215_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2574_ dispFSM.guesses\[67\] _1072_ _1078_ dispFSM.guesses\[11\] vssd1 vssd1 vccd1
+ vccd1 _1149_ sky130_fd_sc_hd__a22o_1
X_1525_ keypadFSMPlayer.prev_key\[1\] net148 net154 vssd1 vssd1 vccd1 vccd1 _0473_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_10_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1456_ hostdisp.curr_word\[23\] vssd1 vssd1 vccd1 vccd1 _0409_ sky130_fd_sc_hd__inv_2
XFILLER_0_184_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3126_ clknet_leaf_18_clk uart_transmitter.next_clk_count\[6\] net220 vssd1 vssd1
+ vccd1 vccd1 uart_transmitter.clk_count\[6\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_179_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3057_ clknet_leaf_16_clk net333 _0019_ vssd1 vssd1 vccd1 vccd1 keypadFSMPlayer.prev_key\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_38_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2008_ hostdisp.curr_guesses\[22\] net94 net79 hostdisp.curr_guesses\[14\] vssd1
+ vssd1 vccd1 vccd1 hostdisp.next_curr_guesses\[14\] sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_120_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_21_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_172_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_279 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_324 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_45_Left_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_185_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2017__B1 net80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_193_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_54_Left_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_190_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3412__CLK clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2290_ lcdPlayer.cnt_500hz\[0\] lcdPlayer.cnt_500hz\[1\] vssd1 vssd1 vccd1 vccd1
+ _0958_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_63_Left_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_160_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2705__A net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_191_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2008__B1 net79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_72_Left_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2424__B _0827_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_268 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2626_ net113 _1193_ _1198_ _1190_ vssd1 vssd1 vccd1 vccd1 _1199_ sky130_fd_sc_hd__a211o_1
XFILLER_0_2_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3092__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_81_Left_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2557_ dispFSM.guesses\[26\] net114 _1086_ dispFSM.guesses\[74\] vssd1 vssd1 vccd1
+ vccd1 _1133_ sky130_fd_sc_hd__a22o_1
X_1508_ net148 _0415_ net154 _0429_ vssd1 vssd1 vccd1 vccd1 _0458_ sky130_fd_sc_hd__o211ai_1
X_2488_ _1066_ lcdPlayer.lcd_rs _0764_ vssd1 vssd1 vccd1 vccd1 _1067_ sky130_fd_sc_hd__mux2_1
X_1439_ gamelogic.setWord\[9\] vssd1 vssd1 vccd1 vccd1 _0393_ sky130_fd_sc_hd__inv_2
X_3109_ clknet_leaf_28_clk _0099_ vssd1 vssd1 vccd1 vccd1 lcdPlayer.cnt_500hz\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_167_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_167_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_90_Left_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_175_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_166 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3219__Q gamelogic.indexCorrect\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2722__A1 net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1790_ clock_div.count\[11\] clock_div.count\[13\] clock_div.count\[12\] clock_div.count\[10\]
+ vssd1 vssd1 vccd1 vccd1 _0688_ sky130_fd_sc_hd__or4b_1
XFILLER_0_181_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_141_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_172_Right_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3460_ clknet_leaf_5_clk _0338_ net191 vssd1 vssd1 vccd1 vccd1 gamelogic.setWord\[22\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_149_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3391_ clknet_leaf_22_clk _0280_ net202 vssd1 vssd1 vccd1 vccd1 dispFSM.guesses\[45\]
+ sky130_fd_sc_hd__dfrtp_1
X_2411_ _0828_ net123 vssd1 vssd1 vccd1 vccd1 _1031_ sky130_fd_sc_hd__nand2_2
X_2342_ net150 _0621_ _0619_ vssd1 vssd1 vccd1 vccd1 _0990_ sky130_fd_sc_hd__a21oi_1
XANTENNA__2713__A1 gamelogic.indexCorrect\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2273_ dispFSM.msg\[7\] _0941_ _0942_ net324 vssd1 vssd1 vccd1 vccd1 _0082_ sky130_fd_sc_hd__a22o_1
XFILLER_0_165_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_165_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_316 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_191_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_172_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_12_clk_A clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout227_A net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2401__B1 _0017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1988_ _0816_ _0820_ vssd1 vssd1 vccd1 vccd1 _0821_ sky130_fd_sc_hd__nor2_2
XFILLER_0_130_60 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2609_ lcdPlayer.nextState\[3\] hostdisp.bottom\[101\] _1061_ _1069_ vssd1 vssd1
+ vccd1 vccd1 _1182_ sky130_fd_sc_hd__and4b_1
X_3589_ net261 vssd1 vssd1 vccd1 vccd1 gpio_oeb[22] sky130_fd_sc_hd__buf_2
XANTENNA_clkbuf_leaf_27_clk_A clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_2_2__f_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_2_2__leaf_clk sky130_fd_sc_hd__clkbuf_16
XPHY_EDGE_ROW_119_Left_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_126_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_178_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2640__B1 net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_128_Left_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2943__A1 dispFSM.msg\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1424__A net144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_137_Left_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout190 net225 vssd1 vssd1 vccd1 vccd1 net190 sky130_fd_sc_hd__buf_2
XFILLER_0_135_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkload5_A clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2960_ host_message_reg.setLetter\[7\] net55 _1394_ gamelogic.setWord\[7\] vssd1
+ vssd1 vccd1 vccd1 _0323_ sky130_fd_sc_hd__a22o_1
XFILLER_0_139_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2891_ dispFSM.guesses\[31\] net88 net65 net406 vssd1 vssd1 vccd1 vccd1 _0258_ sky130_fd_sc_hd__a22o_1
XANTENNA__2631__B1 net110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1911_ lcdPlayer.cnt_500hz\[13\] _0752_ _0754_ _0763_ vssd1 vssd1 vccd1 vccd1 _0764_
+ sky130_fd_sc_hd__or4_4
XFILLER_0_173_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1842_ net411 _0719_ vssd1 vssd1 vccd1 vccd1 clock_div.next_count\[20\] sky130_fd_sc_hd__xor2_1
XFILLER_0_56_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_146_Left_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1773_ uart_transmitter.bit_index\[2\] _0665_ _0669_ _0672_ vssd1 vssd1 vccd1 vccd1
+ uart_transmitter.next_state\[2\] sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_155_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3512_ clknet_leaf_31_clk hostdisp.next_curr_word\[34\] net165 vssd1 vssd1 vccd1
+ vccd1 hostdisp.curr_word\[34\] sky130_fd_sc_hd__dfstp_1
XFILLER_0_69_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3443_ clknet_leaf_13_clk _0321_ net207 vssd1 vssd1 vccd1 vccd1 gamelogic.setWord\[5\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__3324__RESET_B net218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_114_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3374_ clknet_leaf_21_clk _0263_ net203 vssd1 vssd1 vccd1 vccd1 dispFSM.guesses\[28\]
+ sky130_fd_sc_hd__dfstp_1
X_2325_ net561 _0977_ _0979_ vssd1 vssd1 vccd1 vccd1 _0097_ sky130_fd_sc_hd__o21a_1
XFILLER_0_85_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2256_ net300 buffer.temp_guess\[2\] net127 vssd1 vssd1 vccd1 vccd1 _0069_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_192_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout177_A net179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2187_ gamelogic.setWord\[36\] hostdisp.curr_guesses\[36\] net123 vssd1 vssd1 vccd1
+ vccd1 _0896_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_189_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3280__CLK clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_164_116 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout132_X net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_8_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3232__Q host_message_reg.setLetter\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2208__A3 net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_291 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2803__A gamelogic.letter\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_146_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold2 keypadFSMHost.strobe vssd1 vssd1 vccd1 vccd1 net266 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_146_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3090_ clknet_leaf_21_clk _0080_ net211 vssd1 vssd1 vccd1 vccd1 message_reg.msg\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_2110_ hostdisp.curr_word\[38\] net99 _0855_ gamelogic.letter\[6\] vssd1 vssd1 vccd1
+ vccd1 hostdisp.next_curr_word\[38\] sky130_fd_sc_hd__o22a_1
X_2041_ net140 net95 net80 net428 vssd1 vssd1 vccd1 vccd1 hostdisp.next_curr_guesses\[47\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_55_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2852__A0 net144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_146_127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2943_ dispFSM.msg\[3\] net84 net58 net501 vssd1 vssd1 vccd1 vccd1 _0310_ sky130_fd_sc_hd__o22a_1
XFILLER_0_139_190 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_283 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2874_ dispFSM.guesses\[14\] net85 net60 net413 vssd1 vssd1 vccd1 vccd1 _0241_ sky130_fd_sc_hd__o22a_1
XANTENNA__2080__B2 gamelogic.letter\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1825_ net455 _0709_ vssd1 vssd1 vccd1 vccd1 clock_div.next_count\[13\] sky130_fd_sc_hd__xor2_1
XFILLER_0_25_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2432__B net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1756_ _0658_ _0659_ vssd1 vssd1 vccd1 vccd1 uart_receiver.next_clk_count\[9\] sky130_fd_sc_hd__nor2_1
XFILLER_0_4_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1687_ keypadFSMHost.state\[4\] keypadFSMHost.state\[0\] _0608_ _0609_ _0597_ vssd1
+ vssd1 vccd1 vccd1 _0610_ sky130_fd_sc_hd__o32a_1
X_3426_ clknet_leaf_29_clk _0000_ vssd1 vssd1 vccd1 vccd1 lcdPlayer.nextState\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_96_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3357_ clknet_leaf_25_clk _0246_ net183 vssd1 vssd1 vccd1 vccd1 dispFSM.guesses\[11\]
+ sky130_fd_sc_hd__dfstp_1
X_2308_ lcdPlayer.cnt_500hz\[8\] _0965_ _0968_ vssd1 vssd1 vccd1 vccd1 _0091_ sky130_fd_sc_hd__o21a_1
X_3288_ clknet_leaf_6_clk hostdisp.nextBottom\[86\] net192 vssd1 vssd1 vccd1 vccd1
+ hostdisp.bottom\[86\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_136_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2239_ lcdPlayer.cnt_500hz\[4\] _0755_ lcdPlayer.cnt_500hz\[10\] lcdPlayer.cnt_500hz\[9\]
+ lcdPlayer.cnt_500hz\[8\] vssd1 vssd1 vccd1 vccd1 _0931_ sky130_fd_sc_hd__o2111a_1
XTAP_TAPCELL_ROW_123_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_330 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_175_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2071__B2 gamelogic.letter\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_160_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3176__CLK clknet_leaf_30_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_27_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_70_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_193_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_193_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1610_ net4 net3 net229 vssd1 vssd1 vccd1 vccd1 _0545_ sky130_fd_sc_hd__o21ba_2
X_2590_ hostdisp.bottom\[84\] net118 _1095_ hostdisp.top\[76\] _1163_ vssd1 vssd1
+ vccd1 vccd1 _1164_ sky130_fd_sc_hd__a221o_1
XFILLER_0_1_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1541_ _0483_ _0488_ vssd1 vssd1 vccd1 vccd1 _0489_ sky130_fd_sc_hd__and2_1
XFILLER_0_151_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1472_ net148 keypadplayer.scan_col\[0\] keypadplayer.scan_col\[3\] net147 vssd1
+ vssd1 vccd1 vccd1 _0424_ sky130_fd_sc_hd__or4_1
XFILLER_0_5_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3211_ clknet_leaf_29_clk _0187_ vssd1 vssd1 vccd1 vccd1 lcdPlayer.currentState\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_181_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2522__C1 _1099_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3142_ clknet_leaf_26_clk _0118_ vssd1 vssd1 vccd1 vccd1 lcdPlayer.cnt_20ms\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_78_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3073_ clknet_leaf_17_clk keypadFSMPlayer.next_state\[0\] _0035_ vssd1 vssd1 vccd1
+ vccd1 _1399_ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_163_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2708__A net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1628__A1 net6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2024_ hostdisp.curr_guesses\[38\] net94 net79 net519 vssd1 vssd1 vccd1 vccd1 hostdisp.next_curr_guesses\[30\]
+ sky130_fd_sc_hd__o22a_1
XANTENNA__3049__CLK clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2926_ dispFSM.guesses\[66\] net83 net61 net502 vssd1 vssd1 vccd1 vccd1 _0293_ sky130_fd_sc_hd__o22a_1
XANTENNA__3199__CLK clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2053__B2 net144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2857_ net66 _1385_ vssd1 vssd1 vccd1 vccd1 _0230_ sky130_fd_sc_hd__and2_1
XFILLER_0_72_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1808_ clock_div.count\[4\] clock_div.count\[5\] clock_div.count\[6\] _0696_ vssd1
+ vssd1 vccd1 vccd1 _0700_ sky130_fd_sc_hd__and4_1
XFILLER_0_31_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2788_ host_message_reg.setLetter\[5\] _1336_ net104 vssd1 vssd1 vccd1 vccd1 _0210_
+ sky130_fd_sc_hd__a21o_1
Xhold210 dispFSM.guesses\[67\] vssd1 vssd1 vccd1 vccd1 net474 sky130_fd_sc_hd__dlygate4sd3_1
Xhold221 dispFSM.guesses\[62\] vssd1 vssd1 vccd1 vccd1 net485 sky130_fd_sc_hd__dlygate4sd3_1
Xhold243 dispFSM.guesses\[28\] vssd1 vssd1 vccd1 vccd1 net507 sky130_fd_sc_hd__dlygate4sd3_1
X_1739_ uart_receiver.clk_count\[4\] _0646_ _0641_ vssd1 vssd1 vccd1 vccd1 _0648_
+ sky130_fd_sc_hd__o21ai_1
Xhold232 hostdisp.top\[64\] vssd1 vssd1 vccd1 vccd1 net496 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_170_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold287 hostdisp.curr_guesses\[8\] vssd1 vssd1 vccd1 vccd1 net551 sky130_fd_sc_hd__dlygate4sd3_1
Xhold254 dispFSM.guesses\[22\] vssd1 vssd1 vccd1 vccd1 net518 sky130_fd_sc_hd__dlygate4sd3_1
Xhold276 dispFSM.guesses\[38\] vssd1 vssd1 vccd1 vccd1 net540 sky130_fd_sc_hd__dlygate4sd3_1
Xhold265 dispFSM.guesses\[42\] vssd1 vssd1 vccd1 vccd1 net529 sky130_fd_sc_hd__dlygate4sd3_1
X_3409_ clknet_leaf_21_clk _0298_ net209 vssd1 vssd1 vccd1 vccd1 dispFSM.guesses\[63\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold298 dispFSM.guesses\[14\] vssd1 vssd1 vccd1 vccd1 net562 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2618__A net226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_181_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2595__A2 net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_101_Left_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1432__A net140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_156_222 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3341__CLK clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2035__A1 net144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_119 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2711_ _1266_ _1268_ _1274_ vssd1 vssd1 vccd1 vccd1 _1275_ sky130_fd_sc_hd__and3b_1
XFILLER_0_124_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3491__CLK clknet_leaf_30_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2642_ _1209_ _1211_ _1213_ _0360_ vssd1 vssd1 vccd1 vccd1 _1214_ sky130_fd_sc_hd__o31a_1
XFILLER_0_14_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2573_ dispFSM.guesses\[27\] net114 net109 dispFSM.guesses\[35\] vssd1 vssd1 vccd1
+ vccd1 _1148_ sky130_fd_sc_hd__a22o_1
X_1524_ keypadFSMPlayer.prev_key\[2\] _0460_ vssd1 vssd1 vccd1 vccd1 _0472_ sky130_fd_sc_hd__xor2_1
XFILLER_0_10_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_77 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1455_ hostdisp.curr_word\[21\] vssd1 vssd1 vccd1 vccd1 _0408_ sky130_fd_sc_hd__inv_2
XFILLER_0_10_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3125_ clknet_leaf_18_clk uart_transmitter.next_clk_count\[5\] net220 vssd1 vssd1
+ vccd1 vccd1 uart_transmitter.clk_count\[5\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_6_clk_X clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2510__A2 _1078_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3056_ clknet_leaf_15_clk net265 _0018_ vssd1 vssd1 vccd1 vccd1 keypadFSMPlayer.strobe_edge
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_96_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2007_ net400 net95 net80 net409 vssd1 vssd1 vccd1 vccd1 hostdisp.next_curr_guesses\[13\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_187_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_186_Right_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_82 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2577__A2 net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2909_ dispFSM.guesses\[49\] net87 net62 net526 vssd1 vssd1 vccd1 vccd1 _0276_ sky130_fd_sc_hd__o22a_1
XFILLER_0_5_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_131_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout72_A net73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3364__CLK clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_153_Right_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2568__A2 _1096_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_190_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_49 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_160_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_120 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_203 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_120_Right_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2559__A2 net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2625_ net109 _1186_ _1188_ _1084_ vssd1 vssd1 vccd1 vccd1 _1198_ sky130_fd_sc_hd__a22o_1
XFILLER_0_2_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2556_ dispFSM.guesses\[66\] _1072_ net117 dispFSM.guesses\[58\] vssd1 vssd1 vccd1
+ vccd1 _1132_ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1507_ dispFSM.msg\[6\] _0456_ vssd1 vssd1 vccd1 vccd1 _0457_ sky130_fd_sc_hd__nand2b_1
X_2487_ lcdPlayer.nextState\[3\] _1058_ _1059_ _1064_ net139 vssd1 vssd1 vccd1 vccd1
+ _1066_ sky130_fd_sc_hd__o32a_1
XANTENNA__3387__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1438_ gamelogic.indexCorrect\[0\] vssd1 vssd1 vccd1 vccd1 _0392_ sky130_fd_sc_hd__inv_2
XFILLER_0_179_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3108_ clknet_leaf_28_clk _0098_ vssd1 vssd1 vccd1 vccd1 lcdPlayer.cnt_500hz\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_167_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3039_ clknet_leaf_8_clk clock_div.next_count\[19\] net213 vssd1 vssd1 vccd1 vccd1
+ clock_div.count\[19\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_182_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3235__Q host_message_reg.setLetter\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout75_X net75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_57_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2238__B2 _0607_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_185_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2961__A2 net53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2410_ _0829_ net119 vssd1 vssd1 vccd1 vccd1 _1030_ sky130_fd_sc_hd__nor2_1
XANTENNA__2174__A0 gamelogic.setWord\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3390_ clknet_leaf_23_clk _0279_ net188 vssd1 vssd1 vccd1 vccd1 dispFSM.guesses\[44\]
+ sky130_fd_sc_hd__dfstp_1
X_2341_ net310 _0988_ _0989_ vssd1 vssd1 vccd1 vccd1 _0103_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_149_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2272_ dispFSM.msg\[6\] _0941_ _0942_ net289 vssd1 vssd1 vccd1 vccd1 _0081_ sky130_fd_sc_hd__a22o_1
XANTENNA__1604__B net6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_165_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_108_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_181_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2435__B net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_62 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_370 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1987_ gamelogic.rights\[2\] _0818_ _0819_ vssd1 vssd1 vccd1 vccd1 _0820_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_119_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2608_ dispFSM.guesses\[77\] _1086_ _1178_ _1180_ vssd1 vssd1 vccd1 vccd1 _1181_
+ sky130_fd_sc_hd__a211o_1
X_3588_ net260 vssd1 vssd1 vccd1 vccd1 gpio_oeb[21] sky130_fd_sc_hd__buf_2
X_2539_ dispFSM.guesses\[65\] _1072_ net117 dispFSM.guesses\[57\] vssd1 vssd1 vccd1
+ vccd1 _1116_ sky130_fd_sc_hd__a22o_1
XANTENNA__2704__A2 gamelogic.setWord\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_92 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_126_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_182_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_178_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3402__CLK clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_362 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_31_clk_X clknet_leaf_31_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout191 net192 vssd1 vssd1 vccd1 vccd1 net191 sky130_fd_sc_hd__clkbuf_4
Xfanout180 net190 vssd1 vssd1 vccd1 vccd1 net180 sky130_fd_sc_hd__clkbuf_2
XANTENNA__2459__B2 _0828_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_45_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_146_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3082__CLK clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2890_ dispFSM.guesses\[30\] net85 net62 net518 vssd1 vssd1 vccd1 vccd1 _0257_ sky130_fd_sc_hd__o22a_1
X_1910_ _0755_ _0761_ _0762_ vssd1 vssd1 vccd1 vccd1 _0763_ sky130_fd_sc_hd__or3_1
XFILLER_0_56_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1841_ _0718_ _0719_ vssd1 vssd1 vccd1 vccd1 clock_div.next_count\[19\] sky130_fd_sc_hd__nor2_1
XFILLER_0_56_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_181_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1772_ _0671_ vssd1 vssd1 vccd1 vccd1 _0672_ sky130_fd_sc_hd__inv_2
XFILLER_0_107_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_340 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_155_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3511_ clknet_leaf_32_clk hostdisp.next_curr_word\[33\] net164 vssd1 vssd1 vccd1
+ vccd1 hostdisp.curr_word\[33\] sky130_fd_sc_hd__dfstp_1
X_3442_ clknet_leaf_4_clk _0320_ net194 vssd1 vssd1 vccd1 vccd1 gamelogic.setWord\[4\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_69_67 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3373_ clknet_leaf_25_clk _0262_ net183 vssd1 vssd1 vccd1 vccd1 dispFSM.guesses\[27\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_114_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2324_ net74 _0978_ vssd1 vssd1 vccd1 vccd1 _0979_ sky130_fd_sc_hd__nor2_1
XFILLER_0_40_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_166_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2255_ net326 buffer.temp_guess\[1\] net127 vssd1 vssd1 vccd1 vccd1 _0068_ sky130_fd_sc_hd__mux2_1
X_2186_ gamelogic.setWord\[27\] _0895_ net131 vssd1 vssd1 vccd1 vccd1 hostdisp.nextBottom\[75\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_189_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3425__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_164_128 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2622__A1 net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout125_X net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_180 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_170_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_146_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3 keypadFSMPlayer.strobe_edge vssd1 vssd1 vccd1 vccd1 net267 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3448__CLK clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2040_ gamelogic.letter\[6\] net94 net79 net517 vssd1 vssd1 vccd1 vccd1 hostdisp.next_curr_guesses\[46\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_55_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_11_clk_A clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2942_ dispFSM.msg\[2\] net85 net60 dispFSM.guesses\[74\] vssd1 vssd1 vccd1 vccd1
+ _0309_ sky130_fd_sc_hd__o22a_1
XANTENNA_clkbuf_leaf_26_clk_A clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_146_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2873_ dispFSM.guesses\[13\] net90 net64 net321 vssd1 vssd1 vccd1 vccd1 _0240_ sky130_fd_sc_hd__a22o_1
X_3591__263 vssd1 vssd1 vccd1 vccd1 net263 _3591__263/LO sky130_fd_sc_hd__conb_1
XFILLER_0_84_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1824_ _0708_ _0709_ vssd1 vssd1 vccd1 vccd1 clock_div.next_count\[12\] sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_116_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1755_ uart_receiver.clk_count\[9\] _0656_ _0642_ vssd1 vssd1 vccd1 vccd1 _0659_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_20_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1686_ _0538_ _0601_ vssd1 vssd1 vccd1 vccd1 _0609_ sky130_fd_sc_hd__or2_1
XANTENNA__1591__B2 dispFSM.msg\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3425_ clknet_leaf_21_clk _0314_ net210 vssd1 vssd1 vccd1 vccd1 dispFSM.guesses\[79\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_110_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3356_ clknet_leaf_24_clk _0245_ net187 vssd1 vssd1 vccd1 vccd1 dispFSM.guesses\[10\]
+ sky130_fd_sc_hd__dfstp_1
X_3287_ clknet_leaf_14_clk hostdisp.nextBottom\[85\] net207 vssd1 vssd1 vccd1 vccd1
+ hostdisp.bottom\[85\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__2540__B1 net110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2307_ net74 _0967_ vssd1 vssd1 vccd1 vccd1 _0968_ sky130_fd_sc_hd__nor2_1
XFILLER_0_31_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2238_ _0911_ _0915_ _0930_ _0607_ vssd1 vssd1 vccd1 vccd1 gamelogic.nextState\[3\]
+ sky130_fd_sc_hd__a22o_1
X_2169_ gamelogic.setWord\[27\] hostdisp.curr_guesses\[27\] net121 vssd1 vssd1 vccd1
+ vccd1 _0887_ sky130_fd_sc_hd__mux2_1
XFILLER_0_165_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_175_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_145_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_160_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_134_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_165_Left_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_160_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_95_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_186_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_174_Left_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_183_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2598__B1 net226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_70_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_193_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_193_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_183_Left_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1558__D1 net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1540_ _0472_ _0477_ _0486_ _0487_ vssd1 vssd1 vccd1 vccd1 _0488_ sky130_fd_sc_hd__and4_1
XFILLER_0_151_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1573__A1 dispFSM.msg\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1471_ net148 _0415_ vssd1 vssd1 vccd1 vccd1 _0423_ sky130_fd_sc_hd__nor2_1
XFILLER_0_157_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3270__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3210_ clknet_leaf_29_clk _0186_ vssd1 vssd1 vccd1 vccd1 lcdPlayer.currentState\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__2522__B1 net109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3141_ clknet_leaf_26_clk _0117_ vssd1 vssd1 vccd1 vccd1 lcdPlayer.cnt_20ms\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_174_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_192_Left_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_167_Right_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_163_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3072_ clknet_leaf_21_clk _0065_ _0034_ vssd1 vssd1 vccd1 vccd1 dispFSM.msg\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_173_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2023_ hostdisp.curr_guesses\[37\] _0823_ _0825_ net391 vssd1 vssd1 vccd1 vccd1 hostdisp.next_curr_guesses\[29\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_106_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2589__B1 net109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2925_ dispFSM.guesses\[65\] net86 net63 net530 vssd1 vssd1 vccd1 vccd1 _0292_ sky130_fd_sc_hd__o22a_1
XFILLER_0_17_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2856_ net143 buffer.temp_guess\[3\] _0918_ vssd1 vssd1 vccd1 vccd1 _1385_ sky130_fd_sc_hd__mux2_1
X_1807_ _0693_ _0698_ _0699_ vssd1 vssd1 vccd1 vccd1 clock_div.next_count\[5\] sky130_fd_sc_hd__and3_1
XFILLER_0_31_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2787_ _0609_ _1288_ _0592_ vssd1 vssd1 vccd1 vccd1 _1336_ sky130_fd_sc_hd__a21o_1
Xhold211 hostdisp.curr_guesses\[41\] vssd1 vssd1 vccd1 vccd1 net475 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold200 dispFSM.guesses\[0\] vssd1 vssd1 vccd1 vccd1 net464 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold233 keypadFSMPlayer.prev_key\[6\] vssd1 vssd1 vccd1 vccd1 net497 sky130_fd_sc_hd__dlygate4sd3_1
Xhold244 dispFSM.guesses\[46\] vssd1 vssd1 vccd1 vccd1 net508 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout202_A net206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold222 dispFSM.guesses\[18\] vssd1 vssd1 vccd1 vccd1 net486 sky130_fd_sc_hd__dlygate4sd3_1
X_1738_ _0646_ _0647_ _0642_ vssd1 vssd1 vccd1 vccd1 uart_receiver.next_clk_count\[3\]
+ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_170_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1669_ _0556_ _0559_ vssd1 vssd1 vccd1 vccd1 _0594_ sky130_fd_sc_hd__nor2_1
Xhold277 dispFSM.guesses\[33\] vssd1 vssd1 vccd1 vccd1 net541 sky130_fd_sc_hd__dlygate4sd3_1
Xhold266 dispFSM.guesses\[57\] vssd1 vssd1 vccd1 vccd1 net530 sky130_fd_sc_hd__dlygate4sd3_1
Xhold255 hostdisp.curr_guesses\[30\] vssd1 vssd1 vccd1 vccd1 net519 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold288 gamelogic.setWord\[13\] vssd1 vssd1 vccd1 vccd1 net552 sky130_fd_sc_hd__dlygate4sd3_1
Xhold299 dispFSM.guesses\[49\] vssd1 vssd1 vccd1 vccd1 net563 sky130_fd_sc_hd__dlygate4sd3_1
X_3408_ clknet_leaf_20_clk _0297_ net205 vssd1 vssd1 vccd1 vccd1 dispFSM.guesses\[62\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_0_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input7_A gpio_in[33] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2513__B1 _1086_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3339_ clknet_leaf_33_clk _0228_ net162 vssd1 vssd1 vccd1 vccd1 gamelogic.letter\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_147_92 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_181_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_134_Right_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_84_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_24_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3238__Q host_message_reg.setLetter\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3293__CLK clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_186 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3481__SET_B net164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_101_Right_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_75_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2247__C _0693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_156_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_156_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2440__C1 net71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2710_ _1263_ _1264_ _1270_ _1273_ vssd1 vssd1 vccd1 vccd1 _1274_ sky130_fd_sc_hd__a211oi_1
XANTENNA__2991__B1 net48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2641_ hostdisp.bottom\[46\] net105 net110 hostdisp.bottom\[62\] _1212_ vssd1 vssd1
+ vccd1 vccd1 _1213_ sky130_fd_sc_hd__a221o_1
XFILLER_0_124_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2572_ hostdisp.bottom\[83\] net117 _1142_ _1143_ _1146_ vssd1 vssd1 vccd1 vccd1
+ _1147_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_168_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1523_ _0469_ _0470_ vssd1 vssd1 vccd1 vccd1 _0471_ sky130_fd_sc_hd__nand2_1
XFILLER_0_22_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1454_ hostdisp.curr_word\[15\] vssd1 vssd1 vccd1 vccd1 _0407_ sky130_fd_sc_hd__inv_2
XFILLER_0_77_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3124_ clknet_leaf_18_clk uart_transmitter.next_clk_count\[4\] net220 vssd1 vssd1
+ vccd1 vccd1 uart_transmitter.clk_count\[4\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_179_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3055_ clknet_leaf_15_clk net267 _0017_ vssd1 vssd1 vccd1 vccd1 keypadFSMPlayer.strobe_edge1
+ sky130_fd_sc_hd__dfrtp_1
X_2006_ hostdisp.curr_guesses\[20\] net92 net77 hostdisp.curr_guesses\[12\] vssd1
+ vssd1 vccd1 vccd1 hostdisp.next_curr_guesses\[12\] sky130_fd_sc_hd__o22a_1
XANTENNA__3166__CLK clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_94 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2908_ dispFSM.guesses\[48\] net81 net56 net537 vssd1 vssd1 vccd1 vccd1 _0275_ sky130_fd_sc_hd__o22a_1
XFILLER_0_162_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_21_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2839_ _1370_ _1371_ _1374_ vssd1 vssd1 vccd1 vccd1 _1375_ sky130_fd_sc_hd__and3_1
XFILLER_0_130_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3554__SET_B net179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3509__CLK clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2017__A2 net95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_278 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_190_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3230__RESET_B net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3189__CLK clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_29_clk clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_29_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_188_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_170_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2008__A2 net94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_215 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_179_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2624_ hostdisp.top\[101\] _1177_ _1192_ _1078_ _1196_ vssd1 vssd1 vccd1 vccd1 _1197_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_70_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1905__X _0758_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2555_ _1127_ _1130_ _0360_ vssd1 vssd1 vccd1 vccd1 _1131_ sky130_fd_sc_hd__o21a_1
X_1506_ dispFSM.msg\[7\] _0455_ _0456_ vssd1 vssd1 vccd1 vccd1 _0065_ sky130_fd_sc_hd__and3_1
X_2486_ net106 _1064_ vssd1 vssd1 vccd1 vccd1 _1065_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1437_ gamelogic.setWord\[7\] vssd1 vssd1 vccd1 vccd1 _0391_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_169_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3107_ clknet_leaf_28_clk _0097_ vssd1 vssd1 vccd1 vccd1 lcdPlayer.cnt_500hz\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__3341__Q gamelogic.letter\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3038_ clknet_leaf_8_clk clock_div.next_count\[18\] net214 vssd1 vssd1 vccd1 vccd1
+ clock_div.count\[18\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__2101__D1 gamelogic.indexCorrect\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_190_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2955__B1 net48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3331__CLK clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3251__Q hostdisp.bottom\[49\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_193_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_5_clk_X clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2340_ net310 _0988_ net74 vssd1 vssd1 vccd1 vccd1 _0989_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_58_58 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2271_ dispFSM.msg\[5\] _0941_ _0942_ net352 vssd1 vssd1 vccd1 vccd1 _0080_ sky130_fd_sc_hd__a22o_1
XFILLER_0_165_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_149_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_67 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1986_ gamelogic.rights\[1\] gamelogic.rights\[0\] vssd1 vssd1 vccd1 vccd1 _0819_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_172_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_9_clk clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_9_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_125_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout115_A _1076_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3354__CLK clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2607_ dispFSM.guesses\[21\] _1081_ _1179_ _0360_ vssd1 vssd1 vccd1 vccd1 _1180_
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_61_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3587_ net259 vssd1 vssd1 vccd1 vccd1 gpio_oeb[20] sky130_fd_sc_hd__buf_2
X_2538_ _1112_ _1113_ _1114_ _0360_ vssd1 vssd1 vccd1 vccd1 _1115_ sky130_fd_sc_hd__o31a_1
XFILLER_0_100_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1912__A1 net139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2469_ hostdisp.curr_word\[33\] net72 net69 net312 vssd1 vssd1 vccd1 vccd1 _0165_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_155_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3071__Q dispFSM.msg\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_167_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_54_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_178_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2640__A2 net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_319 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_190_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_374 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_189_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout192 net200 vssd1 vssd1 vccd1 vccd1 net192 sky130_fd_sc_hd__buf_2
Xfanout181 net184 vssd1 vssd1 vccd1 vccd1 net181 sky130_fd_sc_hd__clkbuf_4
XANTENNA__2459__A2 net71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout170 net171 vssd1 vssd1 vccd1 vccd1 net170 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_45_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2631__A2 _1078_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1840_ clock_div.count\[17\] clock_div.count\[19\] clock_div.count\[18\] _0714_ vssd1
+ vssd1 vccd1 vccd1 _0719_ sky130_fd_sc_hd__and4_1
XFILLER_0_154_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3377__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1771_ _0397_ uart_transmitter.state\[0\] uart_transmitter.state\[1\] vssd1 vssd1
+ vccd1 vccd1 _0671_ sky130_fd_sc_hd__or3_1
XFILLER_0_107_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_352 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3510_ clknet_leaf_31_clk hostdisp.next_curr_word\[32\] net164 vssd1 vssd1 vccd1
+ vccd1 hostdisp.curr_word\[32\] sky130_fd_sc_hd__dfstp_1
XFILLER_0_69_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3441_ clknet_leaf_4_clk _0319_ net178 vssd1 vssd1 vccd1 vccd1 gamelogic.setWord\[3\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_69_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3372_ clknet_leaf_24_clk _0261_ net187 vssd1 vssd1 vccd1 vccd1 dispFSM.guesses\[26\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_114_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2323_ lcdPlayer.cnt_500hz\[14\] _0977_ vssd1 vssd1 vccd1 vccd1 _0978_ sky130_fd_sc_hd__and2_1
X_2254_ net317 buffer.temp_guess\[0\] net127 vssd1 vssd1 vccd1 vccd1 _0067_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_166_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2185_ gamelogic.setWord\[35\] hostdisp.curr_guesses\[35\] net121 vssd1 vssd1 vccd1
+ vccd1 _0895_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_69_Left_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_189_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3458__SET_B net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2607__C1 _0360_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2622__A2 hostdisp.bottom\[101\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout232_A net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_310 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1969_ net2 buffer.Rx_byte\[4\] _0805_ vssd1 vssd1 vccd1 vccd1 _0806_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_78_Left_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_160_346 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout118_X net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3066__Q dispFSM.msg\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_184_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_87_Left_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_67_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_183_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_96_Left_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_148_Right_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4 keypadFSMHost.strobe_edge vssd1 vssd1 vccd1 vccd1 net268 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_159_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_186_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_186_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2941_ dispFSM.msg\[1\] net86 net62 net515 vssd1 vssd1 vccd1 vccd1 _0308_ sky130_fd_sc_hd__o22a_1
XFILLER_0_29_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2872_ dispFSM.guesses\[12\] net83 net60 net432 vssd1 vssd1 vccd1 vccd1 _0239_ sky130_fd_sc_hd__o22a_1
X_1823_ clock_div.count\[11\] clock_div.count\[10\] clock_div.count\[12\] _0703_ vssd1
+ vssd1 vccd1 vccd1 _0709_ sky130_fd_sc_hd__and4_1
XFILLER_0_127_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_116_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1754_ uart_receiver.clk_count\[9\] uart_receiver.clk_count\[8\] _0654_ vssd1 vssd1
+ vccd1 vccd1 _0658_ sky130_fd_sc_hd__and3_1
XFILLER_0_40_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1685_ _0538_ _0594_ vssd1 vssd1 vccd1 vccd1 _0608_ sky130_fd_sc_hd__nor2_1
X_3424_ clknet_leaf_20_clk _0313_ net203 vssd1 vssd1 vccd1 vccd1 dispFSM.guesses\[78\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_40_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_115_Right_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3355_ clknet_leaf_21_clk _0244_ net204 vssd1 vssd1 vccd1 vccd1 dispFSM.guesses\[9\]
+ sky130_fd_sc_hd__dfstp_1
X_3286_ clknet_leaf_4_clk hostdisp.nextBottom\[84\] net177 vssd1 vssd1 vccd1 vccd1
+ hostdisp.bottom\[84\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2306_ lcdPlayer.cnt_500hz\[7\] lcdPlayer.cnt_500hz\[8\] _0964_ vssd1 vssd1 vccd1
+ vccd1 _0967_ sky130_fd_sc_hd__and3_1
X_2237_ _0929_ vssd1 vssd1 vccd1 vccd1 _0930_ sky130_fd_sc_hd__inv_2
XFILLER_0_136_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3542__CLK clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2168_ gamelogic.setWord\[18\] _0886_ net131 vssd1 vssd1 vccd1 vccd1 hostdisp.nextBottom\[66\]
+ sky130_fd_sc_hd__mux2_1
X_2099_ hostdisp.curr_word\[36\] hostdisp.curr_word\[38\] _0413_ net99 vssd1 vssd1
+ vccd1 vccd1 _0852_ sky130_fd_sc_hd__a31o_1
XFILLER_0_152_60 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_17_Right_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_30_clk_X clknet_leaf_30_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_160_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_134_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_95_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout95_A _0823_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_186_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3072__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_26_Right_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout50_X net50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_27_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_183_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_35_Right_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_70_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_193_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_255 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2770__A1 host_message_reg.setLetter\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3415__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1470_ _0415_ net154 net148 vssd1 vssd1 vccd1 vccd1 _0422_ sky130_fd_sc_hd__a21o_1
XFILLER_0_157_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_44_Right_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_111_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3140_ clknet_leaf_26_clk _0116_ vssd1 vssd1 vccd1 vccd1 lcdPlayer.cnt_20ms\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_66_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3565__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3071_ clknet_leaf_15_clk _0064_ _0033_ vssd1 vssd1 vccd1 vccd1 dispFSM.msg\[6\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_167_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_163_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2022_ hostdisp.curr_guesses\[36\] net92 net77 net477 vssd1 vssd1 vccd1 vccd1 hostdisp.next_curr_guesses\[28\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_159_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2038__B1 net77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_235 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_122_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_53_Right_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_174_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2924_ dispFSM.guesses\[64\] net82 net56 net513 vssd1 vssd1 vccd1 vccd1 _0291_ sky130_fd_sc_hd__o22a_1
XFILLER_0_127_173 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2855_ net66 _1384_ vssd1 vssd1 vccd1 vccd1 _0229_ sky130_fd_sc_hd__and2_1
X_1806_ clock_div.count\[4\] _0696_ clock_div.count\[5\] vssd1 vssd1 vccd1 vccd1 _0699_
+ sky130_fd_sc_hd__a21o_1
X_2786_ host_message_reg.setLetter\[4\] _1290_ _1310_ _1335_ vssd1 vssd1 vccd1 vccd1
+ _0209_ sky130_fd_sc_hd__o22a_1
Xhold201 hostdisp.curr_guesses\[38\] vssd1 vssd1 vccd1 vccd1 net465 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_115_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold223 hostdisp.curr_guesses\[17\] vssd1 vssd1 vccd1 vccd1 net487 sky130_fd_sc_hd__dlygate4sd3_1
Xhold212 hostdisp.curr_guesses\[32\] vssd1 vssd1 vccd1 vccd1 net476 sky130_fd_sc_hd__dlygate4sd3_1
Xhold234 dispFSM.guesses\[36\] vssd1 vssd1 vccd1 vccd1 net498 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1737_ uart_receiver.clk_count\[1\] uart_receiver.clk_count\[0\] uart_receiver.clk_count\[2\]
+ uart_receiver.clk_count\[3\] vssd1 vssd1 vccd1 vccd1 _0647_ sky130_fd_sc_hd__a31o_1
Xhold267 clock_div.count\[11\] vssd1 vssd1 vccd1 vccd1 net531 sky130_fd_sc_hd__dlygate4sd3_1
X_1668_ keypadFSMHost.state\[1\] keypadFSMHost.state\[5\] keypadFSMHost.state\[2\]
+ keypadFSMHost.state\[3\] vssd1 vssd1 vccd1 vccd1 _0593_ sky130_fd_sc_hd__or4_1
XPHY_EDGE_ROW_62_Right_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold256 lcdPlayer.cnt_20ms\[0\] vssd1 vssd1 vccd1 vccd1 net520 sky130_fd_sc_hd__dlygate4sd3_1
Xhold278 hostdisp.curr_guesses\[35\] vssd1 vssd1 vccd1 vccd1 net542 sky130_fd_sc_hd__dlygate4sd3_1
Xhold245 dispFSM.guesses\[11\] vssd1 vssd1 vccd1 vccd1 net509 sky130_fd_sc_hd__dlygate4sd3_1
X_3407_ clknet_leaf_21_clk _0296_ net201 vssd1 vssd1 vccd1 vccd1 dispFSM.guesses\[61\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold289 hostdisp.curr_guesses\[36\] vssd1 vssd1 vccd1 vccd1 net553 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3344__Q gamelogic.letter\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1599_ net377 net147 _0535_ vssd1 vssd1 vccd1 vccd1 _0052_ sky130_fd_sc_hd__mux2_1
X_3338_ clknet_leaf_33_clk _0227_ net163 vssd1 vssd1 vccd1 vccd1 gamelogic.letter\[0\]
+ sky130_fd_sc_hd__dfrtp_4
X_3269_ clknet_leaf_0_clk hostdisp.nextBottom\[67\] net170 vssd1 vssd1 vccd1 vccd1
+ hostdisp.bottom\[67\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_181_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_71_Right_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3514__SET_B net165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_10_clk_A clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_198 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_80_Right_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_25_clk_A clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_75_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_102_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2640_ hostdisp.bottom\[86\] net118 net112 hostdisp.bottom\[78\] vssd1 vssd1 vccd1
+ vccd1 _1212_ sky130_fd_sc_hd__a22o_1
XFILLER_0_109_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1447__Y _0017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2571_ hostdisp.bottom\[43\] net105 _1144_ _1145_ vssd1 vssd1 vccd1 vccd1 _1146_
+ sky130_fd_sc_hd__a211o_1
X_1522_ keypadFSMPlayer.state\[5\] keypadFSMPlayer.state\[4\] keypadFSMPlayer.state\[1\]
+ _1400_ vssd1 vssd1 vccd1 vccd1 _0470_ sky130_fd_sc_hd__or4b_1
X_1453_ hostdisp.curr_word\[13\] vssd1 vssd1 vccd1 vccd1 _0406_ sky130_fd_sc_hd__inv_2
XANTENNA__3177__RESET_B net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3123_ clknet_leaf_18_clk uart_transmitter.next_clk_count\[3\] net220 vssd1 vssd1
+ vccd1 vccd1 uart_transmitter.clk_count\[3\] sky130_fd_sc_hd__dfrtp_1
X_3054_ clknet_leaf_11_clk _0049_ net216 vssd1 vssd1 vccd1 vccd1 keypadHostt.scan_col\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_179_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2005_ hostdisp.curr_guesses\[19\] net92 net77 net516 vssd1 vssd1 vccd1 vccd1 hostdisp.next_curr_guesses\[11\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_89_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_187_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2454__B net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout145_A gamelogic.letter\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2907_ net384 net88 net65 dispFSM.guesses\[39\] vssd1 vssd1 vccd1 vccd1 _0274_ sky130_fd_sc_hd__a22o_1
XANTENNA__3339__Q gamelogic.letter\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2431__B1 net67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2982__A1 gamelogic.setWord\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2982__B2 gamelogic.setWord\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2838_ gamelogic.correct\[2\] gamelogic.rights\[2\] vssd1 vssd1 vccd1 vccd1 _1374_
+ sky130_fd_sc_hd__xor2_1
X_2769_ host_message_reg.setLetter\[1\] _0601_ _0604_ _1321_ _1310_ vssd1 vssd1 vccd1
+ vccd1 _1322_ sky130_fd_sc_hd__a221o_1
XFILLER_0_130_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_269 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout100_X net100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_29_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_14_Left_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_80_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3260__CLK clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_153_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_260 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_23_Left_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_32_Left_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_169_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_227 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_41_Left_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_271 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2623_ net111 _1194_ _1195_ lcdPlayer.nextState\[4\] vssd1 vssd1 vccd1 vccd1 _1196_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_179_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2716__A1 gamelogic.letter\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2554_ hostdisp.bottom\[50\] net114 net109 hostdisp.bottom\[58\] _1129_ vssd1 vssd1
+ vccd1 vccd1 _1130_ sky130_fd_sc_hd__a221o_1
X_1505_ _0430_ _0440_ keypadFSMPlayer.state\[4\] _0374_ _0426_ vssd1 vssd1 vccd1 vccd1
+ _0456_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_10_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2485_ _1062_ _1063_ vssd1 vssd1 vccd1 vccd1 _1064_ sky130_fd_sc_hd__or2_1
X_1436_ gamelogic.setWord\[0\] vssd1 vssd1 vccd1 vccd1 _0390_ sky130_fd_sc_hd__inv_2
XANTENNA__2449__B net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_169_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3106_ clknet_leaf_27_clk _0096_ vssd1 vssd1 vccd1 vccd1 lcdPlayer.cnt_500hz\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_50_Left_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_179_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3037_ clknet_leaf_8_clk clock_div.next_count\[17\] net213 vssd1 vssd1 vccd1 vccd1
+ clock_div.count\[17\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__3283__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_72 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2652__B1 _1085_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3069__Q dispFSM.msg\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2955__A1 host_message_reg.setLetter\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2404__S _0934_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_57_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_166_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2946__A1 dispFSM.msg\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3156__CLK clknet_leaf_31_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2270_ dispFSM.msg\[4\] _0941_ _0942_ net281 vssd1 vssd1 vccd1 vccd1 _0079_ sky130_fd_sc_hd__a22o_1
XFILLER_0_165_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_181_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2634__B1 net105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_176_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_184_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_172_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1985_ gamelogic.incorrect\[1\] gamelogic.incorrect\[2\] _0817_ vssd1 vssd1 vccd1
+ vccd1 _0818_ sky130_fd_sc_hd__a21o_1
XFILLER_0_172_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2606_ dispFSM.guesses\[29\] net115 net108 dispFSM.msg\[5\] vssd1 vssd1 vccd1 vccd1
+ _1179_ sky130_fd_sc_hd__a22o_1
XANTENNA__3121__RESET_B net223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3586_ net157 vssd1 vssd1 vccd1 vccd1 net16 sky130_fd_sc_hd__clkbuf_1
XANTENNA_fanout108_A _1106_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2537_ hostdisp.top\[73\] _1095_ _1098_ hostdisp.top\[41\] vssd1 vssd1 vccd1 vccd1
+ _1114_ sky130_fd_sc_hd__a22o_1
X_2468_ hostdisp.curr_word\[32\] net72 net68 net330 vssd1 vssd1 vccd1 vccd1 _0164_
+ sky130_fd_sc_hd__a22o_1
X_1419_ keypadFSMPlayer.state\[1\] vssd1 vssd1 vccd1 vccd1 _0373_ sky130_fd_sc_hd__inv_2
X_2399_ lcdPlayer.cnt_20ms\[19\] _1022_ vssd1 vssd1 vccd1 vccd1 _1025_ sky130_fd_sc_hd__nand2_1
XFILLER_0_167_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3029__CLK clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_178_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_148_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_190_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2134__S net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_129_Right_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3179__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_98_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_189_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout80_X net80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout160 net225 vssd1 vssd1 vccd1 vccd1 net160 sky130_fd_sc_hd__buf_2
Xfanout182 net183 vssd1 vssd1 vccd1 vccd1 net182 sky130_fd_sc_hd__buf_2
Xfanout171 net180 vssd1 vssd1 vccd1 vccd1 net171 sky130_fd_sc_hd__buf_2
Xfanout193 net194 vssd1 vssd1 vccd1 vccd1 net193 sky130_fd_sc_hd__clkbuf_4
XANTENNA__2864__A0 net140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_106_Left_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_45_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2616__B1 _1098_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2092__B2 net144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1770_ message_reg.state\[0\] _0670_ _0667_ vssd1 vssd1 vccd1 vccd1 uart_transmitter.next_state\[1\]
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_64_180 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3440_ clknet_leaf_4_clk _0318_ net194 vssd1 vssd1 vccd1 vccd1 gamelogic.setWord\[2\]
+ sky130_fd_sc_hd__dfstp_1
X_3371_ clknet_leaf_20_clk _0260_ net210 vssd1 vssd1 vccd1 vccd1 dispFSM.guesses\[25\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_176_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2322_ _0977_ _0956_ _0976_ vssd1 vssd1 vccd1 vccd1 _0096_ sky130_fd_sc_hd__and3b_1
XFILLER_0_85_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2253_ net285 _0537_ _0605_ vssd1 vssd1 vccd1 vccd1 _0066_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_166_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2184_ gamelogic.setWord\[26\] _0894_ net131 vssd1 vssd1 vccd1 vccd1 hostdisp.nextBottom\[74\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_149_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_125_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2083__B2 net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_157_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_145_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1968_ net149 net150 uart_receiver.bit_index\[2\] vssd1 vssd1 vccd1 vccd1 _0805_
+ sky130_fd_sc_hd__or3b_1
XFILLER_0_43_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout225_A net8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3471__CLK clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1899_ lcdPlayer.cnt_500hz\[4\] _0751_ vssd1 vssd1 vccd1 vccd1 _0752_ sky130_fd_sc_hd__nand2_2
X_3569_ net253 vssd1 vssd1 vccd1 vccd1 gpio_oeb[2] sky130_fd_sc_hd__buf_2
XFILLER_0_11_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_184_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_4_clk_X clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_196 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold5 lcdPlayer.cnt_20ms\[5\] vssd1 vssd1 vccd1 vccd1 net269 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_186_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3344__CLK clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_186_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2065__B2 gamelogic.letter\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2940_ dispFSM.msg\[0\] net84 net58 net521 vssd1 vssd1 vccd1 vccd1 _0307_ sky130_fd_sc_hd__o22a_1
XFILLER_0_29_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2871_ dispFSM.guesses\[11\] net82 net57 net405 vssd1 vssd1 vccd1 vccd1 _0238_ sky130_fd_sc_hd__o22a_1
X_1822_ net468 _0707_ vssd1 vssd1 vccd1 vccd1 _0708_ sky130_fd_sc_hd__nor2_1
XANTENNA__3494__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_128 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1753_ _0656_ _0657_ vssd1 vssd1 vccd1 vccd1 uart_receiver.next_clk_count\[8\] sky130_fd_sc_hd__nor2_1
X_1684_ _0538_ _0598_ vssd1 vssd1 vccd1 vccd1 _0607_ sky130_fd_sc_hd__nor2_2
XFILLER_0_20_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1907__A net139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3423_ clknet_leaf_21_clk _0312_ net202 vssd1 vssd1 vccd1 vccd1 dispFSM.guesses\[77\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_110_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_96_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3354_ clknet_leaf_23_clk _0243_ net182 vssd1 vssd1 vccd1 vccd1 dispFSM.guesses\[8\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__2540__A2 _1086_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2305_ net319 _0964_ _0966_ vssd1 vssd1 vccd1 vccd1 _0090_ sky130_fd_sc_hd__o21a_1
X_3285_ clknet_leaf_30_clk hostdisp.nextBottom\[83\] net184 vssd1 vssd1 vccd1 vccd1
+ hostdisp.bottom\[83\] sky130_fd_sc_hd__dfrtp_1
X_2236_ gamelogic.state\[2\] _0928_ vssd1 vssd1 vccd1 vccd1 _0929_ sky130_fd_sc_hd__or2_1
XFILLER_0_17_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout175_A net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2167_ gamelogic.setWord\[26\] hostdisp.curr_guesses\[26\] net121 vssd1 vssd1 vccd1
+ vccd1 _0886_ sky130_fd_sc_hd__mux2_1
XFILLER_0_177_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2098_ hostdisp.curr_word\[31\] net96 _0851_ net140 vssd1 vssd1 vccd1 vccd1 hostdisp.next_curr_word\[31\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__2056__B2 net142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_192_214 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_72 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout130_X net130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout228_X net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_134_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3217__CLK clknet_leaf_31_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_186_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_203 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_183_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3224__RESET_B net223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_181_Right_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_286 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_10_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2522__A2 net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3070_ clknet_leaf_21_clk _0063_ _0032_ vssd1 vssd1 vccd1 vccd1 dispFSM.msg\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_78_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2021_ hostdisp.curr_guesses\[35\] net91 net76 net472 vssd1 vssd1 vccd1 vccd1 hostdisp.next_curr_guesses\[27\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_159_200 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_18_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2038__A1 net142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2589__A2 net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2923_ dispFSM.guesses\[63\] net88 net65 net425 vssd1 vssd1 vccd1 vccd1 _0290_ sky130_fd_sc_hd__a22o_1
XFILLER_0_122_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2854_ gamelogic.letter\[2\] buffer.temp_guess\[2\] _0918_ vssd1 vssd1 vccd1 vccd1
+ _1384_ sky130_fd_sc_hd__mux2_1
X_1805_ clock_div.count\[4\] clock_div.count\[5\] _0696_ vssd1 vssd1 vccd1 vccd1 _0698_
+ sky130_fd_sc_hd__nand3_1
X_2785_ _1327_ _1331_ _1334_ vssd1 vssd1 vccd1 vccd1 _1335_ sky130_fd_sc_hd__a21o_1
XFILLER_0_127_185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2210__A1 net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold202 dispFSM.guesses\[34\] vssd1 vssd1 vccd1 vccd1 net466 sky130_fd_sc_hd__dlygate4sd3_1
X_1736_ uart_receiver.clk_count\[1\] uart_receiver.clk_count\[0\] uart_receiver.clk_count\[2\]
+ uart_receiver.clk_count\[3\] vssd1 vssd1 vccd1 vccd1 _0646_ sky130_fd_sc_hd__and4_1
Xhold224 clock_div.count\[21\] vssd1 vssd1 vccd1 vccd1 net488 sky130_fd_sc_hd__dlygate4sd3_1
Xhold213 hostdisp.curr_guesses\[28\] vssd1 vssd1 vccd1 vccd1 net477 sky130_fd_sc_hd__dlygate4sd3_1
Xhold235 dispFSM.guesses\[52\] vssd1 vssd1 vccd1 vccd1 net499 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1667_ _0538_ _0564_ vssd1 vssd1 vccd1 vccd1 _0592_ sky130_fd_sc_hd__nor2_1
Xhold268 dispFSM.guesses\[9\] vssd1 vssd1 vccd1 vccd1 net532 sky130_fd_sc_hd__dlygate4sd3_1
Xhold246 dispFSM.guesses\[54\] vssd1 vssd1 vccd1 vccd1 net510 sky130_fd_sc_hd__dlygate4sd3_1
Xhold257 dispFSM.guesses\[72\] vssd1 vssd1 vccd1 vccd1 net521 sky130_fd_sc_hd__dlygate4sd3_1
X_1598_ net342 net146 _0535_ vssd1 vssd1 vccd1 vccd1 _0053_ sky130_fd_sc_hd__mux2_1
Xhold279 dispFSM.guesses\[70\] vssd1 vssd1 vccd1 vccd1 net543 sky130_fd_sc_hd__dlygate4sd3_1
X_3406_ clknet_leaf_23_clk _0295_ net188 vssd1 vssd1 vccd1 vccd1 dispFSM.guesses\[60\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_40_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3337_ clknet_leaf_0_clk _0226_ net171 vssd1 vssd1 vccd1 vccd1 gamelogic.incorrect\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__2513__A2 net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3268_ clknet_leaf_2_clk hostdisp.nextBottom\[66\] net170 vssd1 vssd1 vccd1 vccd1
+ hostdisp.bottom\[66\] sky130_fd_sc_hd__dfrtp_1
X_3199_ clknet_leaf_24_clk _0175_ vssd1 vssd1 vccd1 vccd1 net44 sky130_fd_sc_hd__dfxtp_1
X_2219_ _0913_ _0914_ vssd1 vssd1 vccd1 vccd1 _0915_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_181_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2407__S _0934_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_60 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_24_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2142__S net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1960__A0 net2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2268__A1 dispFSM.msg\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2440__A1 net130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2440__B2 net73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2991__A2 net52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3532__CLK clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2570_ hostdisp.bottom\[67\] net111 net109 hostdisp.bottom\[59\] vssd1 vssd1 vccd1
+ vccd1 _1145_ sky130_fd_sc_hd__a22o_1
XFILLER_0_168_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1521_ keypadFSMPlayer.state\[2\] keypadFSMPlayer.state\[3\] vssd1 vssd1 vccd1 vccd1
+ _0469_ sky130_fd_sc_hd__nor2_1
XFILLER_0_105_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1452_ hostdisp.curr_word\[7\] vssd1 vssd1 vccd1 vccd1 _0405_ sky130_fd_sc_hd__inv_2
XFILLER_0_184_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3122_ clknet_leaf_18_clk uart_transmitter.next_clk_count\[2\] net224 vssd1 vssd1
+ vccd1 vccd1 uart_transmitter.clk_count\[2\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__3520__SET_B net180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3053_ clknet_leaf_11_clk _0048_ net216 vssd1 vssd1 vccd1 vccd1 keypadHostt.scan_col\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_117_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2004_ hostdisp.curr_guesses\[18\] net91 net77 net494 vssd1 vssd1 vccd1 vccd1 hostdisp.next_curr_guesses\[10\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_187_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2906_ dispFSM.guesses\[46\] net87 net61 net540 vssd1 vssd1 vccd1 vccd1 _0273_ sky130_fd_sc_hd__o22a_1
XFILLER_0_9_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2837_ _1373_ gamelogic.correct\[1\] _1366_ vssd1 vssd1 vccd1 vccd1 _0222_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2768_ _1314_ _1320_ _1300_ vssd1 vssd1 vccd1 vccd1 _1321_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_131_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2699_ net140 gamelogic.setWord\[23\] vssd1 vssd1 vccd1 vccd1 _1263_ sky130_fd_sc_hd__nand2_1
X_1719_ uart_receiver.clk_count\[1\] uart_receiver.clk_count\[0\] vssd1 vssd1 vccd1
+ vccd1 _0635_ sky130_fd_sc_hd__or2_1
XFILLER_0_111_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3555__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2600__S net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_17 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_176_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_239 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2177__A0 gamelogic.setWord\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2622_ net228 hostdisp.bottom\[101\] _1070_ _1082_ vssd1 vssd1 vccd1 vccd1 _1195_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_2_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2553_ hostdisp.bottom\[42\] net105 _1097_ hostdisp.top\[50\] _1128_ vssd1 vssd1
+ vccd1 vccd1 _1129_ sky130_fd_sc_hd__a221o_1
X_1504_ _0434_ _0447_ vssd1 vssd1 vccd1 vccd1 _0455_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_189_Left_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2484_ net138 lcdPlayer.nextState\[2\] vssd1 vssd1 vccd1 vccd1 _1063_ sky130_fd_sc_hd__nand2b_1
X_1435_ gamelogic.setWord\[17\] vssd1 vssd1 vccd1 vccd1 _0389_ sky130_fd_sc_hd__inv_2
XFILLER_0_10_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_169_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3105_ clknet_leaf_27_clk _0095_ vssd1 vssd1 vccd1 vccd1 lcdPlayer.cnt_500hz\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__3428__CLK clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3036_ clknet_leaf_8_clk clock_div.next_count\[16\] net213 vssd1 vssd1 vccd1 vccd1
+ clock_div.count\[16\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_179_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2101__B1 net75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2465__B net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_190_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_24_clk_A clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_190_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2955__A2 net52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout70_A net71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2643__A1 dispFSM.msg\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_40_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_165_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_181_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1984_ gamelogic.correct\[0\] gamelogic.correct\[1\] gamelogic.correct\[2\] vssd1
+ vssd1 vccd1 vccd1 _0817_ sky130_fd_sc_hd__o21a_1
XFILLER_0_172_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2605_ dispFSM.guesses\[69\] _1072_ net117 dispFSM.guesses\[61\] _1177_ vssd1 vssd1
+ vccd1 vccd1 _1178_ sky130_fd_sc_hd__a221o_1
XANTENNA__3100__CLK clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3585_ net156 vssd1 vssd1 vccd1 vccd1 net15 sky130_fd_sc_hd__clkbuf_1
X_2536_ hostdisp.bottom\[49\] net114 _1097_ hostdisp.top\[49\] _1110_ vssd1 vssd1
+ vccd1 vccd1 _1113_ sky130_fd_sc_hd__a221o_1
XFILLER_0_2_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3250__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2467_ hostdisp.curr_word\[31\] net73 net68 net415 vssd1 vssd1 vccd1 vccd1 _0163_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__2570__B1 net109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1418_ keypadFSMPlayer.state\[4\] vssd1 vssd1 vccd1 vccd1 _0372_ sky130_fd_sc_hd__inv_2
XFILLER_0_47_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2398_ lcdPlayer.cnt_20ms\[19\] _1022_ vssd1 vssd1 vccd1 vccd1 _1024_ sky130_fd_sc_hd__or2_1
X_3603__237 vssd1 vssd1 vccd1 vccd1 _3603__237/HI net237 sky130_fd_sc_hd__conb_1
XFILLER_0_3_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3019_ net223 vssd1 vssd1 vccd1 vccd1 _0044_ sky130_fd_sc_hd__inv_2
XANTENNA__2625__A1 net109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2625__B2 _1084_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_172 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_228 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_137_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_190_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_189_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3249__RESET_B net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2561__B1 net226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout150 uart_receiver.bit_index\[0\] vssd1 vssd1 vccd1 vccd1 net150 sky130_fd_sc_hd__clkbuf_2
Xfanout161 net162 vssd1 vssd1 vccd1 vccd1 net161 sky130_fd_sc_hd__clkbuf_4
Xfanout183 net184 vssd1 vssd1 vccd1 vccd1 net183 sky130_fd_sc_hd__clkbuf_4
Xfanout172 net174 vssd1 vssd1 vccd1 vccd1 net172 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout73_X net73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout194 net200 vssd1 vssd1 vccd1 vccd1 net194 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_44_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_45_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2616__A1 net226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3010__A net223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3273__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3370_ clknet_leaf_25_clk _0259_ net182 vssd1 vssd1 vccd1 vccd1 dispFSM.guesses\[24\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_176_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2321_ lcdPlayer.cnt_500hz\[13\] lcdPlayer.cnt_500hz\[12\] _0973_ vssd1 vssd1 vccd1
+ vccd1 _0977_ sky130_fd_sc_hd__and3_1
XANTENNA__2552__B1 _1098_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2252_ _0550_ keypadHostt.scan_col\[3\] _0937_ vssd1 vssd1 vccd1 vccd1 _0049_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_166_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2183_ gamelogic.setWord\[34\] hostdisp.curr_guesses\[34\] net121 vssd1 vssd1 vccd1
+ vccd1 _0894_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_125_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2083__A2 net97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_145_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1967_ _0618_ _0804_ vssd1 vssd1 vccd1 vccd1 uart_receiver.temp_byte\[3\] sky130_fd_sc_hd__and2_1
XFILLER_0_50_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout218_A net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1594__A1 net6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1898_ lcdPlayer.cnt_500hz\[3\] _0750_ vssd1 vssd1 vccd1 vccd1 _0751_ sky130_fd_sc_hd__and2_1
XFILLER_0_70_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3568_ net252 vssd1 vssd1 vccd1 vccd1 gpio_oeb[1] sky130_fd_sc_hd__buf_2
XANTENNA__2543__B1 _1084_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2519_ _1060_ _1093_ vssd1 vssd1 vccd1 vccd1 _1097_ sky130_fd_sc_hd__nor2_4
X_3499_ clknet_leaf_14_clk hostdisp.next_curr_word\[21\] net201 vssd1 vssd1 vccd1
+ vccd1 hostdisp.curr_word\[21\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_89_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_91 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_184_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_162_Right_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2145__S net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2534__B1 net109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold6 _0112_ vssd1 vssd1 vccd1 vccd1 net270 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_186_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_162_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2870_ dispFSM.guesses\[10\] net83 net58 net419 vssd1 vssd1 vccd1 vccd1 _0237_ sky130_fd_sc_hd__o22a_1
XANTENNA__2470__C1 _1034_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1821_ _0706_ _0707_ vssd1 vssd1 vccd1 vccd1 clock_div.next_count\[11\] sky130_fd_sc_hd__nor2_1
XFILLER_0_37_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_10_clk clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_10_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_154_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1752_ uart_receiver.clk_count\[8\] _0654_ _0641_ vssd1 vssd1 vccd1 vccd1 _0657_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_187_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1683_ _0582_ _0605_ vssd1 vssd1 vccd1 vccd1 _0606_ sky130_fd_sc_hd__and2_1
XFILLER_0_20_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1907__B net106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3422_ clknet_leaf_23_clk _0311_ net187 vssd1 vssd1 vccd1 vccd1 dispFSM.guesses\[76\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_20_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2525__B1 _1097_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3353_ clknet_leaf_21_clk net316 net204 vssd1 vssd1 vccd1 vccd1 dispFSM.guesses\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2304_ _0957_ _0965_ vssd1 vssd1 vccd1 vccd1 _0966_ sky130_fd_sc_hd__nor2_1
X_3284_ clknet_leaf_2_clk hostdisp.nextBottom\[82\] net170 vssd1 vssd1 vccd1 vccd1
+ hostdisp.bottom\[82\] sky130_fd_sc_hd__dfrtp_1
X_2235_ gamelogic.state\[0\] gamelogic.state\[1\] gamelogic.state\[3\] vssd1 vssd1
+ vccd1 vccd1 _0928_ sky130_fd_sc_hd__or3_1
X_2166_ gamelogic.setWord\[17\] _0885_ net135 vssd1 vssd1 vccd1 vccd1 hostdisp.nextBottom\[65\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3169__CLK clknet_leaf_30_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_177_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout168_A net169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2097_ hostdisp.curr_word\[30\] net101 _0850_ gamelogic.letter\[6\] vssd1 vssd1 vccd1
+ vccd1 hostdisp.next_curr_word\[30\] sky130_fd_sc_hd__o22a_1
XFILLER_0_0_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_226 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_3_Right_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_160_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2999_ net221 vssd1 vssd1 vccd1 vccd1 _0024_ sky130_fd_sc_hd__inv_2
XFILLER_0_133_304 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_125_Left_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_160_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout123_X net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_186_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_134_Left_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_145_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2452__C1 net71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_143_Left_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3616__247 vssd1 vssd1 vccd1 vccd1 _3616__247/HI net247 sky130_fd_sc_hd__conb_1
XFILLER_0_19_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_70_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_191_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_152_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_152_Left_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_111_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3311__CLK clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2020_ hostdisp.curr_guesses\[34\] net91 net76 net548 vssd1 vssd1 vccd1 vccd1 hostdisp.next_curr_guesses\[26\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_173_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3461__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_18_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2038__A2 net92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_161_Left_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_122_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2922_ dispFSM.guesses\[62\] net85 net60 net510 vssd1 vssd1 vccd1 vccd1 _0289_ sky130_fd_sc_hd__o22a_1
XFILLER_0_97_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_61_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2443__C1 net70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2853_ net66 _1383_ vssd1 vssd1 vccd1 vccd1 _0228_ sky130_fd_sc_hd__and2_1
X_1804_ net461 _0696_ vssd1 vssd1 vccd1 vccd1 clock_div.next_count\[4\] sky130_fd_sc_hd__xor2_1
X_2784_ _0541_ _0543_ _0551_ _0601_ host_message_reg.setLetter\[4\] vssd1 vssd1 vccd1
+ vccd1 _1334_ sky130_fd_sc_hd__a32o_1
XANTENNA__3543__SET_B net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_268 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1735_ _0641_ _0644_ _0645_ vssd1 vssd1 vccd1 vccd1 uart_receiver.next_clk_count\[2\]
+ sky130_fd_sc_hd__and3_1
XANTENNA_clkbuf_leaf_3_clk_X clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold203 clock_div.count\[22\] vssd1 vssd1 vccd1 vccd1 net467 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold225 hostdisp.curr_guesses\[20\] vssd1 vssd1 vccd1 vccd1 net489 sky130_fd_sc_hd__dlygate4sd3_1
Xhold214 dispFSM.guesses\[60\] vssd1 vssd1 vccd1 vccd1 net478 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_170_Left_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1666_ _0590_ _0012_ vssd1 vssd1 vccd1 vccd1 keypadFSMPlayer.next_state\[2\] sky130_fd_sc_hd__or2_1
Xhold236 hostdisp.curr_guesses\[22\] vssd1 vssd1 vccd1 vccd1 net500 sky130_fd_sc_hd__dlygate4sd3_1
Xhold247 dispFSM.guesses\[26\] vssd1 vssd1 vccd1 vccd1 net511 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold269 lcdPlayer.cnt_500hz\[1\] vssd1 vssd1 vccd1 vccd1 net533 sky130_fd_sc_hd__dlygate4sd3_1
Xhold258 dispFSM.guesses\[19\] vssd1 vssd1 vccd1 vccd1 net522 sky130_fd_sc_hd__dlygate4sd3_1
X_1597_ net386 _0418_ _0535_ vssd1 vssd1 vccd1 vccd1 _0054_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3405_ clknet_leaf_25_clk _0294_ net184 vssd1 vssd1 vccd1 vccd1 dispFSM.guesses\[59\]
+ sky130_fd_sc_hd__dfstp_1
X_3336_ clknet_leaf_0_clk _0225_ net171 vssd1 vssd1 vccd1 vccd1 gamelogic.incorrect\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_147_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3267_ clknet_leaf_15_clk hostdisp.nextBottom\[65\] net209 vssd1 vssd1 vccd1 vccd1
+ hostdisp.bottom\[65\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_71 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2218_ buffer.temp_guess\[0\] buffer.temp_guess\[1\] buffer.temp_guess\[2\] buffer.temp_guess\[3\]
+ vssd1 vssd1 vccd1 vccd1 _0914_ sky130_fd_sc_hd__or4_1
X_3198_ clknet_leaf_25_clk _0174_ vssd1 vssd1 vccd1 vccd1 net43 sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_181_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2149_ gamelogic.setWord\[17\] hostdisp.curr_guesses\[17\] net125 vssd1 vssd1 vccd1
+ vccd1 _0877_ sky130_fd_sc_hd__mux2_1
XFILLER_0_163_72 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2985__B1 net49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_192_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3484__CLK clknet_leaf_31_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2681__X _1247_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2440__A2 host_message_reg.setLetter\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1520_ net6 _0416_ _0467_ net128 vssd1 vssd1 vccd1 vccd1 _0468_ sky130_fd_sc_hd__or4b_1
XFILLER_0_22_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1451_ hostdisp.curr_word\[5\] vssd1 vssd1 vccd1 vccd1 _0404_ sky130_fd_sc_hd__inv_2
XFILLER_0_184_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3121_ clknet_leaf_18_clk net291 net223 vssd1 vssd1 vccd1 vccd1 uart_transmitter.clk_count\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_172_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3052_ clknet_leaf_11_clk _0047_ net216 vssd1 vssd1 vccd1 vccd1 keypadHostt.scan_col\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_117_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_179_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2003_ hostdisp.curr_guesses\[17\] net94 net79 net457 vssd1 vssd1 vccd1 vccd1 hostdisp.next_curr_guesses\[9\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_26_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2967__B1 net49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2905_ net373 net90 net64 dispFSM.guesses\[37\] vssd1 vssd1 vccd1 vccd1 _0272_ sky130_fd_sc_hd__a22o_1
XANTENNA__2431__A2 _1031_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2836_ _0815_ _1371_ _1372_ vssd1 vssd1 vccd1 vccd1 _1373_ sky130_fd_sc_hd__and3_1
XFILLER_0_170_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2767_ _1312_ _1318_ vssd1 vssd1 vccd1 vccd1 _1320_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_115_178 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout200_A net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1718_ uart_receiver.state\[0\] _0617_ vssd1 vssd1 vccd1 vccd1 _0634_ sky130_fd_sc_hd__or2_1
XFILLER_0_77_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2698_ _1236_ _1262_ vssd1 vssd1 vccd1 vccd1 _0194_ sky130_fd_sc_hd__and2_1
X_1649_ _0541_ _0553_ _0555_ vssd1 vssd1 vccd1 vccd1 _0584_ sky130_fd_sc_hd__and3_1
XANTENNA_input5_A gpio_in[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3319_ clknet_leaf_12_clk _0005_ net215 vssd1 vssd1 vccd1 vccd1 keypadFSMHost.state\[0\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA_fanout190_X net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2110__B2 gamelogic.letter\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_43_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2621_ hostdisp.bottom\[69\] dispFSM.guesses\[45\] net227 vssd1 vssd1 vccd1 vccd1
+ _1194_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2552_ hostdisp.bottom\[66\] net111 _1098_ hostdisp.top\[42\] vssd1 vssd1 vccd1 vccd1
+ _1128_ sky130_fd_sc_hd__a22o_1
X_1503_ _0434_ _0443_ vssd1 vssd1 vccd1 vccd1 _0454_ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_282 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2483_ lcdPlayer.nextState\[3\] _1061_ vssd1 vssd1 vccd1 vccd1 _1062_ sky130_fd_sc_hd__nand2_1
X_1434_ gamelogic.indexCorrect\[3\] vssd1 vssd1 vccd1 vccd1 _0388_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_169_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3104_ clknet_leaf_28_clk _0094_ vssd1 vssd1 vccd1 vccd1 lcdPlayer.cnt_500hz\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_179_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3035_ clknet_leaf_7_clk clock_div.next_count\[15\] net213 vssd1 vssd1 vccd1 vccd1
+ clock_div.count\[15\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_128_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2652__A2 net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_187_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2481__B net139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2819_ message_reg.state\[0\] net89 _0370_ vssd1 vssd1 vccd1 vccd1 _0216_ sky130_fd_sc_hd__o21a_1
XFILLER_0_33_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input8_X net8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_185_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout63_A _1391_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3522__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_166_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_330 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3008__A net221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_176_Right_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_181_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2634__A2 _1072_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_354 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_31_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1983_ gamelogic.state\[2\] _0813_ vssd1 vssd1 vccd1 vccd1 _0816_ sky130_fd_sc_hd__nand2_1
XFILLER_0_172_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2604_ lcdPlayer.nextState\[3\] _1060_ _1061_ _1063_ _1156_ vssd1 vssd1 vccd1 vccd1
+ _1177_ sky130_fd_sc_hd__a41o_1
XFILLER_0_23_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3584_ net157 vssd1 vssd1 vccd1 vccd1 net14 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_140_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2535_ hostdisp.bottom\[41\] net105 _1106_ hostdisp.top\[57\] _1111_ vssd1 vssd1
+ vccd1 vccd1 _1112_ sky130_fd_sc_hd__a221o_1
XFILLER_0_100_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_143_Right_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2466_ net344 net70 _1055_ _0828_ vssd1 vssd1 vccd1 vccd1 _0162_ sky130_fd_sc_hd__a22o_1
X_1417_ keypadFSMPlayer.state\[2\] vssd1 vssd1 vccd1 vccd1 _0371_ sky130_fd_sc_hd__inv_2
XFILLER_0_48_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2397_ net278 _1020_ _1023_ vssd1 vssd1 vccd1 vccd1 _0125_ sky130_fd_sc_hd__o21a_1
XFILLER_0_97_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3018_ net219 vssd1 vssd1 vccd1 vccd1 _0043_ sky130_fd_sc_hd__inv_2
XANTENNA__1833__B1 _0693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_184 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_137_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_98_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_189_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_110_Right_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout140 gamelogic.letter\[7\] vssd1 vssd1 vccd1 vccd1 net140 sky130_fd_sc_hd__clkbuf_4
Xfanout151 keypadHostt.scan_col\[2\] vssd1 vssd1 vccd1 vccd1 net151 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_148_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout162 net165 vssd1 vssd1 vccd1 vccd1 net162 sky130_fd_sc_hd__clkbuf_4
Xfanout173 net174 vssd1 vssd1 vccd1 vccd1 net173 sky130_fd_sc_hd__clkbuf_2
Xfanout195 net196 vssd1 vssd1 vccd1 vccd1 net195 sky130_fd_sc_hd__clkbuf_4
Xfanout184 net190 vssd1 vssd1 vccd1 vccd1 net184 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_107_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_53_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3418__CLK clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2001__B1 net80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_29_Left_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2320_ lcdPlayer.cnt_500hz\[11\] lcdPlayer.cnt_500hz\[12\] _0971_ lcdPlayer.cnt_500hz\[13\]
+ vssd1 vssd1 vccd1 vccd1 _0976_ sky130_fd_sc_hd__a31o_1
XFILLER_0_85_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2251_ _0938_ net151 _0937_ vssd1 vssd1 vccd1 vccd1 _0048_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_114_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_23_clk_A clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2182_ gamelogic.setWord\[25\] _0893_ net135 vssd1 vssd1 vccd1 vccd1 hostdisp.nextBottom\[73\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_192_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_177_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_125_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2607__A2 _1081_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_38_Left_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1966_ buffer.Rx_byte\[3\] net2 _0803_ vssd1 vssd1 vccd1 vccd1 _0804_ sky130_fd_sc_hd__mux2_1
XFILLER_0_172_176 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1897_ lcdPlayer.cnt_500hz\[0\] lcdPlayer.cnt_500hz\[1\] lcdPlayer.cnt_500hz\[2\]
+ vssd1 vssd1 vccd1 vccd1 _0750_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_47_Left_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3567_ net251 vssd1 vssd1 vccd1 vccd1 gpio_oeb[0] sky130_fd_sc_hd__buf_2
X_2518_ net138 net139 _1094_ vssd1 vssd1 vccd1 vccd1 _1096_ sky130_fd_sc_hd__and3_2
X_3498_ clknet_leaf_4_clk hostdisp.next_curr_word\[20\] net194 vssd1 vssd1 vccd1 vccd1
+ hostdisp.curr_word\[20\] sky130_fd_sc_hd__dfstp_1
X_2449_ hostdisp.curr_word\[22\] net120 vssd1 vssd1 vccd1 vccd1 _1047_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_184_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_56_Left_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_255 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2950__A host_message_reg.Cstate vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2782__A1 host_message_reg.setLetter\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2161__S net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold7 clock_div.count\[29\] vssd1 vssd1 vccd1 vccd1 net271 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_230 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_263 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1820_ clock_div.count\[11\] clock_div.count\[10\] _0703_ vssd1 vssd1 vccd1 vccd1
+ _0707_ sky130_fd_sc_hd__and3_1
XFILLER_0_127_357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1751_ uart_receiver.clk_count\[8\] _0654_ vssd1 vssd1 vccd1 vccd1 _0656_ sky130_fd_sc_hd__and2_1
XFILLER_0_52_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1682_ _0537_ _0564_ _0604_ vssd1 vssd1 vccd1 vccd1 _0605_ sky130_fd_sc_hd__and3_1
XFILLER_0_25_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3390__CLK clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3421_ clknet_leaf_23_clk _0310_ net187 vssd1 vssd1 vccd1 vccd1 dispFSM.guesses\[75\]
+ sky130_fd_sc_hd__dfstp_1
X_3352_ clknet_leaf_20_clk _0241_ net203 vssd1 vssd1 vccd1 vccd1 dispFSM.guesses\[6\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_110_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2303_ lcdPlayer.cnt_500hz\[7\] _0964_ vssd1 vssd1 vccd1 vccd1 _0965_ sky130_fd_sc_hd__and2_1
X_3283_ clknet_leaf_5_clk hostdisp.nextBottom\[81\] net196 vssd1 vssd1 vccd1 vccd1
+ hostdisp.bottom\[81\] sky130_fd_sc_hd__dfrtp_1
X_2234_ _0920_ _0927_ vssd1 vssd1 vccd1 vccd1 gamelogic.nextState\[2\] sky130_fd_sc_hd__or2_1
X_2165_ gamelogic.setWord\[25\] hostdisp.curr_guesses\[25\] net124 vssd1 vssd1 vccd1
+ vccd1 _0885_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2096_ net421 net96 _0851_ net141 vssd1 vssd1 vccd1 vccd1 hostdisp.next_curr_word\[29\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_177_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_177_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_192_238 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout230_A net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2998_ net221 vssd1 vssd1 vccd1 vccd1 _0023_ sky130_fd_sc_hd__inv_2
XFILLER_0_133_316 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1949_ _0184_ _0786_ _0793_ _0779_ vssd1 vssd1 vccd1 vccd1 _0002_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_134_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3619_ net248 vssd1 vssd1 vccd1 vccd1 gpio_out[27] sky130_fd_sc_hd__buf_2
XFILLER_0_141_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_145_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2156__S net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_183_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3016__A net223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_13_Right_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_18_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_211 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3459__Q gamelogic.setWord\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2921_ dispFSM.guesses\[61\] net90 net64 net388 vssd1 vssd1 vccd1 vccd1 _0288_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_61_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2852_ net144 buffer.temp_guess\[1\] _0918_ vssd1 vssd1 vccd1 vccd1 _1383_ sky130_fd_sc_hd__mux2_1
X_1803_ _0696_ _0697_ vssd1 vssd1 vccd1 vccd1 clock_div.next_count\[3\] sky130_fd_sc_hd__nor2_1
X_2783_ host_message_reg.setLetter\[3\] _1290_ _1332_ _1333_ vssd1 vssd1 vccd1 vccd1
+ _0208_ sky130_fd_sc_hd__o22a_1
XFILLER_0_142_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_22_Right_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1734_ uart_receiver.clk_count\[1\] uart_receiver.clk_count\[0\] uart_receiver.clk_count\[2\]
+ vssd1 vssd1 vccd1 vccd1 _0645_ sky130_fd_sc_hd__a21o_1
Xhold204 clock_div.count\[12\] vssd1 vssd1 vccd1 vccd1 net468 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2210__A3 net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold226 hostdisp.top\[75\] vssd1 vssd1 vccd1 vccd1 net490 sky130_fd_sc_hd__dlygate4sd3_1
Xhold215 dispFSM.guesses\[59\] vssd1 vssd1 vccd1 vccd1 net479 sky130_fd_sc_hd__dlygate4sd3_1
Xhold259 uart_transmitter.clk_count\[5\] vssd1 vssd1 vccd1 vccd1 net523 sky130_fd_sc_hd__dlygate4sd3_1
X_1665_ _0591_ keypadFSMPlayer.state\[1\] _0452_ vssd1 vssd1 vccd1 vccd1 _0012_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3404_ clknet_leaf_24_clk _0293_ net189 vssd1 vssd1 vccd1 vccd1 dispFSM.guesses\[58\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_40_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold248 dispFSM.guesses\[8\] vssd1 vssd1 vccd1 vccd1 net512 sky130_fd_sc_hd__dlygate4sd3_1
Xhold237 dispFSM.guesses\[75\] vssd1 vssd1 vccd1 vccd1 net501 sky130_fd_sc_hd__dlygate4sd3_1
X_1596_ net369 net4 _0535_ vssd1 vssd1 vccd1 vccd1 _0055_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3335_ clknet_leaf_0_clk _0224_ net171 vssd1 vssd1 vccd1 vccd1 gamelogic.incorrect\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_3266_ clknet_leaf_5_clk hostdisp.nextBottom\[64\] net199 vssd1 vssd1 vccd1 vccd1
+ hostdisp.bottom\[64\] sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_31_Right_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2217_ buffer.temp_guess\[4\] buffer.temp_guess\[5\] buffer.temp_guess\[6\] buffer.temp_guess\[7\]
+ vssd1 vssd1 vccd1 vccd1 _0913_ sky130_fd_sc_hd__or4_1
XFILLER_0_56_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3286__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3197_ clknet_leaf_23_clk _0173_ vssd1 vssd1 vccd1 vccd1 lcdPlayer.lcd_rs sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout180_A net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_181_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2148_ gamelogic.setWord\[8\] _0876_ net134 vssd1 vssd1 vccd1 vccd1 hostdisp.nextBottom\[56\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_163_84 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2079_ hostdisp.curr_word\[17\] net103 _0845_ gamelogic.letter\[1\] vssd1 vssd1 vccd1
+ vccd1 hostdisp.next_curr_word\[17\] sky130_fd_sc_hd__o22a_1
XFILLER_0_95_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2434__B1 net70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_140_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout233_X net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_40_Right_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_192_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout93_A net94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2122__C1 net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2673__B1 gamelogic.setWord\[37\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_199 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_168_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1450_ hostdisp.curr_word\[0\] vssd1 vssd1 vccd1 vccd1 _0403_ sky130_fd_sc_hd__inv_2
XFILLER_0_120_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3120_ clknet_leaf_18_clk uart_transmitter.next_clk_count\[0\] net223 vssd1 vssd1
+ vccd1 vccd1 uart_transmitter.clk_count\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_93_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3051_ clknet_leaf_10_clk _0046_ net216 vssd1 vssd1 vccd1 vccd1 keypadHostt.scan_col\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_165_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2002_ hostdisp.curr_guesses\[16\] net93 net78 net551 vssd1 vssd1 vccd1 vccd1 hostdisp.next_curr_guesses\[8\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_26_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_147_238 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2416__B1 net69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_0_clk_X clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2904_ dispFSM.guesses\[44\] net83 net60 net498 vssd1 vssd1 vccd1 vccd1 _0271_ sky130_fd_sc_hd__o22a_1
XFILLER_0_42_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3397__SET_B net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2835_ gamelogic.correct\[0\] gamelogic.rights\[0\] _1369_ _1370_ vssd1 vssd1 vccd1
+ vccd1 _1372_ sky130_fd_sc_hd__a22o_1
XFILLER_0_170_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2719__A1 net140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2766_ _1312_ _1316_ _1317_ vssd1 vssd1 vccd1 vccd1 _1319_ sky130_fd_sc_hd__nor3_1
XFILLER_0_13_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1717_ uart_receiver.state\[0\] _0617_ vssd1 vssd1 vccd1 vccd1 _0633_ sky130_fd_sc_hd__nor2_1
X_2697_ _1260_ _1261_ gamelogic.indexCorrect\[3\] vssd1 vssd1 vccd1 vccd1 _1262_ sky130_fd_sc_hd__a21o_1
X_1648_ keypadHostt.scan_col\[0\] _0548_ _0559_ vssd1 vssd1 vccd1 vccd1 _0583_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_6_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1579_ _0514_ _0515_ _0512_ vssd1 vssd1 vccd1 vccd1 _0525_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3318_ clknet_leaf_35_clk uart_receiver.next_clk_count\[10\] net159 vssd1 vssd1 vccd1
+ vccd1 uart_receiver.clk_count\[10\] sky130_fd_sc_hd__dfrtp_1
X_3249_ clknet_leaf_22_clk hostdisp.nextBottom\[47\] net202 vssd1 vssd1 vccd1 vccd1
+ hostdisp.bottom\[47\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_174_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2655__B1 net108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_193_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_193_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_157_Right_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1574__A dispFSM.msg\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout96_X net96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2646__B1 _1096_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_160_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_2_clk_X clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_184_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2620_ hostdisp.bottom\[77\] dispFSM.guesses\[53\] net227 vssd1 vssd1 vccd1 vccd1
+ _1193_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_179_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_124_Right_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2551_ hostdisp.top\[74\] _1095_ _1096_ hostdisp.top\[66\] _1126_ vssd1 vssd1 vccd1
+ vccd1 _1127_ sky130_fd_sc_hd__a221o_1
X_1502_ _0434_ _0443_ vssd1 vssd1 vccd1 vccd1 _0453_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_10_Left_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2482_ lcdPlayer.nextState\[5\] lcdPlayer.nextState\[4\] vssd1 vssd1 vccd1 vccd1
+ _1061_ sky130_fd_sc_hd__and2b_2
XANTENNA__2867__X _1391_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1433_ gamelogic.setWord\[25\] vssd1 vssd1 vccd1 vccd1 _0387_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_169_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3103_ clknet_leaf_28_clk _0093_ vssd1 vssd1 vccd1 vccd1 lcdPlayer.cnt_500hz\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_179_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3034_ clknet_leaf_10_clk clock_div.next_count\[14\] net213 vssd1 vssd1 vccd1 vccd1
+ clock_div.count\[14\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__2637__B1 _1097_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_128_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_40 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout143_A gamelogic.letter\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3474__CLK clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2818_ gamelogic.rights\[2\] _1358_ _1359_ _1361_ vssd1 vssd1 vccd1 vccd1 _0215_
+ sky130_fd_sc_hd__a22o_1
X_2749_ net152 _0363_ _0546_ keypadHostt.scan_col\[3\] vssd1 vssd1 vccd1 vccd1 _1303_
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_143_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2672__B net144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2800__B1 _0394_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2687__X _1252_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2619__A0 hostdisp.bottom\[101\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3347__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_294 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2095__B2 net142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2582__B net139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_184_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_366 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3497__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_157_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1982_ gamelogic.state\[2\] _0813_ vssd1 vssd1 vccd1 vccd1 _0815_ sky130_fd_sc_hd__and2_1
XANTENNA__3467__Q gamelogic.setWord\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2603_ net295 net106 _1176_ net188 vssd1 vssd1 vccd1 vccd1 _0178_ sky130_fd_sc_hd__o211a_1
X_3583_ net157 vssd1 vssd1 vccd1 vccd1 net13 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2534_ hostdisp.bottom\[81\] net118 net109 hostdisp.bottom\[57\] vssd1 vssd1 vccd1
+ vccd1 _1111_ sky130_fd_sc_hd__a22o_1
XFILLER_0_23_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_108 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2465_ hostdisp.curr_word\[30\] net119 vssd1 vssd1 vccd1 vccd1 _1055_ sky130_fd_sc_hd__or2_1
XANTENNA__2570__A2 net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1416_ message_reg.state\[1\] vssd1 vssd1 vccd1 vccd1 _0370_ sky130_fd_sc_hd__inv_2
XANTENNA__2858__A0 net142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2396_ _0017_ _1022_ vssd1 vssd1 vccd1 vccd1 _1023_ sky130_fd_sc_hd__nor2_1
X_3017_ net223 vssd1 vssd1 vccd1 vccd1 _0042_ sky130_fd_sc_hd__inv_2
XFILLER_0_64_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3517__RESET_B net169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_190_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_190_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_189_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout130 _0375_ vssd1 vssd1 vccd1 vccd1 net130 sky130_fd_sc_hd__buf_2
Xfanout152 net153 vssd1 vssd1 vccd1 vccd1 net152 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_148_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout163 net164 vssd1 vssd1 vccd1 vccd1 net163 sky130_fd_sc_hd__clkbuf_4
Xfanout141 gamelogic.letter\[5\] vssd1 vssd1 vccd1 vccd1 net141 sky130_fd_sc_hd__buf_4
Xfanout174 net180 vssd1 vssd1 vccd1 vccd1 net174 sky130_fd_sc_hd__clkbuf_4
Xfanout196 net200 vssd1 vssd1 vccd1 vccd1 net196 sky130_fd_sc_hd__clkbuf_4
Xfanout185 net190 vssd1 vssd1 vccd1 vccd1 net185 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_45_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_69_Right_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_154_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_53_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_181_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3019__A net223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_78_Right_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_176_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2552__A2 net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2250_ _0362_ _0559_ vssd1 vssd1 vccd1 vccd1 _0938_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_114_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2181_ gamelogic.setWord\[33\] hostdisp.curr_guesses\[33\] net124 vssd1 vssd1 vccd1
+ vccd1 _0893_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2068__B2 gamelogic.letter\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_87_Right_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_347 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1965_ uart_receiver.bit_index\[2\] net149 uart_receiver.bit_index\[0\] vssd1 vssd1
+ vccd1 vccd1 _0803_ sky130_fd_sc_hd__and3b_1
XFILLER_0_160_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1896_ net276 net533 vssd1 vssd1 vccd1 vccd1 _0749_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_96_Right_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3566_ clknet_leaf_7_clk hostdisp.next_state net197 vssd1 vssd1 vccd1 vccd1 hostdisp.Cstate
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout106_A _0759_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2543__A2 net114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3497_ clknet_leaf_4_clk hostdisp.next_curr_word\[19\] net179 vssd1 vssd1 vccd1 vccd1
+ hostdisp.curr_word\[19\] sky130_fd_sc_hd__dfstp_1
XANTENNA__3512__CLK clknet_leaf_31_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2517_ _1070_ _1093_ vssd1 vssd1 vccd1 vccd1 _1095_ sky130_fd_sc_hd__nor2_4
X_2448_ net325 net71 _1046_ vssd1 vssd1 vccd1 vccd1 _0153_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_59_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2379_ _1010_ _1011_ vssd1 vssd1 vccd1 vccd1 _0119_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_184_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_3_Left_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2059__B2 net140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_182_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_212 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_267 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_155 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3192__CLK clknet_leaf_31_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2534__A2 net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold8 hostdisp.top\[53\] vssd1 vssd1 vccd1 vccd1 net272 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_159_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3021__RESET_B net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_130 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_166 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_144 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1750_ _0641_ _0653_ _0655_ vssd1 vssd1 vccd1 vccd1 uart_receiver.next_clk_count\[7\]
+ sky130_fd_sc_hd__and3_1
XANTENNA__2222__A1 net100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1476__B net6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3535__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1681_ _0597_ _0603_ vssd1 vssd1 vccd1 vccd1 _0604_ sky130_fd_sc_hd__nor2_1
XFILLER_0_111_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_187_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3420_ clknet_leaf_20_clk _0309_ net203 vssd1 vssd1 vccd1 vccd1 dispFSM.guesses\[74\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_110_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_96_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3351_ clknet_leaf_22_clk net322 net201 vssd1 vssd1 vccd1 vccd1 dispFSM.guesses\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__2525__A2 _1096_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2302_ _0964_ _0956_ _0963_ vssd1 vssd1 vccd1 vccd1 _0089_ sky130_fd_sc_hd__and3b_1
X_3282_ clknet_leaf_6_clk hostdisp.nextBottom\[80\] net191 vssd1 vssd1 vccd1 vccd1
+ hostdisp.bottom\[80\] sky130_fd_sc_hd__dfrtp_1
X_2233_ _0916_ _0926_ vssd1 vssd1 vccd1 vccd1 _0927_ sky130_fd_sc_hd__nand2_1
X_2164_ gamelogic.setWord\[16\] _0884_ net134 vssd1 vssd1 vccd1 vccd1 hostdisp.nextBottom\[64\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_64_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2095_ hostdisp.curr_word\[28\] net101 _0850_ net142 vssd1 vssd1 vccd1 vccd1 hostdisp.next_curr_word\[28\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_61_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_152_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_87 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2997_ net221 vssd1 vssd1 vccd1 vccd1 _0022_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout223_A net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1948_ _0783_ _0786_ _0187_ vssd1 vssd1 vccd1 vccd1 _0793_ sky130_fd_sc_hd__a21oi_1
X_1879_ uart_transmitter.clk_count\[4\] uart_transmitter.clk_count\[3\] _0734_ vssd1
+ vssd1 vccd1 vccd1 _0739_ sky130_fd_sc_hd__and3_1
XFILLER_0_16_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_134_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3618_ lcdPlayer.lcd_rs vssd1 vssd1 vccd1 vccd1 net37 sky130_fd_sc_hd__clkbuf_1
XANTENNA_fanout109_X net109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3549_ clknet_leaf_22_clk hostdisp.next_curr_guesses\[31\] net201 vssd1 vssd1 vccd1
+ vccd1 hostdisp.curr_guesses\[31\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_145_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2452__B2 net73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2452__A1 net130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3558__CLK clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_22_clk_A clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2172__S net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_151_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_151_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2204__A1 net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_151_136 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_2_3__f_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_2_3__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_159_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkload1_A clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_122_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2920_ dispFSM.guesses\[60\] net83 net58 net499 vssd1 vssd1 vccd1 vccd1 _0287_ sky130_fd_sc_hd__o22a_1
XANTENNA__2443__A1 net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2851_ net66 _1382_ vssd1 vssd1 vccd1 vccd1 _0227_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_75_Left_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_170_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1802_ net375 _0694_ vssd1 vssd1 vccd1 vccd1 _0697_ sky130_fd_sc_hd__nor2_1
X_2782_ host_message_reg.setLetter\[3\] _0601_ _1310_ _0597_ vssd1 vssd1 vccd1 vccd1
+ _1333_ sky130_fd_sc_hd__a211o_1
XFILLER_0_110_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3475__Q gamelogic.setWord\[37\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1733_ uart_receiver.clk_count\[1\] uart_receiver.clk_count\[0\] uart_receiver.clk_count\[2\]
+ vssd1 vssd1 vccd1 vccd1 _0644_ sky130_fd_sc_hd__nand3_1
Xhold216 dispFSM.guesses\[66\] vssd1 vssd1 vccd1 vccd1 net480 sky130_fd_sc_hd__dlygate4sd3_1
Xhold205 dispFSM.guesses\[10\] vssd1 vssd1 vccd1 vccd1 net469 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1664_ keypadFSMPlayer.state\[5\] _0489_ _0491_ vssd1 vssd1 vccd1 vccd1 _0591_ sky130_fd_sc_hd__and3_1
X_3403_ clknet_leaf_20_clk _0292_ net205 vssd1 vssd1 vccd1 vccd1 dispFSM.guesses\[57\]
+ sky130_fd_sc_hd__dfstp_1
Xhold238 dispFSM.guesses\[58\] vssd1 vssd1 vccd1 vccd1 net502 sky130_fd_sc_hd__dlygate4sd3_1
Xhold249 dispFSM.guesses\[56\] vssd1 vssd1 vccd1 vccd1 net513 sky130_fd_sc_hd__dlygate4sd3_1
Xhold227 hostdisp.curr_guesses\[18\] vssd1 vssd1 vccd1 vccd1 net491 sky130_fd_sc_hd__dlygate4sd3_1
X_1595_ net497 net232 _0535_ vssd1 vssd1 vccd1 vccd1 _0056_ sky130_fd_sc_hd__mux2_1
XFILLER_0_40_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3334_ clknet_leaf_0_clk _0223_ net171 vssd1 vssd1 vccd1 vccd1 gamelogic.correct\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_3265_ clknet_leaf_22_clk hostdisp.nextBottom\[63\] net186 vssd1 vssd1 vccd1 vccd1
+ hostdisp.bottom\[63\] sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_84_Left_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2216_ gamelogic.state\[0\] gamelogic.state\[1\] _0365_ gamelogic.state\[2\] vssd1
+ vssd1 vccd1 vccd1 _0912_ sky130_fd_sc_hd__or4_2
X_3196_ clknet_leaf_30_clk _0172_ net185 vssd1 vssd1 vccd1 vccd1 hostdisp.top\[101\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_1_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_181_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2147_ gamelogic.setWord\[16\] hostdisp.curr_guesses\[16\] net124 vssd1 vssd1 vccd1
+ vccd1 _0876_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2078_ hostdisp.curr_word\[16\] net103 _0845_ net145 vssd1 vssd1 vccd1 vccd1 hostdisp.next_curr_word\[16\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_72_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_163_96 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_138_Right_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_140_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2985__A2 net53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_93_Left_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_192_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout226_X net226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3380__CLK clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_105_Right_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_15_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2189__A0 gamelogic.setWord\[37\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_331 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_184_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3050_ clknet_leaf_15_clk _0045_ net221 vssd1 vssd1 vccd1 vccd1 keypadFSMPlayer.strobe
+ sky130_fd_sc_hd__dfrtp_1
X_2001_ hostdisp.curr_guesses\[15\] _0823_ net80 net345 vssd1 vssd1 vccd1 vccd1 hostdisp.next_curr_guesses\[7\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_26_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2967__A2 net53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2903_ dispFSM.guesses\[43\] net81 net57 net557 vssd1 vssd1 vccd1 vccd1 _0270_ sky130_fd_sc_hd__o22a_1
XFILLER_0_155_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2834_ gamelogic.correct\[0\] gamelogic.rights\[0\] _1369_ _1370_ vssd1 vssd1 vccd1
+ vccd1 _1371_ sky130_fd_sc_hd__nand4_1
X_2765_ _1316_ _1317_ vssd1 vssd1 vccd1 vccd1 _1318_ sky130_fd_sc_hd__nor2_1
XFILLER_0_115_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1716_ uart_receiver.state\[2\] _0396_ _0621_ net127 _0617_ vssd1 vssd1 vccd1 vccd1
+ _0632_ sky130_fd_sc_hd__o221a_1
X_2696_ gamelogic.state\[0\] _0922_ _1235_ vssd1 vssd1 vccd1 vccd1 _1261_ sky130_fd_sc_hd__o21ai_1
X_1647_ _0579_ _0580_ _0581_ vssd1 vssd1 vccd1 vccd1 _0582_ sky130_fd_sc_hd__nor3_1
XANTENNA__3253__CLK clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1578_ dispFSM.msg\[2\] _0447_ vssd1 vssd1 vccd1 vccd1 _0524_ sky130_fd_sc_hd__and2_1
XFILLER_0_6_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3317_ clknet_leaf_34_clk uart_receiver.next_clk_count\[9\] net159 vssd1 vssd1 vccd1
+ vccd1 uart_receiver.clk_count\[9\] sky130_fd_sc_hd__dfrtp_1
X_3248_ clknet_leaf_5_clk hostdisp.nextBottom\[46\] net193 vssd1 vssd1 vccd1 vccd1
+ hostdisp.bottom\[46\] sky130_fd_sc_hd__dfrtp_1
X_3179_ clknet_leaf_22_clk _0155_ net185 vssd1 vssd1 vccd1 vccd1 hostdisp.top\[63\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout176_X net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_101_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_20_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1590__A dispFSM.msg\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2686__A net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_160_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_184_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_149_Left_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3276__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2550_ hostdisp.bottom\[82\] net118 net112 hostdisp.bottom\[74\] vssd1 vssd1 vccd1
+ vccd1 _1126_ sky130_fd_sc_hd__a22o_1
X_1501_ _0434_ _0444_ vssd1 vssd1 vccd1 vccd1 _0452_ sky130_fd_sc_hd__or2_1
X_2481_ net138 net139 vssd1 vssd1 vccd1 vccd1 _1060_ sky130_fd_sc_hd__or2_4
X_1432_ net140 vssd1 vssd1 vccd1 vccd1 _0386_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_158_Left_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3102_ clknet_leaf_28_clk _0092_ vssd1 vssd1 vccd1 vccd1 lcdPlayer.cnt_500hz\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_3033_ clknet_leaf_10_clk clock_div.next_count\[13\] net213 vssd1 vssd1 vccd1 vccd1
+ clock_div.count\[13\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_128_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_187_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_34_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_167_Left_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout136_A net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3571__255 vssd1 vssd1 vccd1 vccd1 net255 _3571__255/LO sky130_fd_sc_hd__conb_1
XFILLER_0_103_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2817_ gamelogic.rights\[2\] _1360_ vssd1 vssd1 vccd1 vccd1 _1361_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_82_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2748_ net151 _0560_ vssd1 vssd1 vccd1 vccd1 _1302_ sky130_fd_sc_hd__nor2_1
XFILLER_0_169_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2573__B1 net109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2679_ gamelogic.setWord\[38\] _0385_ gamelogic.setWord\[39\] _0386_ vssd1 vssd1
+ vccd1 vccd1 _1245_ sky130_fd_sc_hd__a22oi_1
XPHY_EDGE_ROW_176_Left_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3413__SET_B net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_190_Right_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout49_A net50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2800__B2 gamelogic.letter\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1585__A dispFSM.msg\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_176_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_56_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_184_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_378 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1981_ gamelogic.state\[0\] gamelogic.state\[3\] gamelogic.state\[1\] vssd1 vssd1
+ vccd1 vccd1 _0814_ sky130_fd_sc_hd__or3b_1
XFILLER_0_184_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2602_ _0360_ _1166_ _1172_ _1175_ _1159_ vssd1 vssd1 vccd1 vccd1 _1176_ sky130_fd_sc_hd__a2111o_1
X_3582_ net258 vssd1 vssd1 vccd1 vccd1 gpio_oeb[15] sky130_fd_sc_hd__buf_2
X_2533_ hostdisp.bottom\[73\] net112 _1096_ hostdisp.top\[65\] vssd1 vssd1 vccd1 vccd1
+ _1110_ sky130_fd_sc_hd__a22o_1
XFILLER_0_23_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2555__B1 _0360_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_139_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_7 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2464_ _1029_ _1054_ net67 net350 vssd1 vssd1 vccd1 vccd1 _0161_ sky130_fd_sc_hd__o2bb2a_1
X_1415_ keypadFSMHost.state\[5\] vssd1 vssd1 vccd1 vccd1 _0369_ sky130_fd_sc_hd__inv_2
XFILLER_0_48_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2395_ lcdPlayer.cnt_20ms\[18\] lcdPlayer.cnt_20ms\[17\] lcdPlayer.cnt_20ms\[16\]
+ _1017_ vssd1 vssd1 vccd1 vccd1 _1022_ sky130_fd_sc_hd__and4_1
X_3016_ net223 vssd1 vssd1 vccd1 vccd1 _0041_ sky130_fd_sc_hd__inv_2
XANTENNA__1818__C1 _0693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3441__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout139_X net139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_31_clk clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_31_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_190_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_137_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_2_1__f_clk_X clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout120 _0859_ vssd1 vssd1 vccd1 vccd1 net120 sky130_fd_sc_hd__buf_2
Xfanout131 net132 vssd1 vssd1 vccd1 vccd1 net131 sky130_fd_sc_hd__clkbuf_4
Xfanout153 keypadHostt.scan_col\[1\] vssd1 vssd1 vccd1 vccd1 net153 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_148_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout164 net165 vssd1 vssd1 vccd1 vccd1 net164 sky130_fd_sc_hd__clkbuf_4
Xfanout142 gamelogic.letter\[4\] vssd1 vssd1 vccd1 vccd1 net142 sky130_fd_sc_hd__buf_4
Xfanout197 net199 vssd1 vssd1 vccd1 vccd1 net197 sky130_fd_sc_hd__clkbuf_4
Xfanout186 net190 vssd1 vssd1 vccd1 vccd1 net186 sky130_fd_sc_hd__clkbuf_2
Xfanout175 net176 vssd1 vssd1 vccd1 vccd1 net175 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_69_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2175__S net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_175 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_22_clk clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_22_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_181_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2537__B1 _1098_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2001__A2 _0823_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3314__CLK clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2180_ gamelogic.setWord\[24\] _0892_ net134 vssd1 vssd1 vccd1 vccd1 hostdisp.nextBottom\[72\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_192_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3464__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2473__C1 _1034_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_177_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_13_clk clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_13_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_7_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1964_ net2 _0801_ _0802_ _0618_ vssd1 vssd1 vccd1 vccd1 uart_receiver.temp_byte\[2\]
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_172_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_160_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1895_ _0400_ _0748_ net116 vssd1 vssd1 vccd1 vccd1 uart_transmitter.next_clk_count\[10\]
+ sky130_fd_sc_hd__a21boi_1
XANTENNA__2114__A _0827_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3565_ clknet_leaf_22_clk hostdisp.next_curr_guesses\[47\] net201 vssd1 vssd1 vccd1
+ vccd1 hostdisp.curr_guesses\[47\] sky130_fd_sc_hd__dfrtp_1
X_3496_ clknet_leaf_4_clk hostdisp.next_curr_word\[18\] net194 vssd1 vssd1 vccd1 vccd1
+ hostdisp.curr_word\[18\] sky130_fd_sc_hd__dfstp_1
X_2516_ _1093_ vssd1 vssd1 vccd1 vccd1 _1094_ sky130_fd_sc_hd__inv_2
X_2447_ net136 host_message_reg.setLetter\[5\] hostdisp.curr_word\[21\] _1031_ net67
+ vssd1 vssd1 vccd1 vccd1 _1046_ sky130_fd_sc_hd__o221a_1
XFILLER_0_166_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_59_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2378_ net399 _1008_ net168 vssd1 vssd1 vccd1 vccd1 _1011_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_184_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2059__A2 net96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_143_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3391__RESET_B net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2950__C keypadFSMHost.state\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_104_Left_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3487__CLK clknet_leaf_30_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout71_X net71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold9 lcdPlayer.cnt_20ms\[20\] vssd1 vssd1 vccd1 vccd1 net273 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_57_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2470__A2 net75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_154_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_142_318 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1680_ _0598_ _0602_ vssd1 vssd1 vccd1 vccd1 _0603_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_116_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3350_ clknet_leaf_24_clk _0239_ net188 vssd1 vssd1 vccd1 vccd1 dispFSM.guesses\[4\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_96_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2301_ lcdPlayer.cnt_500hz\[5\] lcdPlayer.cnt_500hz\[4\] lcdPlayer.cnt_500hz\[6\]
+ _0751_ vssd1 vssd1 vccd1 vccd1 _0964_ sky130_fd_sc_hd__and4_1
X_3281_ clknet_leaf_22_clk hostdisp.nextBottom\[79\] net186 vssd1 vssd1 vccd1 vccd1
+ hostdisp.bottom\[79\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_188_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2232_ _0908_ _0922_ vssd1 vssd1 vccd1 vccd1 _0926_ sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_2_clk clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_2_clk
+ sky130_fd_sc_hd__clkbuf_8
X_2163_ gamelogic.setWord\[24\] hostdisp.curr_guesses\[24\] net125 vssd1 vssd1 vccd1
+ vccd1 _0884_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_119_Right_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_88_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2094_ hostdisp.curr_word\[27\] net101 _0850_ net143 vssd1 vssd1 vccd1 vccd1 hostdisp.next_curr_word\[27\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_177_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_64_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_99 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_74 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2996_ net222 vssd1 vssd1 vccd1 vccd1 _0021_ sky130_fd_sc_hd__inv_2
XFILLER_0_145_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1947_ _0779_ _0787_ _0792_ _0773_ vssd1 vssd1 vccd1 vccd1 _0001_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout216_A net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1878_ uart_transmitter.clk_count\[4\] _0736_ vssd1 vssd1 vccd1 vccd1 _0738_ sky130_fd_sc_hd__or2_1
XFILLER_0_31_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1972__A1 net2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3617_ uart_transmitter.tx_serial vssd1 vssd1 vccd1 vccd1 net36 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3548_ clknet_leaf_6_clk hostdisp.next_curr_guesses\[30\] net191 vssd1 vssd1 vccd1
+ vccd1 hostdisp.curr_guesses\[30\] sky130_fd_sc_hd__dfstp_1
XFILLER_0_3_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_177_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3479_ clknet_leaf_32_clk hostdisp.next_curr_word\[1\] net163 vssd1 vssd1 vccd1 vccd1
+ hostdisp.curr_word\[1\] sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_4_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2452__A2 host_message_reg.setLetter\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_112_Left_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2689__A net142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_121_Left_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_163_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2691__A2 gamelogic.setWord\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_122_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2443__A2 host_message_reg.setLetter\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3502__CLK clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_123 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2850_ net145 buffer.temp_guess\[0\] _0918_ vssd1 vssd1 vccd1 vccd1 _1382_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1801_ clock_div.count\[1\] clock_div.count\[0\] clock_div.count\[3\] clock_div.count\[2\]
+ vssd1 vssd1 vccd1 vccd1 _0696_ sky130_fd_sc_hd__and4_1
XFILLER_0_72_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2781_ _1327_ _1331_ vssd1 vssd1 vccd1 vccd1 _1332_ sky130_fd_sc_hd__xor2_1
XPHY_EDGE_ROW_130_Left_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1732_ _0635_ _0641_ _0643_ vssd1 vssd1 vccd1 vccd1 uart_receiver.next_clk_count\[1\]
+ sky130_fd_sc_hd__and3_1
X_1663_ _0016_ _0014_ _0590_ vssd1 vssd1 vccd1 vccd1 keypadFSMPlayer.next_state\[0\]
+ sky130_fd_sc_hd__or3_1
Xhold217 dispFSM.guesses\[17\] vssd1 vssd1 vccd1 vccd1 net481 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold206 hostdisp.top\[74\] vssd1 vssd1 vccd1 vccd1 net470 sky130_fd_sc_hd__dlygate4sd3_1
Xhold239 clock_div.count\[25\] vssd1 vssd1 vccd1 vccd1 net503 sky130_fd_sc_hd__dlygate4sd3_1
Xhold228 hostdisp.curr_guesses\[40\] vssd1 vssd1 vccd1 vccd1 net492 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3402_ clknet_leaf_23_clk _0291_ net184 vssd1 vssd1 vccd1 vccd1 dispFSM.guesses\[56\]
+ sky130_fd_sc_hd__dfstp_1
X_1594_ net378 net6 _0535_ vssd1 vssd1 vccd1 vccd1 _0057_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3333_ clknet_leaf_0_clk _0222_ net171 vssd1 vssd1 vccd1 vccd1 gamelogic.correct\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_3264_ clknet_leaf_5_clk hostdisp.nextBottom\[62\] net193 vssd1 vssd1 vccd1 vccd1
+ hostdisp.bottom\[62\] sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_7_Right_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2215_ gamelogic.state\[0\] gamelogic.state\[1\] _0365_ gamelogic.state\[2\] vssd1
+ vssd1 vccd1 vccd1 _0911_ sky130_fd_sc_hd__nor4_1
XTAP_TAPCELL_ROW_1_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3195_ clknet_leaf_29_clk _0171_ net166 vssd1 vssd1 vccd1 vccd1 hostdisp.top\[79\]
+ sky130_fd_sc_hd__dfrtp_1
X_2146_ gamelogic.setWord\[7\] _0875_ net136 vssd1 vssd1 vccd1 vccd1 hostdisp.nextBottom\[55\]
+ sky130_fd_sc_hd__mux2_1
XANTENNA__2682__A2 _1247_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2077_ _0845_ vssd1 vssd1 vccd1 vccd1 _0846_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout166_A net169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3182__CLK clknet_leaf_31_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2434__A2 net73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_140_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2979_ gamelogic.setWord\[18\] net51 net47 gamelogic.setWord\[26\] vssd1 vssd1 vccd1
+ vccd1 _0342_ sky130_fd_sc_hd__o22a_1
XFILLER_0_16_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_192_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1684__Y _0607_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout79_A _0826_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3581__257 vssd1 vssd1 vccd1 vccd1 net257 _3581__257/LO sky130_fd_sc_hd__conb_1
XANTENNA__3525__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2673__A2 gamelogic.letter\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2425__A2 net70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2000_ hostdisp.curr_guesses\[14\] net94 net78 net390 vssd1 vssd1 vccd1 vccd1 hostdisp.next_curr_guesses\[6\]
+ sky130_fd_sc_hd__o22a_1
XANTENNA__3423__RESET_B net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2902_ dispFSM.guesses\[42\] net84 net59 net466 vssd1 vssd1 vccd1 vccd1 _0269_ sky130_fd_sc_hd__o22a_1
XFILLER_0_42_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2833_ gamelogic.correct\[1\] gamelogic.rights\[1\] vssd1 vssd1 vccd1 vccd1 _1370_
+ sky130_fd_sc_hd__nand2_1
X_2764_ _1298_ _1314_ _1315_ vssd1 vssd1 vccd1 vccd1 _1317_ sky130_fd_sc_hd__nor3_1
XFILLER_0_115_115 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1715_ net127 vssd1 vssd1 vccd1 vccd1 _0631_ sky130_fd_sc_hd__inv_2
XFILLER_0_111_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2695_ _1252_ _1259_ gamelogic.state\[2\] _0814_ vssd1 vssd1 vccd1 vccd1 _1260_ sky130_fd_sc_hd__a211o_1
X_1646_ _0569_ _0570_ _0578_ vssd1 vssd1 vccd1 vccd1 _0581_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_158_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1577_ _0519_ _0521_ _0523_ _0454_ dispFSM.msg\[3\] vssd1 vssd1 vccd1 vccd1 _0061_
+ sky130_fd_sc_hd__o32a_1
XANTENNA_clkload20_A clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_171_Right_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_158_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3316_ clknet_leaf_35_clk uart_receiver.next_clk_count\[8\] net159 vssd1 vssd1 vccd1
+ vccd1 uart_receiver.clk_count\[8\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3548__CLK clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3247_ clknet_leaf_14_clk hostdisp.nextBottom\[45\] net207 vssd1 vssd1 vccd1 vccd1
+ hostdisp.bottom\[45\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_21_clk_A clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2104__B2 net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2655__A2 net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3178_ clknet_leaf_22_clk _0154_ net201 vssd1 vssd1 vccd1 vccd1 hostdisp.top\[62\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_178_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2129_ _0391_ net120 vssd1 vssd1 vccd1 vccd1 _0867_ sky130_fd_sc_hd__nand2_1
XFILLER_0_178_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout169_X net169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_161_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2040__B1 net79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3078__CLK clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2178__S net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2646__A2 net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_160_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2207__A net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_344 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1500_ net380 _0443_ _0451_ vssd1 vssd1 vccd1 vccd1 _0189_ sky130_fd_sc_hd__a21o_1
XFILLER_0_105_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2480_ net138 lcdPlayer.nextState\[0\] vssd1 vssd1 vccd1 vccd1 _1059_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_130_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1431_ gamelogic.letter\[6\] vssd1 vssd1 vccd1 vccd1 _0385_ sky130_fd_sc_hd__inv_2
XFILLER_0_120_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3101_ clknet_leaf_29_clk _0091_ vssd1 vssd1 vccd1 vccd1 lcdPlayer.cnt_500hz\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_170_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3032_ clknet_leaf_9_clk clock_div.next_count\[12\] net214 vssd1 vssd1 vccd1 vccd1
+ clock_div.count\[12\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__2637__A2 _1095_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_175_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2117__A gamelogic.setWord\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_311 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2816_ _0819_ _1359_ _1360_ _1358_ gamelogic.rights\[1\] vssd1 vssd1 vccd1 vccd1
+ _0214_ sky130_fd_sc_hd__a32o_1
XANTENNA__3220__CLK clknet_leaf_31_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2747_ _0612_ _1293_ _1300_ vssd1 vssd1 vccd1 vccd1 _1301_ sky130_fd_sc_hd__or3b_1
XANTENNA__2022__B1 net77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2678_ gamelogic.setWord\[34\] _0379_ gamelogic.setWord\[38\] _0385_ vssd1 vssd1
+ vccd1 vccd1 _1244_ sky130_fd_sc_hd__o22a_1
XFILLER_0_75_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1629_ net153 _0548_ _0556_ _0563_ vssd1 vssd1 vccd1 vccd1 _0564_ sky130_fd_sc_hd__o31a_1
XFILLER_0_78_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3345__RESET_B net164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input3_A gpio_in[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_185_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_178_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_193_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_181_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_182 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_48_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_56_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3243__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1980_ _0364_ gamelogic.state\[1\] _0365_ vssd1 vssd1 vccd1 vccd1 _0813_ sky130_fd_sc_hd__and3_1
XFILLER_0_184_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2601_ net111 _1173_ _1174_ net105 vssd1 vssd1 vccd1 vccd1 _1175_ sky130_fd_sc_hd__a22o_1
X_3581_ net257 vssd1 vssd1 vccd1 vccd1 gpio_oeb[14] sky130_fd_sc_hd__buf_2
XANTENNA__2004__B1 net77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2532_ net292 net106 _1109_ net182 vssd1 vssd1 vccd1 vccd1 _0174_ sky130_fd_sc_hd__o211a_1
XFILLER_0_140_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3482__SET_B net164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_42 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2463_ _0410_ _0827_ vssd1 vssd1 vccd1 vccd1 _1054_ sky130_fd_sc_hd__or2_1
X_1414_ keypadFSMHost.prev_key\[5\] vssd1 vssd1 vccd1 vccd1 _0368_ sky130_fd_sc_hd__inv_2
XFILLER_0_48_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2394_ _1020_ _1021_ vssd1 vssd1 vccd1 vccd1 _0124_ sky130_fd_sc_hd__nor2_1
XFILLER_0_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3015_ net220 vssd1 vssd1 vccd1 vccd1 _0040_ sky130_fd_sc_hd__inv_2
XFILLER_0_155_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_171_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_148_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_171_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout110 _1087_ vssd1 vssd1 vccd1 vccd1 net110 sky130_fd_sc_hd__buf_2
Xfanout121 net122 vssd1 vssd1 vccd1 vccd1 net121 sky130_fd_sc_hd__clkbuf_4
XANTENNA_input6_X net6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout154 net155 vssd1 vssd1 vccd1 vccd1 net154 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_148_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout132 net133 vssd1 vssd1 vccd1 vccd1 net132 sky130_fd_sc_hd__clkbuf_4
Xfanout165 net225 vssd1 vssd1 vccd1 vccd1 net165 sky130_fd_sc_hd__clkbuf_4
Xfanout143 gamelogic.letter\[3\] vssd1 vssd1 vccd1 vccd1 net143 sky130_fd_sc_hd__buf_4
Xfanout198 net199 vssd1 vssd1 vccd1 vccd1 net198 sky130_fd_sc_hd__clkbuf_2
Xfanout176 net179 vssd1 vssd1 vccd1 vccd1 net176 sky130_fd_sc_hd__clkbuf_4
Xfanout187 net189 vssd1 vssd1 vccd1 vccd1 net187 sky130_fd_sc_hd__clkbuf_4
XANTENNA__3266__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_302 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_139_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3619__248 vssd1 vssd1 vccd1 vccd1 _3619__248/HI net248 sky130_fd_sc_hd__conb_1
XFILLER_0_49_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2191__S net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_125_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1963_ buffer.Rx_byte\[2\] _0801_ vssd1 vssd1 vccd1 vccd1 _0802_ sky130_fd_sc_hd__nand2b_1
X_1894_ net116 _0747_ _0748_ vssd1 vssd1 vccd1 vccd1 uart_transmitter.next_clk_count\[9\]
+ sky130_fd_sc_hd__and3_1
XFILLER_0_7_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_180_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_153_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3564_ clknet_leaf_6_clk hostdisp.next_curr_guesses\[46\] net192 vssd1 vssd1 vccd1
+ vccd1 hostdisp.curr_guesses\[46\] sky130_fd_sc_hd__dfstp_1
XFILLER_0_51_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3495_ clknet_leaf_14_clk hostdisp.next_curr_word\[17\] net194 vssd1 vssd1 vccd1
+ vccd1 hostdisp.curr_word\[17\] sky130_fd_sc_hd__dfstp_1
X_2515_ lcdPlayer.nextState\[2\] _1058_ lcdPlayer.nextState\[3\] vssd1 vssd1 vccd1
+ vccd1 _1093_ sky130_fd_sc_hd__or3b_4
X_2446_ net356 _1045_ net67 vssd1 vssd1 vccd1 vccd1 _0152_ sky130_fd_sc_hd__mux2_1
XANTENNA__3289__CLK clknet_leaf_30_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout196_A net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_16_Left_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2377_ lcdPlayer.cnt_20ms\[12\] lcdPlayer.cnt_20ms\[11\] lcdPlayer.cnt_20ms\[10\]
+ _1004_ vssd1 vssd1 vccd1 vccd1 _1010_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_184_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2464__B1 net67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_182_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_143_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_255 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_113_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2758__B2 host_message_reg.setLetter\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_291 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3280_ clknet_leaf_6_clk hostdisp.nextBottom\[78\] net191 vssd1 vssd1 vccd1 vccd1
+ hostdisp.bottom\[78\] sky130_fd_sc_hd__dfrtp_1
X_2300_ lcdPlayer.cnt_500hz\[5\] lcdPlayer.cnt_500hz\[4\] _0751_ lcdPlayer.cnt_500hz\[6\]
+ vssd1 vssd1 vccd1 vccd1 _0963_ sky130_fd_sc_hd__a31o_1
XANTENNA__3431__CLK clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2231_ _0920_ _0921_ _0925_ vssd1 vssd1 vccd1 vccd1 gamelogic.nextState\[1\] sky130_fd_sc_hd__or3_1
X_2162_ gamelogic.setWord\[15\] _0883_ net136 vssd1 vssd1 vccd1 vccd1 hostdisp.nextBottom\[63\]
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_88_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2093_ hostdisp.curr_word\[26\] net101 _0850_ gamelogic.letter\[2\] vssd1 vssd1 vccd1
+ vccd1 hostdisp.next_curr_word\[26\] sky130_fd_sc_hd__o22a_1
XFILLER_0_177_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_64_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_86 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2995_ net222 vssd1 vssd1 vccd1 vccd1 _0020_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_122 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1946_ _0788_ _0791_ vssd1 vssd1 vccd1 vccd1 _0792_ sky130_fd_sc_hd__xnor2_1
X_1877_ _0736_ _0737_ net116 vssd1 vssd1 vccd1 vccd1 uart_transmitter.next_clk_count\[3\]
+ sky130_fd_sc_hd__and3b_1
XFILLER_0_31_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3616_ net247 vssd1 vssd1 vccd1 vccd1 gpio_out[24] sky130_fd_sc_hd__buf_2
XANTENNA_fanout111_A _1085_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3547_ clknet_leaf_14_clk net392 net208 vssd1 vssd1 vccd1 vccd1 hostdisp.curr_guesses\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_101_92 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3478_ clknet_leaf_31_clk hostdisp.next_curr_word\[0\] net163 vssd1 vssd1 vccd1 vccd1
+ hostdisp.curr_word\[0\] sky130_fd_sc_hd__dfstp_1
XFILLER_0_86_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2795__A host_message_reg.setLetter\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2429_ net334 net68 _1037_ _1029_ vssd1 vssd1 vccd1 vccd1 _0143_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_145_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3541__RESET_B net206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3304__CLK clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_185_Right_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3454__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2676__B1 gamelogic.indexCorrect\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_163_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_159_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_18_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1800_ _0694_ _0695_ vssd1 vssd1 vccd1 vccd1 clock_div.next_count\[2\] sky130_fd_sc_hd__nor2_1
XFILLER_0_127_135 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2780_ net232 _0560_ _1323_ vssd1 vssd1 vccd1 vccd1 _1331_ sky130_fd_sc_hd__and3_1
XFILLER_0_25_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1731_ uart_receiver.clk_count\[1\] uart_receiver.clk_count\[0\] vssd1 vssd1 vccd1
+ vccd1 _0643_ sky130_fd_sc_hd__nand2_1
X_1662_ _0443_ _0445_ _0589_ _0453_ keypadFSMPlayer.state\[4\] vssd1 vssd1 vccd1 vccd1
+ _0590_ sky130_fd_sc_hd__a32o_1
XPHY_EDGE_ROW_152_Right_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold207 dispFSM.guesses\[12\] vssd1 vssd1 vccd1 vccd1 net471 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_133_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold218 dispFSM.guesses\[79\] vssd1 vssd1 vccd1 vccd1 net482 sky130_fd_sc_hd__dlygate4sd3_1
X_3401_ clknet_leaf_15_clk net445 net207 vssd1 vssd1 vccd1 vccd1 dispFSM.guesses\[55\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold229 lcdPlayer.cnt_500hz\[9\] vssd1 vssd1 vccd1 vccd1 net493 sky130_fd_sc_hd__dlygate4sd3_1
X_1593_ _0535_ vssd1 vssd1 vccd1 vccd1 _0536_ sky130_fd_sc_hd__inv_2
XFILLER_0_21_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3332_ clknet_leaf_35_clk _0221_ net165 vssd1 vssd1 vccd1 vccd1 gamelogic.correct\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_0_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3263_ clknet_leaf_15_clk hostdisp.nextBottom\[61\] net209 vssd1 vssd1 vccd1 vccd1
+ hostdisp.bottom\[61\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_147_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2214_ net100 _0909_ vssd1 vssd1 vccd1 vccd1 _0910_ sky130_fd_sc_hd__nor2_1
X_3194_ clknet_leaf_31_clk _0170_ net173 vssd1 vssd1 vccd1 vccd1 hostdisp.top\[78\]
+ sky130_fd_sc_hd__dfrtp_1
X_2145_ gamelogic.setWord\[15\] hostdisp.curr_guesses\[15\] net126 vssd1 vssd1 vccd1
+ vccd1 _0875_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_1_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2076_ _0842_ _0844_ vssd1 vssd1 vccd1 vccd1 _0845_ sky130_fd_sc_hd__nand2_2
XFILLER_0_95_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3327__CLK clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2419__B1 net67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_140_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3477__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2978_ gamelogic.setWord\[17\] net54 net50 gamelogic.setWord\[25\] vssd1 vssd1 vccd1
+ vccd1 _0341_ sky130_fd_sc_hd__o22a_1
XFILLER_0_16_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_192_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_138 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1929_ _0185_ _0776_ vssd1 vssd1 vccd1 vccd1 _0777_ sky130_fd_sc_hd__nor2_1
XFILLER_0_114_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout114_X net114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_151_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_110_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2122__A2 net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_23_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2649__B1 net109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold90 hostdisp.top\[66\] vssd1 vssd1 vccd1 vccd1 net354 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2901_ dispFSM.guesses\[41\] net86 net62 net541 vssd1 vssd1 vccd1 vccd1 _0268_ sky130_fd_sc_hd__o22a_1
XFILLER_0_42_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2832_ gamelogic.correct\[1\] gamelogic.rights\[1\] vssd1 vssd1 vccd1 vccd1 _1369_
+ sky130_fd_sc_hd__or2_1
X_2763_ _1298_ _1315_ _1314_ vssd1 vssd1 vccd1 vccd1 _1316_ sky130_fd_sc_hd__o21a_1
XFILLER_0_155_285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1714_ uart_receiver.state\[0\] uart_receiver.state\[1\] uart_receiver.state\[2\]
+ vssd1 vssd1 vccd1 vccd1 _0630_ sky130_fd_sc_hd__or3b_2
XFILLER_0_53_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2694_ _0377_ gamelogic.setWord\[24\] _1253_ _1256_ _1258_ vssd1 vssd1 vccd1 vccd1
+ _1259_ sky130_fd_sc_hd__o2111a_1
X_1645_ _0572_ _0577_ _0566_ _0568_ vssd1 vssd1 vccd1 vccd1 _0580_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_111_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1576_ _0437_ _0522_ _0448_ vssd1 vssd1 vccd1 vccd1 _0523_ sky130_fd_sc_hd__o21a_1
XFILLER_0_158_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkload13_A clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3315_ clknet_leaf_35_clk uart_receiver.next_clk_count\[7\] net161 vssd1 vssd1 vccd1
+ vccd1 uart_receiver.clk_count\[7\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_74 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3246_ clknet_leaf_22_clk hostdisp.nextBottom\[44\] net186 vssd1 vssd1 vccd1 vccd1
+ hostdisp.bottom\[44\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_174_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3177_ clknet_leaf_14_clk _0153_ net202 vssd1 vssd1 vccd1 vccd1 hostdisp.top\[61\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2128_ hostdisp.curr_guesses\[6\] net120 _0866_ net134 vssd1 vssd1 vccd1 vccd1 hostdisp.nextBottom\[46\]
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_95_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_37_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2059_ net514 net96 _0836_ net140 vssd1 vssd1 vccd1 vccd1 hostdisp.next_curr_word\[7\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_190_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_190_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout231_X net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_211 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_90 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2040__A1 gamelogic.letter\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2591__A2 _1097_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_8_Left_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout91_A net92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_160_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2194__S net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_140_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1430_ net141 vssd1 vssd1 vccd1 vccd1 _0384_ sky130_fd_sc_hd__inv_2
XANTENNA__3172__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3100_ clknet_leaf_29_clk _0090_ vssd1 vssd1 vccd1 vccd1 lcdPlayer.cnt_500hz\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_128_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3031_ clknet_leaf_10_clk clock_div.next_count\[11\] net214 vssd1 vssd1 vccd1 vccd1
+ clock_div.count\[11\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__2098__B2 net140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_128_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2117__B net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2270__A1 dispFSM.msg\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2815_ gamelogic.rights\[1\] gamelogic.rights\[0\] vssd1 vssd1 vccd1 vccd1 _1360_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_14_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3612__243 vssd1 vssd1 vccd1 vccd1 _3612__243/HI net243 sky130_fd_sc_hd__conb_1
X_2746_ _1296_ _1298_ _1299_ vssd1 vssd1 vccd1 vccd1 _1300_ sky130_fd_sc_hd__a21oi_1
X_2677_ gamelogic.setWord\[34\] _0379_ gamelogic.setWord\[35\] _0380_ vssd1 vssd1
+ vccd1 vccd1 _1243_ sky130_fd_sc_hd__a22o_1
XANTENNA__3515__CLK clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2573__A2 net114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1628_ net6 _0557_ _0561_ _0562_ vssd1 vssd1 vccd1 vccd1 _0563_ sky130_fd_sc_hd__a211o_1
XFILLER_0_1_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1559_ _0500_ _0506_ vssd1 vssd1 vccd1 vccd1 _0507_ sky130_fd_sc_hd__nand2_1
X_3229_ clknet_leaf_11_clk _0203_ net217 vssd1 vssd1 vccd1 vccd1 keypadFSMHost.prev_key\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_94_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3045__CLK clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_99_Left_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3195__CLK clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2043__A net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2189__S net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout94_X net94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3055__RESET_B _0017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_20_clk_A clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2600_ hostdisp.bottom\[44\] dispFSM.guesses\[20\] net227 vssd1 vssd1 vccd1 vccd1
+ _1174_ sky130_fd_sc_hd__mux2_1
X_3580_ net157 vssd1 vssd1 vccd1 vccd1 net12 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_82_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2531_ _0764_ _1105_ _1108_ vssd1 vssd1 vccd1 vccd1 _1109_ sky130_fd_sc_hd__or3_1
X_2462_ net343 net70 _1053_ _1029_ vssd1 vssd1 vccd1 vccd1 _0160_ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_35_clk_A clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1413_ keypadFSMHost.prev_key\[4\] vssd1 vssd1 vccd1 vccd1 _0367_ sky130_fd_sc_hd__inv_2
XFILLER_0_48_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2393_ net417 _1018_ net182 vssd1 vssd1 vccd1 vccd1 _1021_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_155_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3014_ net219 vssd1 vssd1 vccd1 vccd1 _0039_ sky130_fd_sc_hd__inv_2
XFILLER_0_64_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_175_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_175_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2562__S net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout141_A gamelogic.letter\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2729_ net365 keypadHostt.scan_col\[3\] _1287_ vssd1 vssd1 vccd1 vccd1 _0200_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout111 _1085_ vssd1 vssd1 vccd1 vccd1 net111 sky130_fd_sc_hd__buf_4
Xfanout100 net104 vssd1 vssd1 vccd1 vccd1 net100 sky130_fd_sc_hd__clkbuf_2
Xfanout122 _0858_ vssd1 vssd1 vccd1 vccd1 net122 sky130_fd_sc_hd__buf_2
Xfanout155 _0421_ vssd1 vssd1 vccd1 vccd1 net155 sky130_fd_sc_hd__buf_2
Xfanout133 hostdisp.Cstate vssd1 vssd1 vccd1 vccd1 net133 sky130_fd_sc_hd__buf_2
Xfanout144 gamelogic.letter\[1\] vssd1 vssd1 vccd1 vccd1 net144 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_148_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout199 net200 vssd1 vssd1 vccd1 vccd1 net199 sky130_fd_sc_hd__clkbuf_4
Xfanout188 net189 vssd1 vssd1 vccd1 vccd1 net188 sky130_fd_sc_hd__clkbuf_4
Xfanout177 net179 vssd1 vssd1 vccd1 vccd1 net177 sky130_fd_sc_hd__clkbuf_4
Xfanout166 net169 vssd1 vssd1 vccd1 vccd1 net166 sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_29_Right_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout54_A _1393_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_96_234 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_38_Right_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2537__A2 _1095_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_166_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_47_Right_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_189_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3210__CLK clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_125_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1962_ uart_receiver.bit_index\[2\] uart_receiver.bit_index\[0\] net149 vssd1 vssd1
+ vccd1 vccd1 _0801_ sky130_fd_sc_hd__or3b_1
XPHY_EDGE_ROW_56_Right_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_172_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1893_ uart_transmitter.clk_count\[9\] _0746_ vssd1 vssd1 vccd1 vccd1 _0748_ sky130_fd_sc_hd__nand2_1
XFILLER_0_28_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_44 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_136_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3563_ clknet_leaf_14_clk hostdisp.next_curr_guesses\[45\] net207 vssd1 vssd1 vccd1
+ vccd1 hostdisp.curr_guesses\[45\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_97_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2411__A _0828_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3494_ clknet_leaf_4_clk hostdisp.next_curr_word\[16\] net177 vssd1 vssd1 vccd1 vccd1
+ hostdisp.curr_word\[16\] sky130_fd_sc_hd__dfstp_1
X_2514_ dispFSM.guesses\[56\] net117 _1091_ _1077_ vssd1 vssd1 vccd1 vccd1 _1092_
+ sky130_fd_sc_hd__a211o_1
X_2445_ net130 host_message_reg.setLetter\[4\] hostdisp.curr_word\[20\] _0830_ _1034_
+ vssd1 vssd1 vccd1 vccd1 _1045_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_65_Right_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2376_ lcdPlayer.cnt_20ms\[12\] lcdPlayer.cnt_20ms\[11\] lcdPlayer.cnt_20ms\[10\]
+ _1004_ vssd1 vssd1 vccd1 vccd1 _1009_ sky130_fd_sc_hd__and4_1
XFILLER_0_75_63 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout189_A net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_267 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_166_Right_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_143_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_74_Right_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout144_X net144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_83_Right_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_113_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3383__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2455__B2 _0828_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_92_Right_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_133_Right_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_182_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_116_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2230_ gamelogic.state\[2\] _0814_ _0924_ vssd1 vssd1 vccd1 vccd1 _0925_ sky130_fd_sc_hd__o21ai_1
XANTENNA_clkbuf_2_2__f_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2161_ gamelogic.setWord\[23\] hostdisp.curr_guesses\[23\] net126 vssd1 vssd1 vccd1
+ vccd1 _0883_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_88_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2092_ hostdisp.curr_word\[25\] net101 _0850_ net144 vssd1 vssd1 vccd1 vccd1 hostdisp.next_curr_word\[25\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_177_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_64_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2994_ net222 vssd1 vssd1 vccd1 vccd1 _0019_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_100_Right_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1945_ _0789_ _0790_ _0185_ _0787_ vssd1 vssd1 vccd1 vccd1 _0791_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_28_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_134 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1957__A0 net2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1876_ uart_transmitter.clk_count\[3\] _0734_ vssd1 vssd1 vccd1 vccd1 _0737_ sky130_fd_sc_hd__or2_1
XFILLER_0_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3615_ net246 vssd1 vssd1 vccd1 vccd1 gpio_out[23] sky130_fd_sc_hd__buf_2
XANTENNA__3256__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3546_ clknet_leaf_1_clk hostdisp.next_curr_guesses\[28\] net176 vssd1 vssd1 vccd1
+ vccd1 hostdisp.curr_guesses\[28\] sky130_fd_sc_hd__dfstp_1
X_3477_ clknet_leaf_14_clk _0355_ net194 vssd1 vssd1 vccd1 vccd1 gamelogic.setWord\[39\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_50_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2134__A0 gamelogic.setWord\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2428_ hostdisp.curr_word\[11\] _0827_ vssd1 vssd1 vccd1 vccd1 _1037_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_4_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2359_ lcdPlayer.cnt_20ms\[6\] _0948_ _0953_ vssd1 vssd1 vccd1 vccd1 _0998_ sky130_fd_sc_hd__and3_1
XFILLER_0_193_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_145_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_163_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_35_Left_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_220 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_147 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3279__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1730_ uart_receiver.clk_count\[0\] _0642_ vssd1 vssd1 vccd1 vccd1 uart_receiver.next_clk_count\[0\]
+ sky130_fd_sc_hd__and2b_1
XFILLER_0_80_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1661_ _0443_ _0445_ _0589_ _0453_ keypadFSMPlayer.state\[4\] vssd1 vssd1 vccd1 vccd1
+ _0015_ sky130_fd_sc_hd__a32o_1
XFILLER_0_13_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_44_Left_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold208 hostdisp.curr_guesses\[27\] vssd1 vssd1 vccd1 vccd1 net472 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_150_150 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3400_ clknet_leaf_20_clk _0289_ net205 vssd1 vssd1 vccd1 vccd1 dispFSM.guesses\[54\]
+ sky130_fd_sc_hd__dfstp_1
Xhold219 dispFSM.guesses\[64\] vssd1 vssd1 vccd1 vccd1 net483 sky130_fd_sc_hd__dlygate4sd3_1
X_1592_ keypadFSMPlayer.unlocked net154 net128 vssd1 vssd1 vccd1 vccd1 _0535_ sky130_fd_sc_hd__and3_4
XFILLER_0_21_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3331_ clknet_leaf_3_clk _0220_ net172 vssd1 vssd1 vccd1 vccd1 gamelogic.indexCorrect\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_193_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3567__251 vssd1 vssd1 vccd1 vccd1 net251 _3567__251/LO sky130_fd_sc_hd__conb_1
X_3262_ clknet_leaf_2_clk hostdisp.nextBottom\[60\] net176 vssd1 vssd1 vccd1 vccd1
+ hostdisp.bottom\[60\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2213_ _0812_ _0908_ vssd1 vssd1 vccd1 vccd1 _0909_ sky130_fd_sc_hd__or2_2
X_3193_ clknet_leaf_29_clk _0169_ net181 vssd1 vssd1 vccd1 vccd1 hostdisp.top\[77\]
+ sky130_fd_sc_hd__dfrtp_1
X_2144_ gamelogic.setWord\[6\] _0874_ net136 vssd1 vssd1 vccd1 vccd1 hostdisp.nextBottom\[54\]
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_1_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_53_Left_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_163_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2075_ hostdisp.curr_word\[16\] net103 net75 _0843_ gamelogic.indexCorrect\[2\] vssd1
+ vssd1 vccd1 vccd1 _0844_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_88_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_158_272 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_140_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_114 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2977_ gamelogic.setWord\[16\] net53 net49 gamelogic.setWord\[24\] vssd1 vssd1 vccd1
+ vccd1 _0340_ sky130_fd_sc_hd__o22a_1
XFILLER_0_106_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_192_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout221_A net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_62_Left_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1928_ _0776_ vssd1 vssd1 vccd1 vccd1 _0186_ sky130_fd_sc_hd__inv_2
X_1859_ _0728_ _0729_ vssd1 vssd1 vccd1 vccd1 clock_div.next_count\[27\] sky130_fd_sc_hd__nor2_1
XFILLER_0_16_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_188_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_151_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1914__S _0764_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3529_ clknet_leaf_2_clk hostdisp.next_curr_guesses\[11\] net171 vssd1 vssd1 vccd1
+ vccd1 hostdisp.curr_guesses\[11\] sky130_fd_sc_hd__dfstp_1
XPHY_EDGE_ROW_71_Left_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3421__CLK clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_164_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_80_Left_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2594__B1 _1084_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold91 clock_div.count\[23\] vssd1 vssd1 vccd1 vccd1 net355 sky130_fd_sc_hd__dlygate4sd3_1
Xhold80 hostdisp.top\[70\] vssd1 vssd1 vccd1 vccd1 net344 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2508__X _1086_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_180_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2900_ dispFSM.guesses\[40\] net81 net56 net539 vssd1 vssd1 vccd1 vccd1 _0267_ sky130_fd_sc_hd__o22a_1
XFILLER_0_85_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2821__A1 net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2831_ _1368_ gamelogic.correct\[0\] _1366_ vssd1 vssd1 vccd1 vccd1 _0221_ sky130_fd_sc_hd__mux2_1
X_2762_ _0612_ _1293_ _1297_ vssd1 vssd1 vccd1 vccd1 _1315_ sky130_fd_sc_hd__and3b_1
XFILLER_0_155_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2243__X _0934_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_139 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_256 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1713_ _0628_ _0627_ vssd1 vssd1 vccd1 vccd1 _0629_ sky130_fd_sc_hd__and2b_1
XFILLER_0_170_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2693_ _0377_ gamelogic.setWord\[24\] _1257_ vssd1 vssd1 vccd1 vccd1 _1258_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_13_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1644_ keypadHostt.scan_col\[3\] _0366_ _0546_ _0567_ _0571_ vssd1 vssd1 vccd1 vccd1
+ _0579_ sky130_fd_sc_hd__a311o_1
XFILLER_0_123_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3402__SET_B net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1575_ _0468_ _0516_ vssd1 vssd1 vccd1 vccd1 _0522_ sky130_fd_sc_hd__xor2_1
XANTENNA__3465__SET_B net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3314_ clknet_leaf_35_clk uart_receiver.next_clk_count\[6\] net161 vssd1 vssd1 vccd1
+ vccd1 uart_receiver.clk_count\[6\] sky130_fd_sc_hd__dfrtp_1
X_3245_ clknet_leaf_3_clk hostdisp.nextBottom\[43\] net174 vssd1 vssd1 vccd1 vccd1
+ hostdisp.bottom\[43\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_174_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3176_ clknet_leaf_30_clk _0152_ net185 vssd1 vssd1 vccd1 vccd1 hostdisp.top\[60\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_178_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3444__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2127_ gamelogic.setWord\[6\] net124 vssd1 vssd1 vccd1 vccd1 _0866_ sky130_fd_sc_hd__or2_1
XFILLER_0_13_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout171_A net180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_37_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2058_ hostdisp.curr_word\[6\] net98 _0835_ gamelogic.letter\[6\] vssd1 vssd1 vccd1
+ vccd1 hostdisp.next_curr_word\[6\] sky130_fd_sc_hd__o22a_1
XFILLER_0_190_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_190_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3173__RESET_B net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout224_X net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2576__B1 _1086_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2040__A2 net94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout84_A _0940_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_160_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_109_Left_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2031__A2 net95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_318 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_118_Left_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3538__SET_B net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3030_ clknet_leaf_9_clk clock_div.next_count\[10\] net214 vssd1 vssd1 vccd1 vccd1
+ clock_div.count\[10\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__2098__A2 net96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_128_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_127_Left_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_175_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_9_clk_A clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_42_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2814_ _1359_ _1358_ gamelogic.rights\[0\] vssd1 vssd1 vccd1 vccd1 _0213_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_139_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2558__B1 net105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2745_ _0612_ _1296_ _1298_ vssd1 vssd1 vccd1 vccd1 _1299_ sky130_fd_sc_hd__nor3_1
XANTENNA__2022__A2 net92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_136_Left_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2676_ _0383_ net141 gamelogic.indexCorrect\[4\] _1239_ _1241_ vssd1 vssd1 vccd1
+ vccd1 _1242_ sky130_fd_sc_hd__a2111oi_2
XFILLER_0_78_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1627_ net3 _0541_ _0543_ _0552_ vssd1 vssd1 vccd1 vccd1 _0562_ sky130_fd_sc_hd__or4b_1
XFILLER_0_111_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1558_ net146 _0505_ _0427_ net229 net233 vssd1 vssd1 vccd1 vccd1 _0506_ sky130_fd_sc_hd__o2111ai_2
X_1489_ _0440_ vssd1 vssd1 vccd1 vccd1 _0441_ sky130_fd_sc_hd__inv_2
X_3228_ clknet_leaf_11_clk _0202_ net222 vssd1 vssd1 vccd1 vccd1 keypadFSMHost.prev_key\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_3159_ clknet_leaf_28_clk _0135_ net166 vssd1 vssd1 vccd1 vccd1 hostdisp.top\[43\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_178_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_34_clk clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_34_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_181_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_169_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3024__RESET_B net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_25_clk clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_25_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__2788__B1 net104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_48 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2521__X _1099_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2530_ _1057_ _1068_ _1069_ net108 _1107_ vssd1 vssd1 vccd1 vccd1 _1108_ sky130_fd_sc_hd__a32o_1
X_2461_ hostdisp.curr_word\[28\] _0827_ vssd1 vssd1 vccd1 vccd1 _1053_ sky130_fd_sc_hd__or2_1
X_1412_ keypadFSMHost.prev_key\[3\] vssd1 vssd1 vccd1 vccd1 _0366_ sky130_fd_sc_hd__inv_2
XFILLER_0_139_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2392_ lcdPlayer.cnt_20ms\[17\] _1018_ vssd1 vssd1 vccd1 vccd1 _1020_ sky130_fd_sc_hd__and2_1
XFILLER_0_47_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3013_ net222 vssd1 vssd1 vccd1 vccd1 _0038_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_147_Right_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_98 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_16_clk clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_16_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_171_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout134_A net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_171_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2728_ net376 net151 _1287_ vssd1 vssd1 vccd1 vccd1 _0199_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2659_ net105 _1229_ _1157_ vssd1 vssd1 vccd1 vccd1 _1230_ sky130_fd_sc_hd__a21o_1
XFILLER_0_1_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout112 _1080_ vssd1 vssd1 vccd1 vccd1 net112 sky130_fd_sc_hd__buf_4
Xfanout101 net104 vssd1 vssd1 vccd1 vccd1 net101 sky130_fd_sc_hd__buf_2
Xfanout134 net137 vssd1 vssd1 vccd1 vccd1 net134 sky130_fd_sc_hd__clkbuf_4
Xfanout123 net126 vssd1 vssd1 vccd1 vccd1 net123 sky130_fd_sc_hd__clkbuf_4
Xfanout156 net157 vssd1 vssd1 vccd1 vccd1 net156 sky130_fd_sc_hd__clkbuf_2
Xfanout145 gamelogic.letter\[0\] vssd1 vssd1 vccd1 vccd1 net145 sky130_fd_sc_hd__buf_4
XANTENNA__3521__SET_B net180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_148_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout167 net169 vssd1 vssd1 vccd1 vccd1 net167 sky130_fd_sc_hd__buf_2
Xfanout189 net190 vssd1 vssd1 vccd1 vccd1 net189 sky130_fd_sc_hd__clkbuf_2
Xfanout178 net179 vssd1 vssd1 vccd1 vccd1 net178 sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_114_Right_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_107_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout47_A net48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_139_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_159_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3162__CLK clknet_leaf_31_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_110 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_316 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2501__B net139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_166_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2473__A2 net75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3505__CLK clknet_leaf_31_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1961_ _0618_ _0800_ vssd1 vssd1 vccd1 vccd1 uart_receiver.temp_byte\[1\] sky130_fd_sc_hd__and2_1
X_1892_ uart_transmitter.clk_count\[9\] _0746_ vssd1 vssd1 vccd1 vccd1 _0747_ sky130_fd_sc_hd__or2_1
XFILLER_0_50_56 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3562_ clknet_leaf_1_clk hostdisp.next_curr_guesses\[44\] net175 vssd1 vssd1 vccd1
+ vccd1 hostdisp.curr_guesses\[44\] sky130_fd_sc_hd__dfstp_1
XFILLER_0_70_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2513_ dispFSM.guesses\[40\] net111 _1086_ dispFSM.guesses\[72\] _1090_ vssd1 vssd1
+ vccd1 vccd1 _1091_ sky130_fd_sc_hd__a221o_1
XFILLER_0_121_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2411__B net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3493_ clknet_leaf_30_clk hostdisp.next_curr_word\[15\] net185 vssd1 vssd1 vccd1
+ vccd1 hostdisp.curr_word\[15\] sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_5_clk clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_5_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_121_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2444_ net362 net67 _1044_ vssd1 vssd1 vccd1 vccd1 _0151_ sky130_fd_sc_hd__o21a_1
XFILLER_0_11_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3035__CLK clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2375_ _1008_ net168 _1007_ vssd1 vssd1 vccd1 vccd1 _0118_ sky130_fd_sc_hd__and3b_1
XFILLER_0_75_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_67_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3185__CLK clknet_leaf_30_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_182_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_143_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_163_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout137_X net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1975__A1 net2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1917__S _0764_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_154_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3528__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2455__A2 net71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_34_clk_A clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2612__C1 net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1966__A1 net2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_343 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2658__S net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2160_ gamelogic.setWord\[14\] _0882_ net134 vssd1 vssd1 vccd1 vccd1 hostdisp.nextBottom\[62\]
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_88_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2091_ hostdisp.curr_word\[24\] net101 _0850_ net145 vssd1 vssd1 vccd1 vccd1 hostdisp.next_curr_word\[24\]
+ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_183_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_100_Left_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_185_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2993_ net208 vssd1 vssd1 vccd1 vccd1 _0018_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_148 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1944_ net166 _0765_ _0770_ _0185_ vssd1 vssd1 vccd1 vccd1 _0790_ sky130_fd_sc_hd__a31o_1
X_3614_ net245 vssd1 vssd1 vccd1 vccd1 gpio_out[22] sky130_fd_sc_hd__buf_2
X_1875_ uart_transmitter.clk_count\[3\] _0734_ vssd1 vssd1 vccd1 vccd1 _0736_ sky130_fd_sc_hd__and2_1
XFILLER_0_153_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_146 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2422__A net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3545_ clknet_leaf_0_clk hostdisp.next_curr_guesses\[27\] net170 vssd1 vssd1 vccd1
+ vccd1 hostdisp.curr_guesses\[27\] sky130_fd_sc_hd__dfstp_1
X_3476_ clknet_leaf_6_clk _0354_ net192 vssd1 vssd1 vccd1 vccd1 gamelogic.setWord\[38\]
+ sky130_fd_sc_hd__dfstp_1
X_2427_ net337 net70 _1036_ _0828_ vssd1 vssd1 vccd1 vccd1 _0142_ sky130_fd_sc_hd__a22o_1
XFILLER_0_43_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_96 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2358_ _0358_ _0947_ _0997_ _0017_ vssd1 vssd1 vccd1 vccd1 _0112_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_193_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2289_ net276 net74 vssd1 vssd1 vccd1 vccd1 _0083_ sky130_fd_sc_hd__nor2_1
XFILLER_0_193_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_218 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_191_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3350__CLK clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2676__A2 net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_163_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_26_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_232 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_174_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1660_ keypadFSMPlayer.state\[5\] keypadFSMPlayer.state\[2\] keypadFSMPlayer.state\[3\]
+ keypadFSMPlayer.state\[1\] vssd1 vssd1 vccd1 vccd1 _0589_ sky130_fd_sc_hd__or4_1
XANTENNA__2242__A _0360_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1591_ _0519_ _0533_ _0534_ _0454_ dispFSM.msg\[0\] vssd1 vssd1 vccd1 vccd1 _0058_
+ sky130_fd_sc_hd__o32a_1
XTAP_TAPCELL_ROW_133_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold209 dispFSM.guesses\[76\] vssd1 vssd1 vccd1 vccd1 net473 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_150_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3330_ clknet_leaf_35_clk _0219_ net161 vssd1 vssd1 vccd1 vccd1 gamelogic.red sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3261_ clknet_leaf_2_clk hostdisp.nextBottom\[59\] net170 vssd1 vssd1 vccd1 vccd1
+ hostdisp.bottom\[59\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_186_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2212_ gamelogic.state\[0\] gamelogic.state\[1\] vssd1 vssd1 vccd1 vccd1 _0908_ sky130_fd_sc_hd__nand2_1
X_3192_ clknet_leaf_31_clk _0168_ net172 vssd1 vssd1 vccd1 vccd1 hostdisp.top\[76\]
+ sky130_fd_sc_hd__dfrtp_1
X_2143_ gamelogic.setWord\[14\] hostdisp.curr_guesses\[14\] net124 vssd1 vssd1 vccd1
+ vccd1 _0874_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_1_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2074_ hostdisp.curr_word\[17\] hostdisp.curr_word\[19\] hostdisp.curr_word\[20\]
+ _0409_ net103 vssd1 vssd1 vccd1 vccd1 _0843_ sky130_fd_sc_hd__a41o_1
XANTENNA__2419__A2 _1031_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_284 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2976_ gamelogic.setWord\[15\] net55 _1394_ gamelogic.setWord\[23\] vssd1 vssd1 vccd1
+ vccd1 _0339_ sky130_fd_sc_hd__a22o_1
XFILLER_0_8_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1927_ net181 _0775_ vssd1 vssd1 vccd1 vccd1 _0776_ sky130_fd_sc_hd__nand2_2
XANTENNA_fanout214_A net218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1858_ clock_div.count\[27\] clock_div.count\[26\] _0727_ vssd1 vssd1 vccd1 vccd1
+ _0729_ sky130_fd_sc_hd__and3_1
XFILLER_0_126_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_188_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_151_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1789_ _0682_ _0683_ _0684_ _0686_ vssd1 vssd1 vccd1 vccd1 _0687_ sky130_fd_sc_hd__or4_1
XFILLER_0_12_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3528_ clknet_leaf_2_clk hostdisp.next_curr_guesses\[10\] net175 vssd1 vssd1 vccd1
+ vccd1 hostdisp.curr_guesses\[10\] sky130_fd_sc_hd__dfstp_1
X_3459_ clknet_leaf_13_clk _0337_ net198 vssd1 vssd1 vccd1 vccd1 gamelogic.setWord\[21\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__2107__B2 net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2997__A net221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1406__A net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2649__A2 net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold81 hostdisp.curr_guesses\[7\] vssd1 vssd1 vccd1 vccd1 net345 sky130_fd_sc_hd__dlygate4sd3_1
Xhold92 hostdisp.top\[60\] vssd1 vssd1 vccd1 vccd1 net356 sky130_fd_sc_hd__dlygate4sd3_1
Xhold70 hostdisp.top\[51\] vssd1 vssd1 vccd1 vccd1 net334 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_187_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_180_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3246__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2806__C1 gamelogic.indexCorrect\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2830_ gamelogic.correct\[0\] gamelogic.rights\[0\] _1367_ vssd1 vssd1 vccd1 vccd1
+ _1368_ sky130_fd_sc_hd__a21oi_1
XANTENNA__3396__CLK clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2761_ _1306_ _1313_ _0560_ vssd1 vssd1 vccd1 vccd1 _1314_ sky130_fd_sc_hd__a21boi_1
XANTENNA__2034__B1 net79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2692_ _0384_ gamelogic.setWord\[29\] gamelogic.setWord\[31\] _0386_ vssd1 vssd1
+ vccd1 vccd1 _1257_ sky130_fd_sc_hd__a22o_1
XFILLER_0_13_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1712_ uart_receiver.state\[2\] _0396_ uart_receiver.state\[1\] vssd1 vssd1 vccd1
+ vccd1 _0628_ sky130_fd_sc_hd__or3_1
XANTENNA__2585__B2 net108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2585__A1 net139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1643_ keypadFSMHost.prev_key\[7\] _0560_ vssd1 vssd1 vccd1 vccd1 _0578_ sky130_fd_sc_hd__xor2_1
XFILLER_0_170_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_1 gamelogic.letter\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1574_ dispFSM.msg\[3\] _0447_ vssd1 vssd1 vccd1 vccd1 _0521_ sky130_fd_sc_hd__and2_1
XANTENNA__2700__A net140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3313_ clknet_leaf_35_clk uart_receiver.next_clk_count\[5\] net161 vssd1 vssd1 vccd1
+ vccd1 uart_receiver.clk_count\[5\] sky130_fd_sc_hd__dfrtp_1
X_3244_ clknet_leaf_3_clk hostdisp.nextBottom\[42\] net174 vssd1 vssd1 vccd1 vccd1
+ hostdisp.bottom\[42\] sky130_fd_sc_hd__dfrtp_1
X_3175_ clknet_leaf_22_clk _0151_ net185 vssd1 vssd1 vccd1 vccd1 hostdisp.top\[59\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_174_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2126_ net130 _0865_ vssd1 vssd1 vccd1 vccd1 hostdisp.nextBottom\[45\] sky130_fd_sc_hd__or2_1
XFILLER_0_178_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_37_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout164_A net165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2057_ hostdisp.curr_word\[5\] net96 _0836_ net141 vssd1 vssd1 vccd1 vccd1 hostdisp.next_curr_word\[5\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_193_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_193_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_146_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2959_ host_message_reg.setLetter\[6\] net53 net49 gamelogic.setWord\[6\] vssd1 vssd1
+ vccd1 vccd1 _0322_ sky130_fd_sc_hd__o22a_1
XANTENNA__2025__B1 net80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout217_X net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_335 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout77_A _0826_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_169_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_108 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_171 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2016__B1 net79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_128_Right_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_169_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2007__B1 net80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2813_ _1358_ _0929_ _0909_ vssd1 vssd1 vccd1 vccd1 _1359_ sky130_fd_sc_hd__and3b_1
XFILLER_0_183_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2744_ _0612_ _1293_ _1297_ vssd1 vssd1 vccd1 vccd1 _1298_ sky130_fd_sc_hd__nor3_1
XFILLER_0_143_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_139_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2675_ _0376_ net145 gamelogic.setWord\[36\] _0382_ _1240_ vssd1 vssd1 vccd1 vccd1
+ _1241_ sky130_fd_sc_hd__a221o_1
X_1626_ net153 _0548_ _0557_ _0559_ vssd1 vssd1 vccd1 vccd1 _0561_ sky130_fd_sc_hd__o22a_1
XFILLER_0_78_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1557_ net147 _0461_ vssd1 vssd1 vccd1 vccd1 _0505_ sky130_fd_sc_hd__nor2_1
XFILLER_0_1_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2730__A1 net3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1488_ net148 keypadplayer.scan_col\[0\] net146 net147 vssd1 vssd1 vccd1 vccd1 _0440_
+ sky130_fd_sc_hd__or4b_2
XFILLER_0_94_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3227_ clknet_leaf_16_clk _0201_ net222 vssd1 vssd1 vccd1 vccd1 keypadFSMHost.prev_key\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_94_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3158_ clknet_leaf_31_clk _0134_ net163 vssd1 vssd1 vccd1 vccd1 hostdisp.top\[42\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_178_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2109_ net403 net96 _0856_ net141 vssd1 vssd1 vccd1 vccd1 hostdisp.next_curr_word\[37\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_178_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3089_ clknet_leaf_19_clk _0079_ net211 vssd1 vssd1 vccd1 vccd1 message_reg.msg\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_193_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_180_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2960__A1 host_message_reg.setLetter\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2460_ hostdisp.curr_word\[27\] net75 net71 net371 _1034_ vssd1 vssd1 vccd1 vccd1
+ _0159_ sky130_fd_sc_hd__a221o_1
X_1411_ gamelogic.state\[3\] vssd1 vssd1 vccd1 vccd1 _0365_ sky130_fd_sc_hd__inv_2
XFILLER_0_139_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2391_ _1018_ _1019_ vssd1 vssd1 vccd1 vccd1 _0123_ sky130_fd_sc_hd__nor2_1
X_3012_ net220 vssd1 vssd1 vccd1 vccd1 _0037_ sky130_fd_sc_hd__inv_2
XFILLER_0_155_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2476__B1 net69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_175_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2779__A1 host_message_reg.setLetter\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_306 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2727_ net360 net152 _1287_ vssd1 vssd1 vccd1 vccd1 _0198_ sky130_fd_sc_hd__mux2_1
XFILLER_0_171_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_189_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2658_ hostdisp.bottom\[47\] dispFSM.guesses\[23\] net228 vssd1 vssd1 vccd1 vccd1
+ _1229_ sky130_fd_sc_hd__mux2_1
X_1609_ net229 net3 vssd1 vssd1 vccd1 vccd1 _0544_ sky130_fd_sc_hd__and2b_1
XANTENNA__2703__A1 gamelogic.letter\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2589_ hostdisp.bottom\[52\] net115 net109 hostdisp.bottom\[60\] vssd1 vssd1 vccd1
+ vccd1 _1163_ sky130_fd_sc_hd__a22o_1
Xfanout102 net104 vssd1 vssd1 vccd1 vccd1 net102 sky130_fd_sc_hd__buf_2
XFILLER_0_1_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout113 _1080_ vssd1 vssd1 vccd1 vccd1 net113 sky130_fd_sc_hd__buf_2
Xfanout146 keypadplayer.scan_col\[3\] vssd1 vssd1 vccd1 vccd1 net146 sky130_fd_sc_hd__buf_2
Xfanout135 net137 vssd1 vssd1 vccd1 vccd1 net135 sky130_fd_sc_hd__buf_2
Xfanout124 net125 vssd1 vssd1 vccd1 vccd1 net124 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_148_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input1_A en vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout157 net24 vssd1 vssd1 vccd1 vccd1 net157 sky130_fd_sc_hd__clkbuf_2
Xfanout168 net169 vssd1 vssd1 vccd1 vccd1 net168 sky130_fd_sc_hd__buf_1
Xfanout179 net180 vssd1 vssd1 vccd1 vccd1 net179 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_107_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3307__CLK clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_159_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_181_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_122 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_155 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_328 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2942__A1 dispFSM.msg\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_155_Left_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_8_clk_A clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_166_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_164_Left_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_141_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1960_ net2 buffer.Rx_byte\[1\] _0799_ vssd1 vssd1 vccd1 vccd1 _0800_ sky130_fd_sc_hd__mux2_1
X_1891_ _0746_ net116 _0745_ vssd1 vssd1 vccd1 vccd1 uart_transmitter.next_clk_count\[8\]
+ sky130_fd_sc_hd__and3b_1
XFILLER_0_141_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_136_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3561_ clknet_leaf_0_clk hostdisp.next_curr_guesses\[43\] net170 vssd1 vssd1 vccd1
+ vccd1 hostdisp.curr_guesses\[43\] sky130_fd_sc_hd__dfstp_1
XPHY_EDGE_ROW_180_Right_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2512_ dispFSM.guesses\[0\] _1084_ net109 dispFSM.guesses\[32\] vssd1 vssd1 vccd1
+ vccd1 _1090_ sky130_fd_sc_hd__a22o_1
XFILLER_0_11_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3492_ clknet_leaf_30_clk hostdisp.next_curr_word\[14\] net174 vssd1 vssd1 vccd1
+ vccd1 hostdisp.curr_word\[14\] sky130_fd_sc_hd__dfstp_1
XPHY_EDGE_ROW_173_Left_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2443_ net129 host_message_reg.setLetter\[3\] _1029_ _1043_ net70 vssd1 vssd1 vccd1
+ vccd1 _1044_ sky130_fd_sc_hd__a221o_1
X_2374_ lcdPlayer.cnt_20ms\[11\] lcdPlayer.cnt_20ms\[10\] _1004_ vssd1 vssd1 vccd1
+ vccd1 _1008_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_67_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_182_Left_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_148_168 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_154_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_191_Left_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2688__B1 gamelogic.setWord\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input4_X net4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2860__A0 net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2679__B1 gamelogic.setWord\[39\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2090_ _0850_ vssd1 vssd1 vccd1 vccd1 _0851_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_88_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_183_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2992_ gamelogic.setWord\[31\] net55 _1394_ gamelogic.setWord\[39\] vssd1 vssd1 vccd1
+ vccd1 _0355_ sky130_fd_sc_hd__a22o_1
XFILLER_0_28_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1943_ _0183_ _0182_ vssd1 vssd1 vccd1 vccd1 _0789_ sky130_fd_sc_hd__nor2_1
XFILLER_0_28_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3613_ net244 vssd1 vssd1 vccd1 vccd1 gpio_out[21] sky130_fd_sc_hd__buf_2
X_1874_ _0734_ _0735_ net116 vssd1 vssd1 vccd1 vccd1 uart_transmitter.next_clk_count\[2\]
+ sky130_fd_sc_hd__and3b_1
XFILLER_0_126_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_153_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_141_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2422__B _0822_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3544_ clknet_leaf_1_clk hostdisp.next_curr_guesses\[26\] net175 vssd1 vssd1 vccd1
+ vccd1 hostdisp.curr_guesses\[26\] sky130_fd_sc_hd__dfstp_1
X_3475_ clknet_leaf_14_clk _0353_ net199 vssd1 vssd1 vccd1 vccd1 gamelogic.setWord\[37\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_177_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2426_ hostdisp.curr_word\[10\] net119 vssd1 vssd1 vccd1 vccd1 _1036_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout194_A net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2357_ _0948_ _0953_ vssd1 vssd1 vccd1 vccd1 _0997_ sky130_fd_sc_hd__and2_1
X_2288_ net106 _0955_ vssd1 vssd1 vccd1 vccd1 _0957_ sky130_fd_sc_hd__nand2b_1
XANTENNA__3167__RESET_B net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_176_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_104_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2172__X hostdisp.nextBottom\[68\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_191_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3590__262 vssd1 vssd1 vccd1 vccd1 net262 _3590__262/LO sky130_fd_sc_hd__conb_1
XANTENNA__2070__B2 net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_182 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2358__C1 _0017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3217__Q gamelogic.indexCorrect\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_174_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_182_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2242__B _0693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1590_ dispFSM.msg\[0\] _0447_ vssd1 vssd1 vccd1 vccd1 _0534_ sky130_fd_sc_hd__and2_1
XANTENNA__3175__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2116__A2 net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3260_ clknet_leaf_3_clk hostdisp.nextBottom\[58\] net178 vssd1 vssd1 vccd1 vccd1
+ hostdisp.bottom\[58\] sky130_fd_sc_hd__dfrtp_1
X_2211_ _0607_ net97 net135 vssd1 vssd1 vccd1 vccd1 hostdisp.next_state sky130_fd_sc_hd__mux2_1
X_3191_ clknet_leaf_31_clk _0167_ net172 vssd1 vssd1 vccd1 vccd1 hostdisp.top\[75\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_179_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2142_ net534 _0873_ net136 vssd1 vssd1 vccd1 vccd1 hostdisp.nextBottom\[53\] sky130_fd_sc_hd__mux2_1
X_2073_ hostdisp.curr_word\[18\] _0408_ hostdisp.curr_word\[22\] net103 vssd1 vssd1
+ vccd1 vccd1 _0842_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_1_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_66 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_173_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_161_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2975_ gamelogic.setWord\[14\] net53 net49 gamelogic.setWord\[22\] vssd1 vssd1 vccd1
+ vccd1 _0338_ sky130_fd_sc_hd__o22a_1
XFILLER_0_44_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3518__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1926_ lcdPlayer.nextState\[4\] lcdPlayer.currentState\[4\] _0764_ vssd1 vssd1 vccd1
+ vccd1 _0775_ sky130_fd_sc_hd__mux2_1
X_1857_ clock_div.count\[26\] _0727_ net440 vssd1 vssd1 vccd1 vccd1 _0728_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_21_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_188_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_151_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1788_ clock_div.count\[14\] clock_div.count\[17\] _0685_ vssd1 vssd1 vccd1 vccd1
+ _0686_ sky130_fd_sc_hd__or3b_1
X_3527_ clknet_leaf_5_clk hostdisp.next_curr_guesses\[9\] net197 vssd1 vssd1 vccd1
+ vccd1 hostdisp.curr_guesses\[9\] sky130_fd_sc_hd__dfstp_1
XANTENNA__2579__S net226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3458_ clknet_leaf_1_clk _0336_ net176 vssd1 vssd1 vccd1 vccd1 gamelogic.setWord\[20\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA_clkbuf_leaf_33_clk_A clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3389_ clknet_leaf_25_clk _0278_ net183 vssd1 vssd1 vccd1 vccd1 dispFSM.guesses\[43\]
+ sky130_fd_sc_hd__dfstp_1
X_2409_ _0829_ _0857_ vssd1 vssd1 vccd1 vccd1 _1029_ sky130_fd_sc_hd__nor2_2
XFILLER_0_39_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_83_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3048__CLK clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_109_Right_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2594__A2 net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold71 hostdisp.curr_guesses\[5\] vssd1 vssd1 vccd1 vccd1 net335 sky130_fd_sc_hd__dlygate4sd3_1
Xhold60 message_reg.msg\[7\] vssd1 vssd1 vccd1 vccd1 net324 sky130_fd_sc_hd__dlygate4sd3_1
Xhold82 hostdisp.next_curr_guesses\[7\] vssd1 vssd1 vccd1 vccd1 net346 sky130_fd_sc_hd__dlygate4sd3_1
Xhold93 hostdisp.top\[101\] vssd1 vssd1 vccd1 vccd1 net357 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_170_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2760_ _0540_ _0547_ vssd1 vssd1 vccd1 vccd1 _1313_ sky130_fd_sc_hd__nand2_1
XFILLER_0_155_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2034__A1 net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2691_ _0386_ gamelogic.setWord\[31\] _0388_ _1254_ _1255_ vssd1 vssd1 vccd1 vccd1
+ _1256_ sky130_fd_sc_hd__o2111a_1
X_1711_ net2 net100 host_message_reg.Cstate vssd1 vssd1 vccd1 vccd1 _0627_ sky130_fd_sc_hd__or3b_1
X_1642_ _0573_ _0574_ _0575_ _0576_ vssd1 vssd1 vccd1 vccd1 _0577_ sky130_fd_sc_hd__or4_1
XFILLER_0_53_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1573_ dispFSM.msg\[4\] _0454_ _0518_ _0520_ vssd1 vssd1 vccd1 vccd1 _0062_ sky130_fd_sc_hd__o22a_1
XFILLER_0_21_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3312_ clknet_leaf_35_clk uart_receiver.next_clk_count\[4\] net161 vssd1 vssd1 vccd1
+ vccd1 uart_receiver.clk_count\[4\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3243_ clknet_leaf_14_clk hostdisp.nextBottom\[41\] net199 vssd1 vssd1 vccd1 vccd1
+ hostdisp.bottom\[41\] sky130_fd_sc_hd__dfrtp_1
X_3174_ clknet_leaf_22_clk _0150_ net201 vssd1 vssd1 vccd1 vccd1 hostdisp.top\[58\]
+ sky130_fd_sc_hd__dfrtp_1
X_2125_ gamelogic.setWord\[5\] hostdisp.curr_guesses\[5\] net125 vssd1 vssd1 vccd1
+ vccd1 _0865_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_37_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2056_ hostdisp.curr_word\[4\] net98 _0835_ net142 vssd1 vssd1 vccd1 vccd1 hostdisp.next_curr_word\[4\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_88_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_190_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_101_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3340__CLK clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2958_ host_message_reg.setLetter\[5\] net55 _1394_ net534 vssd1 vssd1 vccd1 vccd1
+ _0321_ sky130_fd_sc_hd__a22o_1
XFILLER_0_8_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_20_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1909_ lcdPlayer.cnt_500hz\[11\] lcdPlayer.cnt_500hz\[10\] vssd1 vssd1 vccd1 vccd1
+ _0762_ sky130_fd_sc_hd__nand2_1
XANTENNA__2576__A2 _1084_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2889_ dispFSM.guesses\[29\] net90 net64 net395 vssd1 vssd1 vccd1 vccd1 _0256_ sky130_fd_sc_hd__a22o_1
XANTENNA__3490__CLK clknet_leaf_30_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout112_X net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_347 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_286 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_160_291 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_169_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2519__Y _1097_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_187_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2812_ _1342_ _1356_ _1357_ vssd1 vssd1 vccd1 vccd1 _1358_ sky130_fd_sc_hd__nand3b_2
X_2743_ _0369_ _1397_ _1294_ keypadFSMHost.state\[2\] keypadFSMHost.state\[3\] vssd1
+ vssd1 vccd1 vccd1 _1297_ sky130_fd_sc_hd__a311o_1
XFILLER_0_143_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2558__A2 _1078_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_139_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2674_ gamelogic.setWord\[32\] _0377_ _1237_ _1238_ vssd1 vssd1 vccd1 vccd1 _1240_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_111_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1625_ _0542_ _0545_ _0552_ _0539_ vssd1 vssd1 vccd1 vccd1 _0560_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_111_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1556_ _0496_ _0503_ _0502_ vssd1 vssd1 vccd1 vccd1 _0504_ sky130_fd_sc_hd__o21a_1
XFILLER_0_111_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1487_ _0426_ _0438_ vssd1 vssd1 vccd1 vccd1 _0439_ sky130_fd_sc_hd__nor2_1
XANTENNA_clkload11_A clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3226_ clknet_leaf_11_clk _0200_ net216 vssd1 vssd1 vccd1 vccd1 keypadFSMHost.prev_key\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_3157_ clknet_leaf_28_clk _0133_ net166 vssd1 vssd1 vccd1 vccd1 hostdisp.top\[41\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_94_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_178_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2108_ hostdisp.curr_word\[36\] net99 _0855_ net142 vssd1 vssd1 vccd1 vccd1 hostdisp.next_curr_word\[36\]
+ sky130_fd_sc_hd__o22a_1
X_3088_ clknet_leaf_18_clk _0078_ net219 vssd1 vssd1 vccd1 vccd1 message_reg.msg\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_193_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2039_ net141 net95 net80 net401 vssd1 vssd1 vccd1 vccd1 hostdisp.next_curr_guesses\[45\]
+ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_59_Left_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_193_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2549__A2 net106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_157_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_68_Left_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2721__A2 gamelogic.setWord\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_77_Left_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_169_188 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_161_Right_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_172_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_86_Left_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2531__A _0764_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1410_ gamelogic.state\[0\] vssd1 vssd1 vccd1 vccd1 _0364_ sky130_fd_sc_hd__inv_2
XANTENNA__2173__A0 gamelogic.setWord\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2390_ net418 _1017_ net168 vssd1 vssd1 vccd1 vccd1 _1019_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_3_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3011_ net223 vssd1 vssd1 vccd1 vccd1 _0036_ sky130_fd_sc_hd__inv_2
XFILLER_0_161_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_175_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_175_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_171_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_190_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3259__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2726_ net408 keypadHostt.scan_col\[0\] _1287_ vssd1 vssd1 vccd1 vccd1 _0197_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2657_ _1224_ _1225_ _1227_ vssd1 vssd1 vccd1 vccd1 _1228_ sky130_fd_sc_hd__or3_1
XFILLER_0_124_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_189_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1608_ net229 net4 vssd1 vssd1 vccd1 vccd1 _0543_ sky130_fd_sc_hd__and2b_1
XFILLER_0_1_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout103 net104 vssd1 vssd1 vccd1 vccd1 net103 sky130_fd_sc_hd__buf_2
X_2588_ hostdisp.bottom\[76\] net112 _1096_ hostdisp.top\[68\] vssd1 vssd1 vccd1 vccd1
+ _1162_ sky130_fd_sc_hd__a22o_1
Xfanout147 keypadplayer.scan_col\[2\] vssd1 vssd1 vccd1 vccd1 net147 sky130_fd_sc_hd__buf_2
X_1539_ _0484_ _0485_ _0478_ _0480_ vssd1 vssd1 vccd1 vccd1 _0487_ sky130_fd_sc_hd__o211a_1
Xfanout136 net137 vssd1 vssd1 vccd1 vccd1 net136 sky130_fd_sc_hd__clkbuf_4
Xfanout125 net126 vssd1 vssd1 vccd1 vccd1 net125 sky130_fd_sc_hd__clkbuf_4
Xfanout114 _1076_ vssd1 vssd1 vccd1 vccd1 net114 sky130_fd_sc_hd__buf_4
Xfanout158 net160 vssd1 vssd1 vccd1 vccd1 net158 sky130_fd_sc_hd__clkbuf_4
Xfanout169 net225 vssd1 vssd1 vccd1 vccd1 net169 sky130_fd_sc_hd__clkbuf_2
X_3209_ clknet_leaf_29_clk _0185_ vssd1 vssd1 vccd1 vccd1 lcdPlayer.currentState\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_107_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1520__A net6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_159_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout92_X net92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold190 gamelogic.incorrect\[2\] vssd1 vssd1 vccd1 vccd1 net454 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_16_Right_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1430__A net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_177_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1969__A0 net2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1890_ uart_transmitter.clk_count\[8\] uart_transmitter.clk_count\[7\] _0742_ vssd1
+ vssd1 vccd1 vccd1 _0746_ sky130_fd_sc_hd__and3_1
XANTENNA__3285__RESET_B net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_178 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_25_Right_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3560_ clknet_leaf_0_clk hostdisp.next_curr_guesses\[42\] net175 vssd1 vssd1 vccd1
+ vccd1 hostdisp.curr_guesses\[42\] sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_136_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3551__CLK clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2511_ dispFSM.guesses\[16\] net105 _1088_ _0360_ vssd1 vssd1 vccd1 vccd1 _1089_
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_11_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3491_ clknet_leaf_30_clk hostdisp.next_curr_word\[13\] net185 vssd1 vssd1 vccd1
+ vccd1 hostdisp.curr_word\[13\] sky130_fd_sc_hd__dfrtp_1
X_2442_ hostdisp.curr_word\[19\] _0827_ vssd1 vssd1 vccd1 vccd1 _1043_ sky130_fd_sc_hd__or2_1
X_2373_ lcdPlayer.cnt_20ms\[10\] _1004_ lcdPlayer.cnt_20ms\[11\] vssd1 vssd1 vccd1
+ vccd1 _1007_ sky130_fd_sc_hd__a21o_1
XFILLER_0_75_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_33 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_34_Right_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_67_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2723__X _1286_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3081__CLK clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_50_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_43_Right_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_171_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_154_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2709_ _0382_ gamelogic.setWord\[20\] _1271_ _1272_ gamelogic.indexCorrect\[2\] vssd1
+ vssd1 vccd1 vccd1 _1273_ sky130_fd_sc_hd__a221o_1
XFILLER_0_112_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_7_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_52_Right_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_58_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout52_A _1393_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_61_Right_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_150 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_70_Right_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1425__A gamelogic.letter\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_88_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_183_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_48 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_142_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2991_ gamelogic.setWord\[30\] net52 net48 gamelogic.setWord\[38\] vssd1 vssd1 vccd1
+ vccd1 _0354_ sky130_fd_sc_hd__o22a_1
XFILLER_0_145_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1942_ _0776_ _0182_ vssd1 vssd1 vccd1 vccd1 _0788_ sky130_fd_sc_hd__nand2_1
X_1873_ uart_transmitter.clk_count\[0\] uart_transmitter.clk_count\[1\] uart_transmitter.clk_count\[2\]
+ vssd1 vssd1 vccd1 vccd1 _0735_ sky130_fd_sc_hd__a21o_1
XFILLER_0_124_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3612_ net243 vssd1 vssd1 vccd1 vccd1 gpio_out[20] sky130_fd_sc_hd__buf_2
XFILLER_0_153_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3543_ clknet_leaf_7_clk hostdisp.next_curr_guesses\[25\] net200 vssd1 vssd1 vccd1
+ vccd1 hostdisp.curr_guesses\[25\] sky130_fd_sc_hd__dfstp_1
XFILLER_0_51_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3474_ clknet_leaf_6_clk _0352_ net192 vssd1 vssd1 vccd1 vccd1 gamelogic.setWord\[36\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_10_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2425_ net383 net70 _1035_ _1029_ vssd1 vssd1 vccd1 vccd1 _0141_ sky130_fd_sc_hd__a22o_1
XFILLER_0_86_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2356_ net167 _0947_ _0996_ _0955_ vssd1 vssd1 vccd1 vccd1 _0111_ sky130_fd_sc_hd__a31o_1
X_2287_ net106 _0955_ vssd1 vssd1 vccd1 vccd1 _0956_ sky130_fd_sc_hd__and2b_1
XFILLER_0_29_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_191_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout142_X net142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2070__A2 net96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_7_clk_A clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_334 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1581__B2 dispFSM.msg\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2530__B1 net108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3233__Q host_message_reg.setLetter\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2804__A net142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_174_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2597__B1 net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1572__A1 dispFSM.msg\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2210_ net133 hostdisp.curr_guesses\[47\] net123 _0907_ vssd1 vssd1 vccd1 vccd1 hostdisp.nextBottom\[87\]
+ sky130_fd_sc_hd__a31o_1
XPHY_EDGE_ROW_13_Left_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3190_ clknet_leaf_31_clk _0166_ net172 vssd1 vssd1 vccd1 vccd1 hostdisp.top\[74\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__2521__B1 _1098_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2141_ gamelogic.setWord\[13\] hostdisp.curr_guesses\[13\] net125 vssd1 vssd1 vccd1
+ vccd1 _0873_ sky130_fd_sc_hd__mux2_1
X_2072_ net560 net96 _0841_ gamelogic.letter\[7\] vssd1 vssd1 vccd1 vccd1 hostdisp.next_curr_word\[15\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_158_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_22_Left_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2974_ net569 _1392_ _1394_ gamelogic.setWord\[21\] vssd1 vssd1 vccd1 vccd1 _0337_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__2714__A net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2588__B1 _1096_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1925_ lcdPlayer.nextState\[3\] _0764_ _0774_ net181 vssd1 vssd1 vccd1 vccd1 _0185_
+ sky130_fd_sc_hd__o211a_2
X_1856_ net363 _0727_ vssd1 vssd1 vccd1 vccd1 clock_div.next_count\[26\] sky130_fd_sc_hd__xor2_1
X_1787_ clock_div.count\[15\] clock_div.count\[16\] vssd1 vssd1 vccd1 vccd1 _0685_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_97_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_151_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3526_ clknet_leaf_7_clk hostdisp.next_curr_guesses\[8\] net196 vssd1 vssd1 vccd1
+ vccd1 hostdisp.curr_guesses\[8\] sky130_fd_sc_hd__dfstp_1
XFILLER_0_97_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout102_A net104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_31_Left_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3457_ clknet_leaf_1_clk _0335_ net176 vssd1 vssd1 vccd1 vccd1 gamelogic.setWord\[19\]
+ sky130_fd_sc_hd__dfstp_1
X_2408_ _0423_ net146 _0934_ vssd1 vssd1 vccd1 vccd1 _0131_ sky130_fd_sc_hd__mux2_1
X_3388_ clknet_leaf_24_clk _0277_ net189 vssd1 vssd1 vccd1 vccd1 dispFSM.guesses\[42\]
+ sky130_fd_sc_hd__dfstp_1
X_2339_ _0988_ _0956_ _0987_ vssd1 vssd1 vccd1 vccd1 _0102_ sky130_fd_sc_hd__and3b_1
XANTENNA__2512__B1 net109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_118 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_2_Right_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_162_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_40_Left_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold50 hostdisp.top\[56\] vssd1 vssd1 vccd1 vccd1 net314 sky130_fd_sc_hd__dlygate4sd3_1
Xhold72 hostdisp.next_curr_guesses\[5\] vssd1 vssd1 vccd1 vccd1 net336 sky130_fd_sc_hd__dlygate4sd3_1
Xhold61 hostdisp.top\[61\] vssd1 vssd1 vccd1 vccd1 net325 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold83 hostdisp.top\[55\] vssd1 vssd1 vccd1 vccd1 net347 sky130_fd_sc_hd__dlygate4sd3_1
Xhold94 lcdPlayer.cnt_20ms\[9\] vssd1 vssd1 vccd1 vccd1 net358 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2518__B net139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_187_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2806__A1 gamelogic.letter\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2034__A2 net94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1710_ _0538_ _0596_ vssd1 vssd1 vccd1 vccd1 _0626_ sky130_fd_sc_hd__or2_2
X_2690_ gamelogic.letter\[2\] gamelogic.setWord\[26\] vssd1 vssd1 vccd1 vccd1 _1255_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_41_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1641_ _0543_ _0552_ _0368_ vssd1 vssd1 vccd1 vccd1 _0576_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_6_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3292__CLK clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1572_ dispFSM.msg\[4\] _0519_ _0455_ vssd1 vssd1 vccd1 vccd1 _0520_ sky130_fd_sc_hd__o21a_1
XFILLER_0_123_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3311_ clknet_leaf_35_clk uart_receiver.next_clk_count\[3\] net159 vssd1 vssd1 vccd1
+ vccd1 uart_receiver.clk_count\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_191_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3242_ clknet_leaf_5_clk hostdisp.nextBottom\[40\] net199 vssd1 vssd1 vccd1 vccd1
+ hostdisp.bottom\[40\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_89 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3173_ clknet_leaf_14_clk _0149_ net202 vssd1 vssd1 vccd1 vccd1 hostdisp.top\[57\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_175_Right_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2124_ hostdisp.curr_guesses\[4\] net120 _0864_ net133 vssd1 vssd1 vccd1 vccd1 hostdisp.nextBottom\[44\]
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_107_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2428__B _0827_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2055_ hostdisp.curr_word\[3\] net98 _0835_ net143 vssd1 vssd1 vccd1 vccd1 hostdisp.next_curr_word\[3\]
+ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_101_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2025__A2 net95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2957_ host_message_reg.setLetter\[4\] net52 net48 gamelogic.setWord\[4\] vssd1 vssd1
+ vccd1 vccd1 _0320_ sky130_fd_sc_hd__o22a_1
XFILLER_0_32_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2888_ dispFSM.guesses\[28\] net85 net60 net554 vssd1 vssd1 vccd1 vccd1 _0255_ sky130_fd_sc_hd__o22a_1
XFILLER_0_96_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1908_ lcdPlayer.cnt_500hz\[8\] lcdPlayer.cnt_500hz\[12\] lcdPlayer.cnt_500hz\[14\]
+ lcdPlayer.cnt_500hz\[9\] vssd1 vssd1 vccd1 vccd1 _0761_ sky130_fd_sc_hd__or4bb_1
X_1839_ clock_div.count\[18\] _0717_ net402 vssd1 vssd1 vccd1 vccd1 _0718_ sky130_fd_sc_hd__a21oi_1
XANTENNA__2981__B1 net48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout105_X net105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3509_ clknet_leaf_29_clk hostdisp.next_curr_word\[31\] net181 vssd1 vssd1 vccd1
+ vccd1 hostdisp.curr_word\[31\] sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_142_Right_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_169_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3165__CLK clknet_leaf_30_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2016__A2 net94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_259 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_298 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2724__B1 _1286_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput40 net40 vssd1 vssd1 vccd1 vccd1 gpio_out[30] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_91_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3508__CLK clknet_leaf_31_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_28_clk clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_28_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_187_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_175_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_34_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_160_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_183_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2007__A2 net95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_32_clk_A clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2811_ _0364_ _0916_ _1286_ _1275_ _0926_ vssd1 vssd1 vccd1 vccd1 _1357_ sky130_fd_sc_hd__o32a_1
X_2742_ keypadFSMHost.state\[2\] keypadFSMHost.state\[3\] _0613_ _1295_ vssd1 vssd1
+ vccd1 vccd1 _1296_ sky130_fd_sc_hd__or4_1
XFILLER_0_143_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_139_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3510__SET_B net164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2673_ _0381_ gamelogic.letter\[4\] gamelogic.setWord\[37\] _0384_ vssd1 vssd1 vccd1
+ vccd1 _1239_ sky130_fd_sc_hd__a22o_1
X_1624_ keypadHostt.scan_col\[0\] net153 net151 vssd1 vssd1 vccd1 vccd1 _0559_ sky130_fd_sc_hd__or3_2
XFILLER_0_169_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1555_ _0471_ _0490_ _0495_ vssd1 vssd1 vccd1 vccd1 _0503_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_99_Right_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3225_ clknet_leaf_11_clk _0199_ net216 vssd1 vssd1 vccd1 vccd1 keypadFSMHost.prev_key\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_1486_ _0415_ net154 keypadplayer.scan_col\[0\] vssd1 vssd1 vccd1 vccd1 _0438_ sky130_fd_sc_hd__a21o_1
XFILLER_0_94_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3156_ clknet_leaf_31_clk _0132_ net163 vssd1 vssd1 vccd1 vccd1 hostdisp.top\[40\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__3188__CLK clknet_leaf_31_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3087_ clknet_leaf_19_clk _0077_ net211 vssd1 vssd1 vccd1 vccd1 message_reg.msg\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_19_clk clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_19_clk
+ sky130_fd_sc_hd__clkbuf_8
X_2107_ hostdisp.curr_word\[35\] net98 _0855_ net143 vssd1 vssd1 vccd1 vccd1 hostdisp.next_curr_word\[35\]
+ sky130_fd_sc_hd__o22a_1
XANTENNA__3331__Q gamelogic.indexCorrect\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2038_ net142 net92 net77 net545 vssd1 vssd1 vccd1 vccd1 hostdisp.next_curr_guesses\[44\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_11_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_91 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2954__B1 net49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_157_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3332__RESET_B net165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout82_A _0940_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_202 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1428__A net142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3330__CLK clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3010_ net223 vssd1 vssd1 vccd1 vccd1 _0035_ sky130_fd_sc_hd__inv_2
XFILLER_0_64_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3480__CLK clknet_leaf_31_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_143 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_156_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_179 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2725_ keypadFSMHost.unlocked _0546_ _0552_ vssd1 vssd1 vccd1 vccd1 _1287_ sky130_fd_sc_hd__and3_4
XFILLER_0_120_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_8_clk clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_8_clk
+ sky130_fd_sc_hd__clkbuf_8
X_2656_ dispFSM.guesses\[71\] _1072_ _1084_ dispFSM.guesses\[7\] _1226_ vssd1 vssd1
+ vccd1 vccd1 _1227_ sky130_fd_sc_hd__a221o_1
X_1607_ net233 net6 net229 vssd1 vssd1 vccd1 vccd1 _0542_ sky130_fd_sc_hd__o21ba_2
Xfanout104 _0625_ vssd1 vssd1 vccd1 vccd1 net104 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_59_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2587_ net293 net107 _1161_ net183 vssd1 vssd1 vccd1 vccd1 _0177_ sky130_fd_sc_hd__o211a_1
X_1538_ keypadFSMPlayer.prev_key\[7\] _0429_ vssd1 vssd1 vccd1 vccd1 _0486_ sky130_fd_sc_hd__xor2_1
Xfanout137 hostdisp.Cstate vssd1 vssd1 vccd1 vccd1 net137 sky130_fd_sc_hd__buf_2
Xfanout115 _1076_ vssd1 vssd1 vccd1 vccd1 net115 sky130_fd_sc_hd__buf_2
Xfanout126 _0858_ vssd1 vssd1 vccd1 vccd1 net126 sky130_fd_sc_hd__buf_2
Xfanout148 keypadplayer.scan_col\[1\] vssd1 vssd1 vccd1 vccd1 net148 sky130_fd_sc_hd__buf_2
X_1469_ net4 net232 net6 net3 net231 vssd1 vssd1 vccd1 vccd1 _0421_ sky130_fd_sc_hd__o41a_1
Xfanout159 net160 vssd1 vssd1 vccd1 vccd1 net159 sky130_fd_sc_hd__buf_2
X_3208_ clknet_leaf_29_clk _0184_ vssd1 vssd1 vccd1 vccd1 lcdPlayer.currentState\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_3139_ clknet_leaf_26_clk _0115_ vssd1 vssd1 vccd1 vccd1 lcdPlayer.cnt_20ms\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__2467__A2 net73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_107_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_148 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_159_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_80 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3203__CLK clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_162_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3353__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold180 dispFSM.guesses\[63\] vssd1 vssd1 vccd1 vccd1 net444 sky130_fd_sc_hd__dlygate4sd3_1
Xhold191 clock_div.count\[13\] vssd1 vssd1 vccd1 vccd1 net455 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1711__A net2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_49 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_177_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_107 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_141_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3490_ clknet_leaf_30_clk hostdisp.next_curr_word\[12\] net178 vssd1 vssd1 vccd1
+ vccd1 hostdisp.curr_word\[12\] sky130_fd_sc_hd__dfstp_1
XFILLER_0_11_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_13 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2510_ dispFSM.guesses\[8\] _1078_ net112 dispFSM.guesses\[48\] vssd1 vssd1 vccd1
+ vccd1 _1088_ sky130_fd_sc_hd__a22o_1
X_2441_ net340 net67 _1042_ vssd1 vssd1 vccd1 vccd1 _0150_ sky130_fd_sc_hd__o21a_1
XFILLER_0_51_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2372_ net422 _1004_ _1006_ vssd1 vssd1 vccd1 vccd1 _0117_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_75_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_188_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout132_A net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2708_ net143 gamelogic.setWord\[19\] vssd1 vssd1 vccd1 vccd1 _1272_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_154_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2639_ hostdisp.bottom\[70\] net111 _1096_ hostdisp.top\[70\] _1210_ vssd1 vssd1
+ vccd1 vccd1 _1211_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_7_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_165_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_139_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2612__A2 _1081_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_162 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_162_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3249__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_142_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2990_ gamelogic.setWord\[29\] net55 _1394_ gamelogic.setWord\[37\] vssd1 vssd1 vccd1
+ vccd1 _0353_ sky130_fd_sc_hd__a22o_1
XANTENNA__3399__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2603__A2 net106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1941_ _0770_ _0182_ _0786_ vssd1 vssd1 vccd1 vccd1 _0787_ sky130_fd_sc_hd__a21o_1
X_1872_ uart_transmitter.clk_count\[0\] uart_transmitter.clk_count\[1\] uart_transmitter.clk_count\[2\]
+ vssd1 vssd1 vccd1 vccd1 _0734_ sky130_fd_sc_hd__and3_1
XFILLER_0_9_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3611_ net242 vssd1 vssd1 vccd1 vccd1 gpio_out[19] sky130_fd_sc_hd__buf_2
XFILLER_0_126_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3542_ clknet_leaf_6_clk hostdisp.next_curr_guesses\[24\] net196 vssd1 vssd1 vccd1
+ vccd1 hostdisp.curr_guesses\[24\] sky130_fd_sc_hd__dfstp_1
XFILLER_0_101_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3473_ clknet_leaf_0_clk _0351_ net175 vssd1 vssd1 vccd1 vccd1 gamelogic.setWord\[35\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_177_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2424_ hostdisp.curr_word\[9\] _0827_ vssd1 vssd1 vccd1 vccd1 _1035_ sky130_fd_sc_hd__or2_1
X_2355_ lcdPlayer.cnt_20ms\[4\] _0945_ vssd1 vssd1 vccd1 vccd1 _0996_ sky130_fd_sc_hd__or2_1
XFILLER_0_86_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_4_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2286_ net167 _0948_ _0954_ vssd1 vssd1 vccd1 vccd1 _0955_ sky130_fd_sc_hd__and3_2
XFILLER_0_126_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_104_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_230 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_115_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_189_Right_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_86_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3541__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout48_X net48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_174_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_156_Right_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_47 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2140_ gamelogic.setWord\[4\] _0872_ net132 vssd1 vssd1 vccd1 vccd1 hostdisp.nextBottom\[52\]
+ sky130_fd_sc_hd__mux2_1
X_2071_ hostdisp.curr_word\[14\] net102 _0840_ gamelogic.letter\[6\] vssd1 vssd1 vccd1
+ vccd1 hostdisp.next_curr_word\[14\] sky130_fd_sc_hd__o22a_1
XFILLER_0_163_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_17_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2973_ gamelogic.setWord\[12\] net51 net47 gamelogic.setWord\[20\] vssd1 vssd1 vccd1
+ vccd1 _0336_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_60_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1924_ lcdPlayer.currentState\[3\] net106 vssd1 vssd1 vccd1 vccd1 _0774_ sky130_fd_sc_hd__or2_1
XFILLER_0_173_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1855_ _0726_ _0727_ vssd1 vssd1 vccd1 vccd1 clock_div.next_count\[25\] sky130_fd_sc_hd__nor2_1
XFILLER_0_112_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1786_ clock_div.count\[19\] clock_div.count\[18\] clock_div.count\[21\] clock_div.count\[20\]
+ vssd1 vssd1 vccd1 vccd1 _0684_ sky130_fd_sc_hd__or4_1
X_3525_ clknet_leaf_14_clk net346 net206 vssd1 vssd1 vccd1 vccd1 hostdisp.curr_guesses\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkload34_A clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_151_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_123_Right_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3414__CLK clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3456_ clknet_leaf_2_clk _0334_ net175 vssd1 vssd1 vccd1 vccd1 gamelogic.setWord\[18\]
+ sky130_fd_sc_hd__dfstp_1
X_2407_ _1028_ net304 _0934_ vssd1 vssd1 vccd1 vccd1 _0130_ sky130_fd_sc_hd__mux2_1
X_3387_ clknet_leaf_21_clk _0276_ net210 vssd1 vssd1 vccd1 vccd1 dispFSM.guesses\[41\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_41_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3564__CLK clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2338_ lcdPlayer.cnt_500hz\[19\] lcdPlayer.cnt_500hz\[18\] _0984_ vssd1 vssd1 vccd1
+ vccd1 _0988_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_179_Left_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2269_ dispFSM.msg\[3\] _0941_ _0942_ net351 vssd1 vssd1 vccd1 vccd1 _0078_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_162_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_344 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2579__A1 dispFSM.msg\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_188_Left_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold40 keypadplayer.scan_col\[2\] vssd1 vssd1 vccd1 vccd1 net304 sky130_fd_sc_hd__dlygate4sd3_1
Xhold51 dispFSM.guesses\[7\] vssd1 vssd1 vccd1 vccd1 net315 sky130_fd_sc_hd__dlygate4sd3_1
Xhold62 buffer.Rx_byte\[1\] vssd1 vssd1 vccd1 vccd1 net326 sky130_fd_sc_hd__dlygate4sd3_1
Xhold73 hostdisp.top\[50\] vssd1 vssd1 vccd1 vccd1 net337 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_187_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold95 clock_div.count\[18\] vssd1 vssd1 vccd1 vccd1 net359 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold84 _0147_ vssd1 vssd1 vccd1 vccd1 net348 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_187_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2806__A2 _0394_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_196 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1640_ _0367_ _0544_ _0552_ vssd1 vssd1 vccd1 vccd1 _0575_ sky130_fd_sc_hd__and3_1
XANTENNA__2990__B2 gamelogic.setWord\[37\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2990__A1 gamelogic.setWord\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1571_ _0372_ keypadFSMPlayer.state\[0\] _0442_ _0453_ vssd1 vssd1 vccd1 vccd1 _0519_
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_158_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3310_ clknet_leaf_34_clk uart_receiver.next_clk_count\[2\] net159 vssd1 vssd1 vccd1
+ vccd1 uart_receiver.clk_count\[2\] sky130_fd_sc_hd__dfrtp_1
X_3241_ clknet_leaf_10_clk keypadFSMHost.next_state\[2\] net215 vssd1 vssd1 vccd1
+ vccd1 _1398_ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_184_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3172_ clknet_leaf_22_clk _0148_ net185 vssd1 vssd1 vccd1 vccd1 hostdisp.top\[56\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_6_clk_A clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2123_ gamelogic.setWord\[4\] net123 vssd1 vssd1 vccd1 vccd1 _0864_ sky130_fd_sc_hd__or2_1
XFILLER_0_83_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2054_ hostdisp.curr_word\[2\] net98 _0835_ gamelogic.letter\[2\] vssd1 vssd1 vccd1
+ vccd1 hostdisp.next_curr_word\[2\] sky130_fd_sc_hd__o22a_1
XFILLER_0_88_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2956_ host_message_reg.setLetter\[3\] net52 net48 gamelogic.setWord\[3\] vssd1 vssd1
+ vccd1 vccd1 _0319_ sky130_fd_sc_hd__o22a_1
XFILLER_0_91_339 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2430__B1 net70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2887_ dispFSM.guesses\[27\] net82 net57 net522 vssd1 vssd1 vccd1 vccd1 _0254_ sky130_fd_sc_hd__o22a_1
X_1907_ net139 net106 vssd1 vssd1 vccd1 vccd1 _0760_ sky130_fd_sc_hd__nand2_1
X_1838_ net359 _0717_ vssd1 vssd1 vccd1 vccd1 clock_div.next_count\[18\] sky130_fd_sc_hd__xor2_1
XANTENNA_fanout212_A net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2733__A1 net6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1769_ _0397_ uart_transmitter.state\[0\] _0399_ vssd1 vssd1 vccd1 vccd1 _0670_ sky130_fd_sc_hd__and3_1
XFILLER_0_12_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3508_ clknet_leaf_31_clk hostdisp.next_curr_word\[30\] net173 vssd1 vssd1 vccd1
+ vccd1 hostdisp.curr_word\[30\] sky130_fd_sc_hd__dfstp_1
X_3439_ clknet_leaf_13_clk _0317_ net197 vssd1 vssd1 vccd1 vccd1 gamelogic.setWord\[1\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_0_169_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3120__RESET_B net223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2421__B1 net69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_130_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput41 net41 vssd1 vssd1 vccd1 vccd1 gpio_out[31] sky130_fd_sc_hd__buf_2
Xoutput30 net30 vssd1 vssd1 vccd1 vccd1 gpio_out[11] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_91_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_160_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2810_ gamelogic.state\[0\] _0916_ _1355_ _1260_ vssd1 vssd1 vccd1 vccd1 _1356_ sky130_fd_sc_hd__o31a_1
XFILLER_0_183_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2741_ _1398_ _1294_ keypadFSMHost.state\[5\] vssd1 vssd1 vccd1 vccd1 _1295_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_26_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_42_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_139_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1608__B net4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2672_ gamelogic.setWord\[33\] net144 vssd1 vssd1 vccd1 vccd1 _1238_ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1623_ _0557_ vssd1 vssd1 vccd1 vccd1 _0558_ sky130_fd_sc_hd__inv_2
XFILLER_0_151_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1554_ _0500_ _0501_ _0428_ vssd1 vssd1 vccd1 vccd1 _0502_ sky130_fd_sc_hd__a21oi_1
X_1485_ _0422_ _0436_ vssd1 vssd1 vccd1 vccd1 _0437_ sky130_fd_sc_hd__nor2_1
XFILLER_0_185_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3224_ clknet_leaf_16_clk _0198_ net223 vssd1 vssd1 vccd1 vccd1 keypadFSMHost.prev_key\[1\]
+ sky130_fd_sc_hd__dfrtp_1
.ends

