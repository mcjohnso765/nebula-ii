* NGSPICE file created from team_04.ext - technology: sky130A

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41ai_2 abstract view
.subckt sky130_fd_sc_hd__o41ai_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_2 abstract view
.subckt sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_4 abstract view
.subckt sky130_fd_sc_hd__o32a_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_2 abstract view
.subckt sky130_fd_sc_hd__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_4 abstract view
.subckt sky130_fd_sc_hd__a32oi_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_1 abstract view
.subckt sky130_fd_sc_hd__a311oi_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_4 abstract view
.subckt sky130_fd_sc_hd__a32o_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_4 abstract view
.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_4 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_16 abstract view
.subckt sky130_fd_sc_hd__clkinv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinvlp_4 abstract view
.subckt sky130_fd_sc_hd__clkinvlp_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_4 abstract view
.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__bufinv_16 abstract view
.subckt sky130_fd_sc_hd__bufinv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_16 abstract view
.subckt sky130_fd_sc_hd__inv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_8 abstract view
.subckt sky130_fd_sc_hd__clkinv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_8 abstract view
.subckt sky130_fd_sc_hd__inv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_12 abstract view
.subckt sky130_fd_sc_hd__inv_12 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_2 abstract view
.subckt sky130_fd_sc_hd__o221ai_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_4 abstract view
.subckt sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311ai_1 abstract view
.subckt sky130_fd_sc_hd__o311ai_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_1 abstract view
.subckt sky130_fd_sc_hd__o2111ai_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_4 abstract view
.subckt sky130_fd_sc_hd__a22o_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_4 abstract view
.subckt sky130_fd_sc_hd__a41o_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_4 abstract view
.subckt sky130_fd_sc_hd__o41a_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_4 abstract view
.subckt sky130_fd_sc_hd__a221o_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_4 abstract view
.subckt sky130_fd_sc_hd__and3b_4 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_2 abstract view
.subckt sky130_fd_sc_hd__o2111ai_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_2 abstract view
.subckt sky130_fd_sc_hd__a32oi_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

.subckt team_04 ACK_I ADR_O[0] ADR_O[10] ADR_O[11] ADR_O[12] ADR_O[13] ADR_O[14] ADR_O[15]
+ ADR_O[16] ADR_O[17] ADR_O[18] ADR_O[19] ADR_O[1] ADR_O[20] ADR_O[21] ADR_O[22] ADR_O[23]
+ ADR_O[24] ADR_O[25] ADR_O[26] ADR_O[27] ADR_O[28] ADR_O[29] ADR_O[2] ADR_O[30] ADR_O[31]
+ ADR_O[3] ADR_O[4] ADR_O[5] ADR_O[6] ADR_O[7] ADR_O[8] ADR_O[9] CYC_O DAT_I[0] DAT_I[10]
+ DAT_I[11] DAT_I[12] DAT_I[13] DAT_I[14] DAT_I[15] DAT_I[16] DAT_I[17] DAT_I[18]
+ DAT_I[19] DAT_I[1] DAT_I[20] DAT_I[21] DAT_I[22] DAT_I[23] DAT_I[24] DAT_I[25] DAT_I[26]
+ DAT_I[27] DAT_I[28] DAT_I[29] DAT_I[2] DAT_I[30] DAT_I[31] DAT_I[3] DAT_I[4] DAT_I[5]
+ DAT_I[6] DAT_I[7] DAT_I[8] DAT_I[9] DAT_O[0] DAT_O[10] DAT_O[11] DAT_O[12] DAT_O[13]
+ DAT_O[14] DAT_O[15] DAT_O[16] DAT_O[17] DAT_O[18] DAT_O[19] DAT_O[1] DAT_O[20] DAT_O[21]
+ DAT_O[22] DAT_O[23] DAT_O[24] DAT_O[25] DAT_O[26] DAT_O[27] DAT_O[28] DAT_O[29]
+ DAT_O[2] DAT_O[30] DAT_O[31] DAT_O[3] DAT_O[4] DAT_O[5] DAT_O[6] DAT_O[7] DAT_O[8]
+ DAT_O[9] SEL_O[0] SEL_O[1] SEL_O[2] SEL_O[3] STB_O WE_O clk en gpio_in[0] gpio_in[10]
+ gpio_in[11] gpio_in[12] gpio_in[13] gpio_in[14] gpio_in[15] gpio_in[16] gpio_in[17]
+ gpio_in[18] gpio_in[19] gpio_in[1] gpio_in[20] gpio_in[21] gpio_in[22] gpio_in[23]
+ gpio_in[24] gpio_in[25] gpio_in[26] gpio_in[27] gpio_in[28] gpio_in[29] gpio_in[2]
+ gpio_in[30] gpio_in[31] gpio_in[32] gpio_in[33] gpio_in[3] gpio_in[4] gpio_in[5]
+ gpio_in[6] gpio_in[7] gpio_in[8] gpio_in[9] gpio_oeb[0] gpio_oeb[10] gpio_oeb[11]
+ gpio_oeb[12] gpio_oeb[13] gpio_oeb[14] gpio_oeb[15] gpio_oeb[16] gpio_oeb[17] gpio_oeb[18]
+ gpio_oeb[19] gpio_oeb[1] gpio_oeb[20] gpio_oeb[21] gpio_oeb[22] gpio_oeb[23] gpio_oeb[24]
+ gpio_oeb[25] gpio_oeb[26] gpio_oeb[27] gpio_oeb[28] gpio_oeb[29] gpio_oeb[2] gpio_oeb[30]
+ gpio_oeb[31] gpio_oeb[32] gpio_oeb[33] gpio_oeb[3] gpio_oeb[4] gpio_oeb[5] gpio_oeb[6]
+ gpio_oeb[7] gpio_oeb[8] gpio_oeb[9] gpio_out[0] gpio_out[10] gpio_out[11] gpio_out[12]
+ gpio_out[13] gpio_out[14] gpio_out[15] gpio_out[16] gpio_out[17] gpio_out[18] gpio_out[19]
+ gpio_out[1] gpio_out[20] gpio_out[21] gpio_out[22] gpio_out[23] gpio_out[24] gpio_out[25]
+ gpio_out[26] gpio_out[27] gpio_out[28] gpio_out[29] gpio_out[2] gpio_out[30] gpio_out[31]
+ gpio_out[32] gpio_out[33] gpio_out[3] gpio_out[4] gpio_out[5] gpio_out[6] gpio_out[7]
+ gpio_out[8] gpio_out[9] mem_adr_start[0] mem_adr_start[10] mem_adr_start[11] mem_adr_start[12]
+ mem_adr_start[13] mem_adr_start[14] mem_adr_start[15] mem_adr_start[16] mem_adr_start[17]
+ mem_adr_start[18] mem_adr_start[19] mem_adr_start[1] mem_adr_start[20] mem_adr_start[21]
+ mem_adr_start[22] mem_adr_start[23] mem_adr_start[24] mem_adr_start[25] mem_adr_start[26]
+ mem_adr_start[27] mem_adr_start[28] mem_adr_start[29] mem_adr_start[2] mem_adr_start[30]
+ mem_adr_start[31] mem_adr_start[3] mem_adr_start[4] mem_adr_start[5] mem_adr_start[6]
+ mem_adr_start[7] mem_adr_start[8] mem_adr_start[9] memory_size[0] memory_size[10]
+ memory_size[11] memory_size[12] memory_size[13] memory_size[14] memory_size[15]
+ memory_size[16] memory_size[17] memory_size[18] memory_size[19] memory_size[1] memory_size[20]
+ memory_size[21] memory_size[22] memory_size[23] memory_size[24] memory_size[25]
+ memory_size[26] memory_size[27] memory_size[28] memory_size[29] memory_size[2] memory_size[30]
+ memory_size[31] memory_size[3] memory_size[4] memory_size[5] memory_size[6] memory_size[7]
+ memory_size[8] memory_size[9] nrst vccd1 vssd1
XFILLER_0_78_1821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06883_ final_design.cpu.reg_window\[211\] final_design.cpu.reg_window\[243\] net911
+ vssd1 vssd1 vccd1 vccd1 _01834_ sky130_fd_sc_hd__mux2_1
X_09671_ net261 _04582_ _04587_ _04589_ vssd1 vssd1 vccd1 vccd1 _04590_ sky130_fd_sc_hd__and4_1
XFILLER_0_74_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10023__B _04940_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11834__S net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08622_ net597 _03257_ _03232_ _02156_ vssd1 vssd1 vccd1 vccd1 _03573_ sky130_fd_sc_hd__o211a_1
XFILLER_0_27_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06928__S net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13840__CLK clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11618__B1 net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08553_ final_design.cpu.reg_window\[897\] final_design.cpu.reg_window\[929\] net833
+ vssd1 vssd1 vccd1 vccd1 _03504_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07504_ _02002_ _02032_ _02449_ _02454_ _02453_ vssd1 vssd1 vccd1 vccd1 _02455_ sky130_fd_sc_hd__o41ai_2
XANTENNA__12291__B1 net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08484_ final_design.cpu.reg_window\[131\] final_design.cpu.reg_window\[163\] net824
+ vssd1 vssd1 vccd1 vccd1 _03435_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_2350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_2361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_2372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07435_ final_design.cpu.reg_window\[513\] final_design.cpu.reg_window\[545\] net912
+ vssd1 vssd1 vccd1 vccd1 _02386_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10396__D _05174_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13990__CLK clknet_leaf_51_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10841__B2 net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout427_A net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07759__S net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1169_A net1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07366_ _02313_ _02314_ _02315_ _02316_ net767 net787 vssd1 vssd1 vccd1 vccd1 _02317_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__06663__S net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07288__A1_N net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09105_ _04026_ _01367_ net254 vssd1 vssd1 vccd1 vccd1 _04027_ sky130_fd_sc_hd__mux2_1
XANTENNA__12594__B2 final_design.data_from_mem\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07297_ net760 _02247_ vssd1 vssd1 vccd1 vccd1 _02248_ sky130_fd_sc_hd__or2_1
XANTENNA__13220__CLK clknet_leaf_54_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout215_X net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1246 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09036_ final_design.CPU_instr_adr\[11\] _03966_ net1037 vssd1 vssd1 vccd1 vccd1
+ _00222_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_57_2143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_2154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout796_A _06333_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_2788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_2165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_2799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_2007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold340 final_design.cpu.reg_window\[737\] vssd1 vssd1 vccd1 vccd1 net1682 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_53_2018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10357__B1 net1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold351 final_design.cpu.reg_window\[878\] vssd1 vssd1 vccd1 vccd1 net1693 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_53_2029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold362 final_design.cpu.reg_window\[455\] vssd1 vssd1 vccd1 vccd1 net1704 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold373 final_design.cpu.reg_window\[140\] vssd1 vssd1 vccd1 vccd1 net1715 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_51_clk_X clknet_leaf_51_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold384 final_design.cpu.reg_window\[452\] vssd1 vssd1 vccd1 vccd1 net1726 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13370__CLK clknet_leaf_58_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout963_A _04036_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold395 final_design.cpu.reg_window\[976\] vssd1 vssd1 vccd1 vccd1 net1737 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout820 net824 vssd1 vssd1 vccd1 vccd1 net820 sky130_fd_sc_hd__clkbuf_4
Xfanout831 net834 vssd1 vssd1 vccd1 vccd1 net831 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12938__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09938_ _04222_ _04581_ _04586_ _04727_ _04856_ vssd1 vssd1 vccd1 vccd1 _04857_ sky130_fd_sc_hd__o221a_1
Xfanout842 _01818_ vssd1 vssd1 vccd1 vccd1 net842 sky130_fd_sc_hd__buf_2
Xfanout853 net854 vssd1 vssd1 vccd1 vccd1 net853 sky130_fd_sc_hd__clkbuf_4
Xfanout864 net865 vssd1 vssd1 vccd1 vccd1 net864 sky130_fd_sc_hd__clkbuf_4
Xfanout875 net876 vssd1 vssd1 vccd1 vccd1 net875 sky130_fd_sc_hd__buf_4
XANTENNA__09514__A2 net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout886 _01437_ vssd1 vssd1 vccd1 vccd1 net886 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_57_1905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09869_ _04770_ _04787_ vssd1 vssd1 vccd1 vccd1 _04788_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_5_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout897 net898 vssd1 vssd1 vccd1 vccd1 net897 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout751_X net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1040 final_design.cpu.reg_window\[98\] vssd1 vssd1 vccd1 vccd1 net2382 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11744__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1051 final_design.cpu.reg_window\[635\] vssd1 vssd1 vccd1 vccd1 net2393 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1062 final_design.cpu.reg_window\[621\] vssd1 vssd1 vccd1 vccd1 net2404 sky130_fd_sc_hd__dlygate4sd3_1
X_11900_ net206 net1952 net272 vssd1 vssd1 vccd1 vccd1 _00642_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_1375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12880_ clknet_leaf_18_clk _00118_ net1111 vssd1 vssd1 vccd1 vccd1 final_design.data_from_mem\[14\]
+ sky130_fd_sc_hd__dfrtp_4
Xhold1073 final_design.cpu.reg_window\[291\] vssd1 vssd1 vccd1 vccd1 net2415 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1084 final_design.cpu.reg_window\[668\] vssd1 vssd1 vccd1 vccd1 net2426 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08619__A net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1095 final_design.cpu.reg_window\[701\] vssd1 vssd1 vccd1 vccd1 net2437 sky130_fd_sc_hd__dlygate4sd3_1
X_11831_ net197 net2219 net266 vssd1 vssd1 vccd1 vccd1 _00583_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12282__B1 net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11762_ net186 net2082 net419 vssd1 vssd1 vccd1 vccd1 _00525_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13501_ clknet_leaf_2_clk _00732_ net1077 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[489\]
+ sky130_fd_sc_hd__dfrtp_1
X_10713_ final_design.CPU_instr_adr\[13\] _05451_ net1053 vssd1 vssd1 vccd1 vccd1
+ _05452_ sky130_fd_sc_hd__mux2_1
XANTENNA__10832__B2 net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11693_ net214 net627 vssd1 vssd1 vccd1 vccd1 _06205_ sky130_fd_sc_hd__and2_1
XFILLER_0_3_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input92_A memory_size[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13432_ clknet_leaf_64_clk _00663_ net1075 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[420\]
+ sky130_fd_sc_hd__dfrtp_1
X_10644_ _05347_ _05385_ _05386_ vssd1 vssd1 vccd1 vccd1 _05387_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11699__B net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06573__S net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12872__Q final_design.data_from_mem\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11388__A2 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12585__B2 final_design.data_from_mem\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10575_ final_design.CPU_instr_adr\[6\] _04002_ net1057 vssd1 vssd1 vccd1 vccd1 _05321_
+ sky130_fd_sc_hd__mux2_1
X_13363_ clknet_leaf_40_clk _00594_ net1211 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[351\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09169__B net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12314_ net1809 net203 net366 vssd1 vssd1 vccd1 vccd1 _01028_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_20_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13294_ clknet_leaf_43_clk _00525_ net1223 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[282\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13713__CLK clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12245_ net558 _06175_ net502 net372 net1485 vssd1 vssd1 vccd1 vccd1 _00962_ sky130_fd_sc_hd__a32o_1
XANTENNA__12163__X _06270_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_19_clk_X clknet_leaf_19_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12176_ net2432 net212 net380 vssd1 vssd1 vccd1 vccd1 _00895_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08961__B1 net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11127_ _01487_ net653 net1013 vssd1 vssd1 vccd1 vccd1 _05842_ sky130_fd_sc_hd__a21o_1
XANTENNA__13863__CLK clknet_leaf_59_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11058_ net89 net1047 vssd1 vssd1 vccd1 vccd1 _05781_ sky130_fd_sc_hd__and2_1
XANTENNA__11848__B1 net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10009_ _04085_ _04685_ _04927_ vssd1 vssd1 vccd1 vccd1 _04928_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_8_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_1773 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12273__B1 net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13243__CLK clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07220_ net749 _02164_ net745 vssd1 vssd1 vccd1 vccd1 _02171_ sky130_fd_sc_hd__o21a_1
XFILLER_0_73_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07151_ final_design.cpu.reg_window\[458\] final_design.cpu.reg_window\[490\] net899
+ vssd1 vssd1 vccd1 vccd1 _02102_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_1544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08244__A2 _03192_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_191 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07082_ _02026_ _02031_ vssd1 vssd1 vccd1 vccd1 _02033_ sky130_fd_sc_hd__or2_1
XANTENNA__13393__CLK clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11829__S net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1733 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08711__B _01630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_2630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_2641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09744__A2 net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1777 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11551__A2 net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07984_ _02932_ _02933_ vssd1 vssd1 vccd1 vccd1 _02935_ sky130_fd_sc_hd__nor2_1
X_09723_ net548 net546 net545 net544 net454 net464 vssd1 vssd1 vccd1 vccd1 _04642_
+ sky130_fd_sc_hd__mux4_1
X_06935_ final_design.cpu.reg_window\[401\] final_design.cpu.reg_window\[433\] net928
+ vssd1 vssd1 vccd1 vccd1 _01886_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout377_A _06271_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09654_ _04189_ _04572_ vssd1 vssd1 vccd1 vccd1 _04573_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_1526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06866_ _01393_ net993 net990 _01380_ vssd1 vssd1 vccd1 vccd1 _01817_ sky130_fd_sc_hd__a31o_2
XTAP_TAPCELL_ROW_69_2570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_2412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_2423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_2434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08605_ _02390_ net460 vssd1 vssd1 vccd1 vccd1 _03556_ sky130_fd_sc_hd__nand2_1
X_06797_ _01744_ _01745_ _01746_ _01747_ net770 net789 vssd1 vssd1 vccd1 vccd1 _01748_
+ sky130_fd_sc_hd__mux4_1
X_09585_ _03199_ _03229_ _04503_ _04140_ vssd1 vssd1 vccd1 vccd1 _04504_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout544_A _01937_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11067__A1 net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12264__A0 net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08536_ net595 _03481_ _03483_ _02356_ vssd1 vssd1 vccd1 vccd1 _03487_ sky130_fd_sc_hd__o211a_1
XFILLER_0_72_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07366__S0 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1879 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout711_A net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12395__S net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08467_ net609 _03415_ _03416_ vssd1 vssd1 vccd1 vccd1 _03418_ sky130_fd_sc_hd__a21oi_2
XANTENNA_fanout332_X net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout809_A net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12016__B1 net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07418_ _02365_ _02366_ _02367_ _02368_ net770 net789 vssd1 vssd1 vccd1 vccd1 _02369_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_64_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08398_ final_design.cpu.reg_window\[518\] final_design.cpu.reg_window\[550\] net823
+ vssd1 vssd1 vccd1 vccd1 _03349_ sky130_fd_sc_hd__mux2_1
XANTENNA__13736__CLK clknet_leaf_40_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_2216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07349_ _02298_ _02299_ vssd1 vssd1 vccd1 vccd1 _02300_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_59_2227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_2238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14200__1258 vssd1 vssd1 vccd1 vccd1 _14200__1258/HI net1258 sky130_fd_sc_hd__conb_1
XFILLER_0_66_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10360_ net33 net1024 net1006 final_design.data_from_mem\[9\] vssd1 vssd1 vccd1 vccd1
+ _00113_ sky130_fd_sc_hd__o22a_1
XANTENNA__12319__A1 net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11739__S net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09019_ net255 _03950_ net1013 vssd1 vssd1 vccd1 vccd1 _03952_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11790__A2 net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10291_ final_design.VGA_data_control.data_to_VGA\[23\] final_design.VGA_data_control.data_to_VGA\[22\]
+ final_design.VGA_data_control.data_to_VGA\[21\] final_design.VGA_data_control.data_to_VGA\[20\]
+ net1050 net1049 vssd1 vssd1 vccd1 vccd1 _05145_ sky130_fd_sc_hd__mux4_1
XANTENNA__13886__CLK clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12030_ net1817 net226 net396 vssd1 vssd1 vccd1 vccd1 _00758_ sky130_fd_sc_hd__mux2_1
Xhold170 final_design.VGA_data_control.ready_data\[3\] vssd1 vssd1 vccd1 vccd1 net1512
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold181 final_design.reqhand.instruction\[6\] vssd1 vssd1 vccd1 vccd1 net1523 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06422__A final_design.data_from_mem\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout966_X net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold192 final_design.VGA_data_control.ready_data\[29\] vssd1 vssd1 vccd1 vccd1 net1534
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_18_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_31_clk_A clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout650 _05849_ vssd1 vssd1 vccd1 vccd1 net650 sky130_fd_sc_hd__buf_4
XANTENNA__13116__CLK clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout661 _02512_ vssd1 vssd1 vccd1 vccd1 net661 sky130_fd_sc_hd__clkbuf_2
Xfanout672 _02329_ vssd1 vssd1 vccd1 vccd1 net672 sky130_fd_sc_hd__buf_2
X_13981_ clknet_leaf_1_clk _01212_ net1077 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[969\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout683 net689 vssd1 vssd1 vccd1 vccd1 net683 sky130_fd_sc_hd__buf_4
Xfanout694 net695 vssd1 vssd1 vccd1 vccd1 net694 sky130_fd_sc_hd__buf_4
XANTENNA__11474__S net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12932_ clknet_leaf_31_clk _00170_ net1233 vssd1 vssd1 vccd1 vccd1 net155 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_77_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12867__Q final_design.data_from_mem\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12863_ clknet_leaf_18_clk _00101_ net1114 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.ready_data\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_1178 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1913 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_46_clk_A clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13266__CLK clknet_leaf_39_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11814_ net227 net2289 net265 vssd1 vssd1 vccd1 vccd1 _00566_ sky130_fd_sc_hd__mux2_1
XANTENNA__12255__B1 net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11745_ net219 net2238 net416 vssd1 vssd1 vccd1 vccd1 _00508_ sky130_fd_sc_hd__mux2_1
XANTENNA__12270__A3 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07399__S net913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1143 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12007__B1 net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11676_ net2424 net295 _06196_ net428 vssd1 vssd1 vccd1 vccd1 _00469_ sky130_fd_sc_hd__a22o_1
X_13415_ clknet_leaf_63_clk _00646_ net1122 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[403\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10627_ _05368_ _05369_ vssd1 vssd1 vccd1 vccd1 _05370_ sky130_fd_sc_hd__nand2_1
XFILLER_0_70_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1717 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13346_ clknet_leaf_10_clk _00577_ net1101 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[334\]
+ sky130_fd_sc_hd__dfrtp_1
X_10558_ _05285_ _05303_ vssd1 vssd1 vccd1 vccd1 _05305_ sky130_fd_sc_hd__nor2_1
XANTENNA__08631__C1 _01996_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11781__A2 net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13277_ clknet_leaf_5_clk _00508_ net1078 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[265\]
+ sky130_fd_sc_hd__dfrtp_1
X_10489_ net1042 final_design.reqhand.current_client\[1\] vssd1 vssd1 vccd1 vccd1
+ _05239_ sky130_fd_sc_hd__nand2_4
XFILLER_0_59_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09726__A2 _01657_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12228_ net580 _06156_ net511 net378 net1852 vssd1 vssd1 vccd1 vccd1 _00946_ sky130_fd_sc_hd__a32o_1
XANTENNA__09282__S0 net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09346__C _04086_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_24 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12159_ net180 net2465 net386 vssd1 vssd1 vccd1 vccd1 _00880_ sky130_fd_sc_hd__mux2_1
XANTENNA__07832__S1 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14041__CLK clknet_leaf_15_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10789__A _05508_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12089__A3 net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11237__X _05941_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11297__A1 final_design.data_from_mem\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06720_ final_design.cpu.reg_window\[472\] final_design.cpu.reg_window\[504\] net944
+ vssd1 vssd1 vccd1 vccd1 _01671_ sky130_fd_sc_hd__mux2_1
XANTENNA__13609__CLK clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06478__S net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12494__B1 net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06651_ final_design.cpu.reg_window\[346\] final_design.cpu.reg_window\[378\] net943
+ vssd1 vssd1 vccd1 vccd1 _01602_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_1109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09370_ _04286_ _04288_ vssd1 vssd1 vccd1 vccd1 _04289_ sky130_fd_sc_hd__nand2_1
X_06582_ _01529_ _01530_ _01531_ _01532_ net777 net783 vssd1 vssd1 vccd1 vccd1 _01533_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__13759__CLK clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08321_ final_design.cpu.reg_window\[136\] final_design.cpu.reg_window\[168\] net812
+ vssd1 vssd1 vccd1 vccd1 _03272_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12261__A3 net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08706__B _01507_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1817 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08252_ final_design.cpu.reg_window\[458\] final_design.cpu.reg_window\[490\] net818
+ vssd1 vssd1 vccd1 vccd1 _03203_ sky130_fd_sc_hd__mux2_1
XANTENNA__06476__A1 final_design.data_from_mem\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07203_ net757 _02153_ vssd1 vssd1 vccd1 vccd1 _02154_ sky130_fd_sc_hd__or2_1
XANTENNA__06957__A1_N net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08183_ _03132_ _03133_ vssd1 vssd1 vccd1 vccd1 _03134_ sky130_fd_sc_hd__nor2_2
X_07134_ final_design.cpu.reg_window\[715\] final_design.cpu.reg_window\[747\] net915
+ vssd1 vssd1 vccd1 vccd1 _02085_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_1817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_77_2850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07425__B1 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10024__A2 net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08622__C1 _02156_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_2703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07065_ final_design.cpu.reg_window\[525\] final_design.cpu.reg_window\[557\] net935
+ vssd1 vssd1 vccd1 vccd1 _02016_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1034_A net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13139__CLK clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout494_A net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1201_A net1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07772__S net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout661_A _02512_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07967_ final_design.cpu.reg_window\[977\] final_design.cpu.reg_window\[1009\] net848
+ vssd1 vssd1 vccd1 vccd1 _02918_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout282_X net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout759_A net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_2507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13289__CLK clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09706_ _03101_ _04497_ vssd1 vssd1 vccd1 vccd1 _04625_ sky130_fd_sc_hd__xnor2_1
X_06918_ final_design.cpu.reg_window\[850\] final_design.cpu.reg_window\[882\] net925
+ vssd1 vssd1 vccd1 vccd1 _01869_ sky130_fd_sc_hd__mux2_1
XANTENNA__12485__B1 net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08689__C1 _02419_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07898_ _02845_ _02846_ _02847_ _02848_ net683 net702 vssd1 vssd1 vccd1 vccd1 _02849_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__07587__S0 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09637_ net319 _04264_ _04275_ net320 _04555_ vssd1 vssd1 vccd1 vccd1 _04556_ sky130_fd_sc_hd__a221o_1
X_06849_ final_design.cpu.reg_window\[148\] final_design.cpu.reg_window\[180\] net948
+ vssd1 vssd1 vccd1 vccd1 _01800_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout1191_X net1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout926_A net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07900__A1 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12237__B1 net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09568_ _04485_ _04486_ net477 vssd1 vssd1 vccd1 vccd1 _04487_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08519_ final_design.cpu.reg_window\[834\] final_design.cpu.reg_window\[866\] net832
+ vssd1 vssd1 vccd1 vccd1 _03470_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_1616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout714_X net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09499_ _02609_ _04050_ vssd1 vssd1 vccd1 vccd1 _04418_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07113__C1 _01821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12252__A3 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11323__A net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06467__A1 final_design.data_from_mem\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11530_ net1791 net187 net524 vssd1 vssd1 vccd1 vccd1 _00397_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06417__A net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07012__S net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11461_ net220 net2351 net306 vssd1 vssd1 vccd1 vccd1 _00347_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13200_ clknet_leaf_33_clk _00431_ net1231 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[188\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11212__A1 net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10412_ _03321_ _05181_ vssd1 vssd1 vccd1 vccd1 _05189_ sky130_fd_sc_hd__nor2_1
XANTENNA__10015__A2 _04693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14180_ clknet_leaf_22_clk _01354_ net1164 vssd1 vssd1 vccd1 vccd1 final_design.VGA_adr\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_11392_ net733 _03811_ _06076_ vssd1 vssd1 vccd1 vccd1 _06077_ sky130_fd_sc_hd__o21a_1
XFILLER_0_61_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11469__S net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_695 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13131_ clknet_leaf_38_clk _00362_ net1191 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[119\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_60_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10343_ net1462 net1011 net989 final_design.data_from_mem\[28\] vssd1 vssd1 vccd1
+ vccd1 _00100_ sky130_fd_sc_hd__a22o_1
XFILLER_0_46_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input55_A mem_adr_start[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10274_ final_design.uart.BAUD_counter\[27\] _05133_ net797 vssd1 vssd1 vccd1 vccd1
+ _05135_ sky130_fd_sc_hd__o21ai_1
X_13062_ clknet_leaf_51_clk _00293_ net1169 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[50\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14064__CLK clknet_leaf_15_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11993__A _05869_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1024 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12013_ _06215_ net289 net403 net2374 vssd1 vssd1 vccd1 vccd1 _00744_ sky130_fd_sc_hd__a22o_1
XANTENNA__08401__A1_N net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10723__B1 net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout480 _03484_ vssd1 vssd1 vccd1 vccd1 net480 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_79_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout491 net493 vssd1 vssd1 vccd1 vccd1 net491 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_45_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11279__A1 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10402__A _03481_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13964_ clknet_leaf_46_clk _01195_ net1215 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[952\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09567__S1 net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12476__B1 net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12915_ clknet_leaf_61_clk _00153_ net1137 vssd1 vssd1 vccd1 vccd1 net137 sky130_fd_sc_hd__dfrtp_1
X_13895_ clknet_leaf_59_clk _01126_ net1126 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[883\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13901__CLK clknet_leaf_44_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09892__A1 _02325_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12228__B1 net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12846_ clknet_leaf_17_clk _00084_ net1108 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.ready_data\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_1721 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1131 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09644__A1 _04342_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12243__A3 net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11728_ net435 net586 _06222_ net296 net2402 vssd1 vssd1 vccd1 vccd1 _00495_ sky130_fd_sc_hd__a32o_1
XFILLER_0_16_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11659_ net184 net632 vssd1 vssd1 vccd1 vccd1 _06187_ sky130_fd_sc_hd__and2_1
XFILLER_0_0_1861 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12400__B1 net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold906 final_design.cpu.reg_window\[604\] vssd1 vssd1 vccd1 vccd1 net2248 sky130_fd_sc_hd__dlygate4sd3_1
Xhold917 final_design.uart.working_data\[3\] vssd1 vssd1 vccd1 vccd1 net2259 sky130_fd_sc_hd__dlygate4sd3_1
Xhold928 final_design.cpu.reg_window\[805\] vssd1 vssd1 vccd1 vccd1 net2270 sky130_fd_sc_hd__dlygate4sd3_1
X_13329_ clknet_leaf_35_clk _00560_ net1241 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[317\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09698__A2_N net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold939 final_design.cpu.reg_window\[605\] vssd1 vssd1 vccd1 vccd1 net2281 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1861 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_3_1_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_3_1_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_0_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13431__CLK clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08870_ net625 _03817_ _03818_ net256 vssd1 vssd1 vccd1 vccd1 _03819_ sky130_fd_sc_hd__a211o_1
XANTENNA__07805__S1 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1889 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07821_ _02610_ _02642_ _02706_ _02771_ vssd1 vssd1 vccd1 vccd1 _02772_ sky130_fd_sc_hd__and4_2
XANTENNA__07591__C1 _02503_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12467__B1 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07752_ net604 _02698_ _02674_ _01626_ vssd1 vssd1 vccd1 vccd1 _02703_ sky130_fd_sc_hd__o211a_1
XANTENNA__10312__A net1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07569__S0 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13581__CLK clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06703_ final_design.cpu.reg_window\[537\] final_design.cpu.reg_window\[569\] net931
+ vssd1 vssd1 vccd1 vccd1 _01654_ sky130_fd_sc_hd__mux2_1
X_07683_ _02628_ _02633_ net713 vssd1 vssd1 vccd1 vccd1 _02634_ sky130_fd_sc_hd__mux2_1
XANTENNA__11842__S net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09422_ net495 _04111_ vssd1 vssd1 vccd1 vccd1 _04341_ sky130_fd_sc_hd__nand2_4
XANTENNA__12219__B1 net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11690__A1 net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06634_ final_design.cpu.reg_window\[795\] final_design.cpu.reg_window\[827\] net943
+ vssd1 vssd1 vccd1 vccd1 _01585_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09353_ net479 _04083_ _04086_ _04269_ _04271_ vssd1 vssd1 vccd1 vccd1 _04272_ sky130_fd_sc_hd__o311a_1
XFILLER_0_19_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06565_ final_design.cpu.reg_window\[93\] final_design.cpu.reg_window\[125\] net949
+ vssd1 vssd1 vccd1 vccd1 _01516_ sky130_fd_sc_hd__mux2_1
XANTENNA__12234__A3 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout242_A _05875_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08304_ _03251_ _03252_ _03253_ _03254_ net674 net696 vssd1 vssd1 vccd1 vccd1 _03255_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_79_2901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06496_ final_design.cpu.reg_window\[670\] final_design.cpu.reg_window\[702\] net932
+ vssd1 vssd1 vccd1 vccd1 _01447_ sky130_fd_sc_hd__mux2_1
X_09284_ net606 net525 _01452_ _02422_ vssd1 vssd1 vccd1 vccd1 _04203_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_79_2912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07110__A2 net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08235_ final_design.cpu.reg_window\[715\] final_design.cpu.reg_window\[747\] net835
+ vssd1 vssd1 vccd1 vccd1 _03186_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout1151_A net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout507_A net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08166_ net707 _03110_ net722 vssd1 vssd1 vccd1 vccd1 _03117_ sky130_fd_sc_hd__o21a_1
XANTENNA__09938__A2 _04581_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14087__CLK clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07117_ final_design.cpu.reg_window\[331\] final_design.cpu.reg_window\[363\] net916
+ vssd1 vssd1 vccd1 vccd1 _02068_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08097_ final_design.cpu.reg_window\[12\] final_design.cpu.reg_window\[44\] net814
+ vssd1 vssd1 vccd1 vccd1 _03048_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout1037_X net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1901 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07048_ final_design.data_from_mem\[14\] net970 _01997_ vssd1 vssd1 vccd1 vccd1 _01999_
+ sky130_fd_sc_hd__o21ai_4
XFILLER_0_45_1480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout497_X net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout876_A _01687_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1204_X net1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input2_X net2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13924__CLK clknet_leaf_52_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08999_ _02452_ _02454_ vssd1 vssd1 vccd1 vccd1 _03934_ sky130_fd_sc_hd__or2_1
XFILLER_0_76_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07007__S net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10961_ net52 _05688_ vssd1 vssd1 vccd1 vccd1 _05689_ sky130_fd_sc_hd__and2_1
XANTENNA__11752__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09874__B2 _04222_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12700_ net1051 _06340_ vssd1 vssd1 vccd1 vccd1 _06341_ sky130_fd_sc_hd__or2_1
XANTENNA__09730__B _04113_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10484__A2 net250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13680_ clknet_leaf_36_clk _00911_ net1237 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[668\]
+ sky130_fd_sc_hd__dfrtp_1
X_10892_ _05600_ _05621_ vssd1 vssd1 vccd1 vccd1 _05623_ sky130_fd_sc_hd__nor2_1
XFILLER_0_74_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12631_ final_design.VGA_data_control.ready_data\[3\] net1022 net976 final_design.data_from_mem\[3\]
+ vssd1 vssd1 vccd1 vccd1 _06303_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_14_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12225__A3 net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12562_ _06225_ net354 net324 net2265 vssd1 vssd1 vccd1 vccd1 _01266_ sky130_fd_sc_hd__a22o_1
XFILLER_0_66_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13304__CLK clknet_leaf_63_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11984__A2 net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11513_ net1922 net215 net522 vssd1 vssd1 vccd1 vccd1 _00382_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_43_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12493_ _06153_ net357 net332 net2515 vssd1 vssd1 vccd1 vccd1 _01199_ sky130_fd_sc_hd__a22o_1
XFILLER_0_81_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_43_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14232_ net1286 vssd1 vssd1 vccd1 vccd1 gpio_out[10] sky130_fd_sc_hd__buf_2
X_11444_ net429 _06094_ vssd1 vssd1 vccd1 vccd1 _06095_ sky130_fd_sc_hd__nand2_4
XANTENNA__06581__S net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11197__B1 net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12880__Q final_design.data_from_mem\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14163_ clknet_leaf_17_clk _01337_ net1109 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.data_to_VGA\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09177__B net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11375_ net663 _03826_ net737 vssd1 vssd1 vccd1 vccd1 _06062_ sky130_fd_sc_hd__a21o_1
XANTENNA__13454__CLK clknet_leaf_43_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08601__A2 _03550_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13114_ clknet_leaf_5_clk _00345_ net1082 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[102\]
+ sky130_fd_sc_hd__dfrtp_1
X_10326_ net1465 net1009 net986 final_design.data_from_mem\[11\] vssd1 vssd1 vccd1
+ vccd1 _00083_ sky130_fd_sc_hd__a22o_1
XANTENNA_input58_X net58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14094_ clknet_leaf_14_clk _01291_ net1104 vssd1 vssd1 vccd1 vccd1 final_design.reqhand.instruction\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13045_ clknet_leaf_57_clk _00276_ net1144 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[33\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09157__A3 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10257_ final_design.uart.BAUD_counter\[21\] _05123_ vssd1 vssd1 vccd1 vccd1 _05124_
+ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_37_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09905__B _04821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1220 net1221 vssd1 vssd1 vccd1 vccd1 net1220 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_37_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09193__A _03617_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1231 net1232 vssd1 vssd1 vccd1 vccd1 net1231 sky130_fd_sc_hd__clkbuf_4
X_10188_ _05072_ _05077_ vssd1 vssd1 vccd1 vccd1 _05078_ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_33_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1242 net1244 vssd1 vssd1 vccd1 vccd1 net1242 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_79_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09314__A0 net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13947_ clknet_leaf_65_clk _01178_ net1070 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[935\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10475__A2 net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13878_ clknet_leaf_58_clk _01109_ net1126 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[866\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_27_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07971__S0 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12829_ net1350 vssd1 vssd1 vccd1 vccd1 _00270_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__09078__C1 net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09617__A1 _04066_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12216__A3 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1901 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1584 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_916 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11424__A1 net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11975__A2 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08020_ _02967_ _02968_ _02969_ _02970_ net679 net699 vssd1 vssd1 vccd1 vccd1 _02971_
+ sky130_fd_sc_hd__mux4_1
Xhold703 final_design.cpu.reg_window\[379\] vssd1 vssd1 vccd1 vccd1 net2045 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12958__RESET_B net1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold714 final_design.cpu.reg_window\[406\] vssd1 vssd1 vccd1 vccd1 net2056 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold725 final_design.cpu.reg_window\[476\] vssd1 vssd1 vccd1 vccd1 net2067 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold736 final_design.cpu.reg_window\[935\] vssd1 vssd1 vccd1 vccd1 net2078 sky130_fd_sc_hd__dlygate4sd3_1
Xhold747 final_design.cpu.reg_window\[213\] vssd1 vssd1 vccd1 vccd1 net2089 sky130_fd_sc_hd__dlygate4sd3_1
Xhold758 final_design.cpu.reg_window\[873\] vssd1 vssd1 vccd1 vccd1 net2100 sky130_fd_sc_hd__dlygate4sd3_1
Xhold769 final_design.cpu.reg_window\[930\] vssd1 vssd1 vccd1 vccd1 net2111 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07800__B1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09971_ net263 _04889_ vssd1 vssd1 vccd1 vccd1 _04890_ sky130_fd_sc_hd__nand2_1
XANTENNA__13947__CLK clknet_leaf_65_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11837__S net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload27_A clknet_leaf_38_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08922_ _02465_ _02466_ vssd1 vssd1 vccd1 vccd1 _03865_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_23_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_1705 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08853_ _03803_ vssd1 vssd1 vccd1 vccd1 _03804_ sky130_fd_sc_hd__inv_2
XANTENNA__11360__B1 net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout192_A _06031_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07804_ final_design.cpu.reg_window\[921\] final_design.cpu.reg_window\[953\] net851
+ vssd1 vssd1 vccd1 vccd1 _02755_ sky130_fd_sc_hd__mux2_1
XANTENNA__12971__CLK clknet_leaf_19_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1749 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08784_ final_design.CPU_instr_adr\[12\] _02064_ _03734_ vssd1 vssd1 vccd1 vccd1
+ _03735_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09390__X _04309_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07735_ net711 _02679_ net723 vssd1 vssd1 vccd1 vccd1 _02686_ sky130_fd_sc_hd__o21a_1
XFILLER_0_75_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09856__A1 _04773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout457_A _03551_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10466__A2 net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07666_ final_design.cpu.reg_window\[94\] final_design.cpu.reg_window\[126\] net856
+ vssd1 vssd1 vccd1 vccd1 _02617_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13327__CLK clknet_leaf_42_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09405_ net451 _04322_ _04323_ _04321_ vssd1 vssd1 vccd1 vccd1 _04324_ sky130_fd_sc_hd__a31o_1
X_06617_ final_design.reqhand.instruction\[28\] final_design.data_from_mem\[28\] net973
+ vssd1 vssd1 vccd1 vccd1 _01568_ sky130_fd_sc_hd__mux2_1
X_07597_ final_design.cpu.reg_window\[413\] final_design.cpu.reg_window\[445\] net870
+ vssd1 vssd1 vccd1 vccd1 _02548_ sky130_fd_sc_hd__mux2_1
XANTENNA__12207__A3 net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout245_X net245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout624_A net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11415__A1 net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09336_ _02673_ _03602_ _04254_ vssd1 vssd1 vccd1 vccd1 _04255_ sky130_fd_sc_hd__or3_1
XANTENNA__12612__B1 net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06548_ net743 net667 vssd1 vssd1 vccd1 vccd1 _01499_ sky130_fd_sc_hd__nor2_1
XFILLER_0_63_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1591 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11966__A2 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09267_ net73 net74 _04185_ vssd1 vssd1 vccd1 vccd1 _04186_ sky130_fd_sc_hd__or3_1
XFILLER_0_1_1444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout412_X net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13477__CLK clknet_leaf_49_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06479_ _01423_ _01424_ _01428_ _01429_ net779 net791 vssd1 vssd1 vccd1 vccd1 _01430_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout1154_X net1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08218_ final_design.cpu.reg_window\[331\] final_design.cpu.reg_window\[363\] net835
+ vssd1 vssd1 vccd1 vccd1 _03169_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09198_ net495 _04054_ vssd1 vssd1 vccd1 vccd1 _04117_ sky130_fd_sc_hd__nand2_2
XFILLER_0_44_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11179__B1 net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11718__A2 net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08149_ net611 _03096_ _03098_ net540 vssd1 vssd1 vccd1 vccd1 _03100_ sky130_fd_sc_hd__a211oi_2
XANTENNA__09792__A0 net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_1428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11160_ final_design.data_from_mem\[2\] net251 _05855_ _05872_ vssd1 vssd1 vccd1
+ vccd1 _05873_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout781_X net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1439 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11747__S net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout879_X net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10111_ final_design.VGA_data_control.v_count\[2\] _05019_ final_design.VGA_data_control.v_count\[3\]
+ vssd1 vssd1 vccd1 vccd1 _05024_ sky130_fd_sc_hd__a21o_1
X_11091_ _05799_ _05810_ _05812_ net59 vssd1 vssd1 vccd1 vccd1 _05813_ sky130_fd_sc_hd__a31oi_1
X_10042_ _04198_ _04253_ _04329_ _04960_ vssd1 vssd1 vccd1 vccd1 _04961_ sky130_fd_sc_hd__and4_2
XFILLER_0_41_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold30 final_design.cpu.reg_window\[20\] vssd1 vssd1 vccd1 vccd1 net1372 sky130_fd_sc_hd__dlygate4sd3_1
Xhold41 final_design.cpu.reg_window\[4\] vssd1 vssd1 vccd1 vccd1 net1383 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_51_1960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold52 final_design.VGA_data_control.data_to_VGA\[0\] vssd1 vssd1 vccd1 vccd1 net1394
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14102__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold63 net127 vssd1 vssd1 vccd1 vccd1 net1405 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold74 net130 vssd1 vssd1 vccd1 vccd1 net1416 sky130_fd_sc_hd__dlygate4sd3_1
Xhold85 net126 vssd1 vssd1 vccd1 vccd1 net1427 sky130_fd_sc_hd__dlygate4sd3_1
Xhold96 net101 vssd1 vssd1 vccd1 vccd1 net1438 sky130_fd_sc_hd__dlygate4sd3_1
X_13801_ clknet_leaf_33_clk _01032_ net1231 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[789\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input18_A DAT_I[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10887__A net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11993_ _05869_ net242 net627 vssd1 vssd1 vccd1 vccd1 _06258_ sky130_fd_sc_hd__and3_1
XANTENNA__11482__S net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13732_ clknet_leaf_54_clk _00963_ net1179 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[720\]
+ sky130_fd_sc_hd__dfrtp_1
X_10944_ _05542_ _05603_ _05668_ vssd1 vssd1 vccd1 vccd1 _05672_ sky130_fd_sc_hd__or3_1
XANTENNA__10457__A2 net1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11654__A1 net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08357__A net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12875__Q final_design.data_from_mem\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13663_ clknet_leaf_8_clk _00894_ net1153 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[651\]
+ sky130_fd_sc_hd__dfrtp_1
X_10875_ _05602_ _05605_ vssd1 vssd1 vccd1 vccd1 _05607_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_45_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12614_ net1398 net1412 _05080_ vssd1 vssd1 vccd1 vccd1 _01307_ sky130_fd_sc_hd__mux2_1
X_13594_ clknet_leaf_64_clk _00825_ net1075 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[582\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_41_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11214__C _05920_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12545_ _06208_ net344 net322 net2217 vssd1 vssd1 vccd1 vccd1 _01249_ sky130_fd_sc_hd__a22o_1
XFILLER_0_13_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08804__B _01722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06833__A1 net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12476_ _06136_ net347 net330 net1958 vssd1 vssd1 vccd1 vccd1 _01182_ sky130_fd_sc_hd__a22o_1
XFILLER_0_65_1620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12844__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14215_ net1273 vssd1 vssd1 vccd1 vccd1 gpio_oeb[27] sky130_fd_sc_hd__buf_2
X_11427_ net1879 net204 net313 vssd1 vssd1 vccd1 vccd1 _00324_ sky130_fd_sc_hd__mux2_1
XANTENNA_5 _05934_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14146_ clknet_leaf_20_clk _01320_ net1162 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.data_to_VGA\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_39_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11358_ net661 _03840_ net733 vssd1 vssd1 vccd1 vccd1 _06047_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_39_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10393__A1 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10393__B2 net167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10309_ net1048 _05155_ _05157_ _05162_ vssd1 vssd1 vccd1 vccd1 _05163_ sky130_fd_sc_hd__o31ai_1
XANTENNA__09194__Y _04113_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10414__X _05190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14077_ clknet_leaf_13_clk _01274_ net1089 vssd1 vssd1 vccd1 vccd1 final_design.uart.working_data\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_11289_ _01909_ net642 _05985_ _05986_ net658 vssd1 vssd1 vccd1 vccd1 _05987_ sky130_fd_sc_hd__a221o_1
XFILLER_0_20_1214 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13028_ clknet_leaf_54_clk _00259_ net1179 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[16\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1050 final_design.VGA_data_control.h_count\[1\] vssd1 vssd1 vccd1 vccd1 net1050
+ sky130_fd_sc_hd__clkbuf_4
Xfanout1061 net1069 vssd1 vssd1 vccd1 vccd1 net1061 sky130_fd_sc_hd__clkbuf_4
Xfanout1072 net1118 vssd1 vssd1 vccd1 vccd1 net1072 sky130_fd_sc_hd__clkbuf_4
Xfanout1083 net1085 vssd1 vssd1 vccd1 vccd1 net1083 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_59_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1094 net1096 vssd1 vssd1 vccd1 vccd1 net1094 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09838__A1 net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07520_ _01662_ _02470_ _01631_ _01632_ vssd1 vssd1 vccd1 vccd1 _02471_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_7_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07451_ final_design.cpu.reg_window\[0\] final_design.cpu.reg_window\[32\] net895
+ vssd1 vssd1 vccd1 vccd1 _02402_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07382_ final_design.cpu.reg_window\[322\] final_design.cpu.reg_window\[354\] net922
+ vssd1 vssd1 vccd1 vccd1 _02333_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_1917 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09121_ _01409_ net992 vssd1 vssd1 vccd1 vccd1 _04040_ sky130_fd_sc_hd__nor2_4
XANTENNA__11948__A2 net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07077__A1 final_design.data_from_mem\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08714__B _01660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09052_ final_design.CPU_instr_adr\[9\] _03787_ vssd1 vssd1 vccd1 vccd1 _03981_ sky130_fd_sc_hd__xor2_1
XFILLER_0_5_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06515__A final_design.data_from_mem\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08003_ _02950_ _02951_ _02952_ _02953_ net682 net702 vssd1 vssd1 vccd1 vccd1 _02954_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_41_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold500 final_design.cpu.reg_window\[692\] vssd1 vssd1 vccd1 vccd1 net1842 sky130_fd_sc_hd__dlygate4sd3_1
Xhold511 final_design.cpu.reg_window\[274\] vssd1 vssd1 vccd1 vccd1 net1853 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout205_A net206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold522 final_design.cpu.reg_window\[744\] vssd1 vssd1 vccd1 vccd1 net1864 sky130_fd_sc_hd__dlygate4sd3_1
Xhold533 final_design.cpu.reg_window\[920\] vssd1 vssd1 vccd1 vccd1 net1875 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_1726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09826__A net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold544 final_design.cpu.reg_window\[1022\] vssd1 vssd1 vccd1 vccd1 net1886 sky130_fd_sc_hd__dlygate4sd3_1
Xhold555 final_design.cpu.reg_window\[361\] vssd1 vssd1 vccd1 vccd1 net1897 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06588__B1 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold566 final_design.cpu.reg_window\[750\] vssd1 vssd1 vccd1 vccd1 net1908 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11581__B1 net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold577 final_design.cpu.reg_window\[793\] vssd1 vssd1 vccd1 vccd1 net1919 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07785__C1 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_2071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold588 final_design.cpu.reg_window\[894\] vssd1 vssd1 vccd1 vccd1 net1930 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_55_2082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14125__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09954_ _03486_ net440 _04872_ net450 vssd1 vssd1 vccd1 vccd1 _04873_ sky130_fd_sc_hd__a211o_1
Xhold599 final_design.cpu.reg_window\[786\] vssd1 vssd1 vccd1 vccd1 net1941 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_55_2093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1114_A net1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08905_ net625 _03847_ vssd1 vssd1 vccd1 vccd1 _03850_ sky130_fd_sc_hd__nor2_1
X_09885_ _03522_ _03640_ vssd1 vssd1 vccd1 vccd1 _04804_ sky130_fd_sc_hd__xor2_1
Xhold1200 final_design.cpu.reg_window\[51\] vssd1 vssd1 vccd1 vccd1 net2542 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout574_A net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1211 wb_manage.curr_state\[2\] vssd1 vssd1 vccd1 vccd1 net2553 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout195_X net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08836_ final_design.CPU_instr_adr\[8\] _03786_ vssd1 vssd1 vccd1 vccd1 _03787_ sky130_fd_sc_hd__and2_1
X_08767_ final_design.CPU_instr_adr\[0\] _02425_ _03716_ _03714_ vssd1 vssd1 vccd1
+ vccd1 _03718_ sky130_fd_sc_hd__a31o_1
XANTENNA__09829__A1 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout362_X net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13580__RESET_B net1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout839_A net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11636__A1 net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07718_ _01599_ net605 vssd1 vssd1 vccd1 vccd1 _02669_ sky130_fd_sc_hd__and2_1
X_08698_ _01486_ _03646_ _03648_ vssd1 vssd1 vccd1 vccd1 _03649_ sky130_fd_sc_hd__nand3_4
XANTENNA__07935__S0 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07081__A _02026_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07649_ _02596_ _02597_ _02598_ _02599_ net687 net694 vssd1 vssd1 vccd1 vccd1 _02600_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_7_1675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout627_X net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10660_ _05400_ _05401_ vssd1 vssd1 vccd1 vccd1 _05402_ sky130_fd_sc_hd__nand2_1
XANTENNA__08905__A net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12867__CLK clknet_leaf_25_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11939__A2 net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09319_ net528 net452 vssd1 vssd1 vccd1 vccd1 _04238_ sky130_fd_sc_hd__nand2_1
X_10591_ _05315_ _05318_ _05335_ vssd1 vssd1 vccd1 vccd1 _05336_ sky130_fd_sc_hd__and3_1
XANTENNA__10298__S1 net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12330_ net671 net647 _06268_ net361 net2011 vssd1 vssd1 vccd1 vccd1 _01043_ sky130_fd_sc_hd__a32o_1
XFILLER_0_17_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07020__S net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06910__S1 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12261_ net578 _06190_ net510 net374 net1491 vssd1 vssd1 vccd1 vccd1 _00977_ sky130_fd_sc_hd__a32o_1
XANTENNA__08112__S0 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14000_ clknet_leaf_33_clk _01231_ net1239 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[988\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_62_1815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_1372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11212_ net645 _05918_ _05916_ net653 vssd1 vssd1 vccd1 vccd1 _05919_ sky130_fd_sc_hd__a211o_1
X_12192_ net2426 net183 net382 vssd1 vssd1 vccd1 vccd1 _00911_ sky130_fd_sc_hd__mux2_1
XANTENNA__10375__B2 final_design.data_from_mem\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11477__S net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11143_ _04939_ net651 net588 _05857_ vssd1 vssd1 vccd1 vccd1 _05858_ sky130_fd_sc_hd__o211a_1
X_11074_ _05793_ _05794_ _05796_ net1034 net1379 vssd1 vssd1 vccd1 vccd1 _00202_ sky130_fd_sc_hd__a32o_1
XFILLER_0_37_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10025_ _04108_ _04398_ net318 vssd1 vssd1 vccd1 vccd1 _04944_ sky130_fd_sc_hd__o21a_1
XFILLER_0_37_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12419__A3 net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13642__CLK clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12101__S net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_47_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10410__A _03352_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11976_ _06178_ net283 net406 net2075 vssd1 vssd1 vccd1 vccd1 _00709_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_47_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13715_ clknet_leaf_40_clk _00946_ net1206 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[703\]
+ sky130_fd_sc_hd__dfrtp_1
X_10927_ _05654_ _05655_ vssd1 vssd1 vccd1 vccd1 _05656_ sky130_fd_sc_hd__nor2_1
XFILLER_0_54_1376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13646_ clknet_leaf_44_clk _00877_ net1208 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[634\]
+ sky130_fd_sc_hd__dfrtp_1
X_10858_ _05588_ _05589_ _05568_ vssd1 vssd1 vccd1 vccd1 _05590_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_6_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13792__CLK clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12052__A1 net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13577_ clknet_leaf_37_clk _00808_ net1228 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[565\]
+ sky130_fd_sc_hd__dfrtp_1
X_10789_ _05508_ _05524_ vssd1 vssd1 vccd1 vccd1 _05525_ sky130_fd_sc_hd__nor2_1
XFILLER_0_26_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08351__S0 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10602__A2 net1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12528_ _06190_ net353 net328 net1532 vssd1 vssd1 vccd1 vccd1 _01233_ sky130_fd_sc_hd__a22o_1
XFILLER_0_48_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_13 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14148__CLK clknet_leaf_19_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12459_ net1957 net185 net337 vssd1 vssd1 vccd1 vccd1 _01166_ sky130_fd_sc_hd__mux2_1
XANTENNA__13022__CLK clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12355__A2 net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10366__B2 final_design.data_from_mem\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11563__B1 net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14129_ clknet_leaf_20_clk final_design.vga.v_next_state\[0\] net1159 vssd1 vssd1
+ vccd1 vccd1 final_design.vga.v_current_state\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout309 _06095_ vssd1 vssd1 vccd1 vccd1 net309 sky130_fd_sc_hd__clkbuf_8
XANTENNA__07782__A2 _02731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06951_ final_design.cpu.reg_window\[721\] final_design.cpu.reg_window\[753\] net928
+ vssd1 vssd1 vccd1 vccd1 _01902_ sky130_fd_sc_hd__mux2_1
XANTENNA__11315__B1 net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1833 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09670_ _02804_ net445 net442 _02800_ _04588_ vssd1 vssd1 vccd1 vccd1 _04589_ sky130_fd_sc_hd__o221a_1
XANTENNA__11866__B2 net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06882_ final_design.cpu.reg_window\[19\] final_design.cpu.reg_window\[51\] net911
+ vssd1 vssd1 vccd1 vccd1 _01833_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_1877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08621_ _03198_ _03571_ _03570_ vssd1 vssd1 vccd1 vccd1 _03572_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_59_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08709__B _01599_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11618__A1 net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08552_ final_design.cpu.reg_window\[961\] final_design.cpu.reg_window\[993\] net833
+ vssd1 vssd1 vccd1 vccd1 _03503_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_1574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07503_ _01969_ _01970_ vssd1 vssd1 vccd1 vccd1 _02454_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_33_1416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08483_ final_design.cpu.reg_window\[195\] final_design.cpu.reg_window\[227\] net820
+ vssd1 vssd1 vccd1 vccd1 _03434_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_2351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_2362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_2373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07434_ final_design.cpu.reg_window\[577\] final_design.cpu.reg_window\[609\] net912
+ vssd1 vssd1 vccd1 vccd1 _02385_ sky130_fd_sc_hd__mux2_1
XANTENNA__08590__S0 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07365_ final_design.cpu.reg_window\[899\] final_design.cpu.reg_window\[931\] net904
+ vssd1 vssd1 vccd1 vccd1 _02316_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_1796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout322_A net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1064_A net1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11151__A net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09104_ _02430_ _04024_ _04025_ net619 vssd1 vssd1 vccd1 vccd1 _04026_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_73_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12594__A2 net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07296_ _02243_ _02244_ _02245_ _02246_ net770 net789 vssd1 vssd1 vccd1 vccd1 _02247_
+ sky130_fd_sc_hd__mux4_1
X_09035_ _03963_ _03965_ net255 vssd1 vssd1 vccd1 vccd1 _03966_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_57_2144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout208_X net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07775__S net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_2155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_2789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12346__A2 net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_2166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold330 final_design.cpu.reg_window\[229\] vssd1 vssd1 vccd1 vccd1 net1672 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_53_2008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10357__A1 net30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13515__CLK clknet_leaf_38_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold341 final_design.cpu.reg_window\[204\] vssd1 vssd1 vccd1 vccd1 net1683 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_53_2019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10357__B2 final_design.data_from_mem\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold352 final_design.cpu.reg_window\[773\] vssd1 vssd1 vccd1 vccd1 net1694 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout691_A net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold363 final_design.cpu.reg_window\[580\] vssd1 vssd1 vccd1 vccd1 net1705 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout789_A net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold374 final_design.cpu.reg_window\[842\] vssd1 vssd1 vccd1 vccd1 net1716 sky130_fd_sc_hd__dlygate4sd3_1
Xhold385 final_design.cpu.reg_window\[82\] vssd1 vssd1 vccd1 vccd1 net1727 sky130_fd_sc_hd__dlygate4sd3_1
Xhold396 final_design.cpu.reg_window\[174\] vssd1 vssd1 vccd1 vccd1 net1738 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout810 net811 vssd1 vssd1 vccd1 vccd1 net810 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout1117_X net1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout821 net823 vssd1 vssd1 vccd1 vccd1 net821 sky130_fd_sc_hd__clkbuf_4
Xfanout832 net833 vssd1 vssd1 vccd1 vccd1 net832 sky130_fd_sc_hd__clkbuf_4
X_09937_ _03388_ net438 _04109_ _04309_ _04855_ vssd1 vssd1 vccd1 vccd1 _04856_ sky130_fd_sc_hd__o221a_1
Xfanout843 net847 vssd1 vssd1 vccd1 vccd1 net843 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11306__B1 _06001_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout956_A net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout577_X net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout854 net872 vssd1 vssd1 vccd1 vccd1 net854 sky130_fd_sc_hd__clkbuf_4
Xfanout865 net872 vssd1 vssd1 vccd1 vccd1 net865 sky130_fd_sc_hd__buf_2
XANTENNA__13665__CLK clknet_leaf_47_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout876 _01687_ vssd1 vssd1 vccd1 vccd1 net876 sky130_fd_sc_hd__buf_6
Xfanout887 net890 vssd1 vssd1 vccd1 vccd1 net887 sky130_fd_sc_hd__clkbuf_4
X_09868_ net728 _04772_ _04786_ vssd1 vssd1 vccd1 vccd1 _04787_ sky130_fd_sc_hd__and3_1
Xfanout898 net899 vssd1 vssd1 vccd1 vccd1 net898 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_5_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1030 final_design.cpu.reg_window\[741\] vssd1 vssd1 vccd1 vccd1 net2372 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11857__B2 net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1041 final_design.cpu.reg_window\[810\] vssd1 vssd1 vccd1 vccd1 net2383 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_57_1917 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1052 final_design.uart.BAUD_counter\[10\] vssd1 vssd1 vccd1 vccd1 net2394 sky130_fd_sc_hd__dlygate4sd3_1
X_08819_ _03668_ _03769_ vssd1 vssd1 vccd1 vccd1 _03770_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_5_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1063 final_design.cpu.reg_window\[102\] vssd1 vssd1 vccd1 vccd1 net2405 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12789__20_A clknet_leaf_30_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1074 final_design.cpu.reg_window\[113\] vssd1 vssd1 vccd1 vccd1 net2416 sky130_fd_sc_hd__dlygate4sd3_1
X_09799_ _03455_ _03557_ _03560_ _03457_ _03424_ vssd1 vssd1 vccd1 vccd1 _04718_ sky130_fd_sc_hd__o311a_1
XANTENNA_fanout744_X net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1085 final_design.VGA_adr\[0\] vssd1 vssd1 vccd1 vccd1 net2427 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13008__RESET_B net1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11830_ net199 net2004 net264 vssd1 vssd1 vccd1 vccd1 _00582_ sky130_fd_sc_hd__mux2_1
Xhold1096 final_design.cpu.reg_window\[301\] vssd1 vssd1 vccd1 vccd1 net2438 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12282__A1 net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11761_ net189 net2118 net419 vssd1 vssd1 vccd1 vccd1 _00524_ sky130_fd_sc_hd__mux2_1
XANTENNA__11760__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13500_ clknet_leaf_2_clk _00731_ net1077 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[488\]
+ sky130_fd_sc_hd__dfrtp_1
X_10712_ _05449_ _05450_ vssd1 vssd1 vccd1 vccd1 _05451_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_36_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06707__X _01658_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11692_ net561 net420 _06204_ net294 net1630 vssd1 vssd1 vccd1 vccd1 _00477_ sky130_fd_sc_hd__a32o_1
XFILLER_0_3_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13431_ clknet_leaf_6_clk _00662_ net1130 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[419\]
+ sky130_fd_sc_hd__dfrtp_1
X_10643_ _05362_ _05383_ vssd1 vssd1 vccd1 vccd1 _05386_ sky130_fd_sc_hd__and2_1
XFILLER_0_3_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13045__CLK clknet_leaf_57_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10045__B1 _04421_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12585__A2 net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input85_A memory_size[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13362_ clknet_leaf_39_clk _00593_ net1206 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[350\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_36_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10574_ final_design.CPU_instr_adr\[6\] _05319_ net1053 vssd1 vssd1 vccd1 vccd1 _05320_
+ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_5_clk_A clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09450__A2 net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10596__B2 net1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11793__B1 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12313_ net2186 net222 net365 vssd1 vssd1 vccd1 vccd1 _01027_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_20_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13293_ clknet_leaf_44_clk _00524_ net1209 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[281\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_39_Left_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_20_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12337__A2 net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13195__CLK clknet_leaf_38_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12244_ net561 _06174_ net498 net372 net1476 vssd1 vssd1 vccd1 vccd1 _00961_ sky130_fd_sc_hd__a32o_1
XANTENNA__11545__B1 net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12175_ net1828 net214 net381 vssd1 vssd1 vccd1 vccd1 _00894_ sky130_fd_sc_hd__mux2_1
XANTENNA__08961__A1 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11126_ _01487_ net654 net1013 vssd1 vssd1 vccd1 vccd1 _05841_ sky130_fd_sc_hd__a21oi_4
X_11057_ net89 net1047 vssd1 vssd1 vccd1 vccd1 _05780_ sky130_fd_sc_hd__nor2_1
XANTENNA__09913__B _04087_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10008_ _03642_ _04045_ _04089_ _03641_ _04926_ vssd1 vssd1 vccd1 vccd1 _04927_ sky130_fd_sc_hd__a221o_1
XFILLER_0_64_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_1416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_48_Left_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07978__A1_N net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11959_ _06160_ net282 net405 net2330 vssd1 vssd1 vccd1 vccd1 _00692_ sky130_fd_sc_hd__a22o_1
XFILLER_0_47_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09140__S net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13629_ clknet_leaf_2_clk _00860_ net1068 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[617\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08229__B1 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07150_ net538 _02098_ vssd1 vssd1 vccd1 vccd1 _02101_ sky130_fd_sc_hd__and2_1
XFILLER_0_82_682 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13538__CLK clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_57_Left_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07081_ _02026_ _02031_ vssd1 vssd1 vccd1 vccd1 _02032_ sky130_fd_sc_hd__and2_1
XFILLER_0_80_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09729__B1 net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10339__B2 final_design.data_from_mem\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1745 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_2620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_2631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07204__A1 net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_2642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13688__CLK clknet_leaf_65_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09744__A3 _02091_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1789 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07983_ net613 _02929_ _02931_ _01908_ vssd1 vssd1 vccd1 vccd1 _02934_ sky130_fd_sc_hd__a211o_1
XANTENNA__11845__S net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09722_ net542 net541 net540 net539 net454 net464 vssd1 vssd1 vccd1 vccd1 _04641_
+ sky130_fd_sc_hd__mux4_1
X_06934_ final_design.cpu.reg_window\[465\] final_design.cpu.reg_window\[497\] net928
+ vssd1 vssd1 vccd1 vccd1 _01885_ sky130_fd_sc_hd__mux2_1
XANTENNA__12500__A2 net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09315__S net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09653_ net78 _04188_ vssd1 vssd1 vccd1 vccd1 _04572_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_69_2560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06865_ _01381_ net1040 net994 net991 vssd1 vssd1 vccd1 vccd1 _01816_ sky130_fd_sc_hd__or4_4
XANTENNA_fanout272_A net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_2571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_1549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_65_2413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08604_ _03520_ _03521_ _03554_ vssd1 vssd1 vccd1 vccd1 _03555_ sky130_fd_sc_hd__o21ai_2
XTAP_TAPCELL_ROW_65_2424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_2435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09584_ _04144_ _04153_ _04154_ _04155_ vssd1 vssd1 vccd1 vccd1 _04503_ sky130_fd_sc_hd__a31o_1
X_06796_ final_design.cpu.reg_window\[918\] final_design.cpu.reg_window\[950\] net919
+ vssd1 vssd1 vccd1 vccd1 _01747_ sky130_fd_sc_hd__mux2_1
X_08535_ net608 _03481_ _03482_ net528 vssd1 vssd1 vccd1 vccd1 _03486_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_38_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13068__CLK clknet_leaf_47_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout537_A _02126_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07366__S1 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08466_ _02297_ net609 vssd1 vssd1 vccd1 vccd1 _03417_ sky130_fd_sc_hd__or2_1
XFILLER_0_49_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12973__Q final_design.CPU_instr_adr\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07417_ final_design.cpu.reg_window\[385\] final_design.cpu.reg_window\[417\] net922
+ vssd1 vssd1 vccd1 vccd1 _02368_ sky130_fd_sc_hd__mux2_1
X_08397_ final_design.cpu.reg_window\[582\] final_design.cpu.reg_window\[614\] net821
+ vssd1 vssd1 vccd1 vccd1 _03348_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout704_A net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout325_X net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_2206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07348_ _02294_ _02297_ vssd1 vssd1 vccd1 vccd1 _02299_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_59_2217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_2228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10578__A1 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_2239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_1599 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07279_ final_design.cpu.reg_window\[966\] final_design.cpu.reg_window\[998\] net904
+ vssd1 vssd1 vccd1 vccd1 _02230_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout1234_X net1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12905__CLK clknet_leaf_60_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09018_ _03950_ vssd1 vssd1 vccd1 vccd1 _03951_ sky130_fd_sc_hd__inv_2
XFILLER_0_27_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10290_ final_design.VGA_data_control.data_to_VGA\[19\] final_design.VGA_data_control.data_to_VGA\[18\]
+ final_design.VGA_data_control.data_to_VGA\[17\] final_design.VGA_data_control.data_to_VGA\[16\]
+ net1050 net1049 vssd1 vssd1 vccd1 vccd1 _05144_ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout694_X net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09196__A1 _02545_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold160 final_design.cpu.reg_window\[713\] vssd1 vssd1 vccd1 vccd1 net1502 sky130_fd_sc_hd__dlygate4sd3_1
Xhold171 final_design.cpu.reg_window\[735\] vssd1 vssd1 vccd1 vccd1 net1513 sky130_fd_sc_hd__dlygate4sd3_1
Xhold182 final_design.VGA_data_control.ready_data\[13\] vssd1 vssd1 vccd1 vccd1 net1524
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold193 final_design.VGA_data_control.ready_data\[9\] vssd1 vssd1 vccd1 vccd1 net1535
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout959_X net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout640 _06093_ vssd1 vssd1 vccd1 vccd1 net640 sky130_fd_sc_hd__buf_4
XANTENNA__11755__S net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout651 net652 vssd1 vssd1 vccd1 vccd1 net651 sky130_fd_sc_hd__clkbuf_4
Xfanout662 net663 vssd1 vssd1 vccd1 vccd1 net662 sky130_fd_sc_hd__clkbuf_4
X_13980_ clknet_leaf_3_clk _01211_ net1079 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[968\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout673 _02328_ vssd1 vssd1 vccd1 vccd1 net673 sky130_fd_sc_hd__buf_2
Xfanout684 net689 vssd1 vssd1 vccd1 vccd1 net684 sky130_fd_sc_hd__buf_4
X_12931_ clknet_leaf_31_clk _00169_ net1233 vssd1 vssd1 vccd1 vccd1 net154 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12862_ clknet_leaf_20_clk _00100_ net1158 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.ready_data\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_34_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07821__X _02772_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11813_ net242 net2236 net265 vssd1 vssd1 vccd1 vccd1 _00565_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12255__A1 net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08554__S0 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11744_ net221 net2033 net416 vssd1 vssd1 vccd1 vccd1 _00507_ sky130_fd_sc_hd__mux2_1
XANTENNA__12883__Q final_design.data_from_mem\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11675_ net566 net241 net627 vssd1 vssd1 vccd1 vccd1 _06196_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_12_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_12_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_1821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13414_ clknet_leaf_51_clk _00645_ net1170 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[402\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12558__A2 net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10626_ net99 final_design.VGA_adr\[7\] vssd1 vssd1 vccd1 vccd1 _05369_ sky130_fd_sc_hd__nand2_1
XFILLER_0_64_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13345_ clknet_leaf_48_clk _00576_ net1200 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[333\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_1827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10557_ _05267_ _05285_ _05303_ _05283_ vssd1 vssd1 vccd1 vccd1 _05304_ sky130_fd_sc_hd__o211a_1
XFILLER_0_64_1729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13830__CLK clknet_leaf_51_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13276_ clknet_leaf_5_clk _00507_ net1078 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[264\]
+ sky130_fd_sc_hd__dfrtp_1
X_10488_ net1018 net1057 vssd1 vssd1 vccd1 vccd1 _05238_ sky130_fd_sc_hd__xnor2_1
X_12227_ net578 _06155_ net510 net378 net1639 vssd1 vssd1 vccd1 vccd1 _00945_ sky130_fd_sc_hd__a32o_1
XANTENNA__09726__A3 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09282__S1 net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09924__A net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12158_ net183 net2489 net386 vssd1 vssd1 vccd1 vccd1 _00879_ sky130_fd_sc_hd__mux2_1
XANTENNA__06945__B1 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13980__CLK clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_36 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11109_ net1539 net1034 net1003 _05829_ vssd1 vssd1 vccd1 vccd1 _00204_ sky130_fd_sc_hd__a22o_1
XFILLER_0_75_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12089_ net581 _06061_ net512 net394 net1720 vssd1 vssd1 vccd1 vccd1 _00814_ sky130_fd_sc_hd__a32o_1
XANTENNA__11297__A2 net235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13210__CLK clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06650_ _01596_ _01599_ vssd1 vssd1 vccd1 vccd1 _01601_ sky130_fd_sc_hd__or2_1
XFILLER_0_73_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_1680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06581_ final_design.cpu.reg_window\[541\] final_design.cpu.reg_window\[573\] net951
+ vssd1 vssd1 vccd1 vccd1 _01532_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_1582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08320_ final_design.cpu.reg_window\[200\] final_design.cpu.reg_window\[232\] net813
+ vssd1 vssd1 vccd1 vccd1 _03271_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_50_clk_X clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13360__CLK clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08251_ final_design.cpu.reg_window\[266\] final_design.cpu.reg_window\[298\] net818
+ vssd1 vssd1 vccd1 vccd1 _03202_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_1829 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12928__CLK clknet_leaf_47_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07202_ _02149_ _02150_ _02151_ _02152_ net764 net785 vssd1 vssd1 vccd1 vccd1 _02153_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__12549__A2 net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08182_ net612 net526 _03131_ net543 vssd1 vssd1 vccd1 vccd1 _03133_ sky130_fd_sc_hd__a211oi_2
XANTENNA__11757__A0 net196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_2840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07425__A1 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07133_ _02080_ _02081_ _02082_ _02083_ net768 net788 vssd1 vssd1 vccd1 vccd1 _02084_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_77_2851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_65_clk_X clknet_leaf_65_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_73_2704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07064_ final_design.cpu.reg_window\[589\] final_design.cpu.reg_window\[621\] net935
+ vssd1 vssd1 vccd1 vccd1 _02015_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_12_Right_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout487_A net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07966_ net721 _02916_ net723 vssd1 vssd1 vccd1 vccd1 _02917_ sky130_fd_sc_hd__o21ai_1
XANTENNA__09045__S net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_2508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09705_ _03102_ net446 _04617_ _04623_ vssd1 vssd1 vccd1 vccd1 _04624_ sky130_fd_sc_hd__o211a_1
X_06917_ net763 _01867_ net747 vssd1 vssd1 vccd1 vccd1 _01868_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07036__S0 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08689__B1 _03523_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07897_ final_design.cpu.reg_window\[151\] final_design.cpu.reg_window\[183\] net849
+ vssd1 vssd1 vccd1 vccd1 _02848_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout275_X net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout654_A net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09350__A1 net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07587__S1 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09636_ _04107_ _04277_ _04116_ vssd1 vssd1 vccd1 vccd1 _04555_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_39_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09840__Y _04759_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06848_ final_design.cpu.reg_window\[212\] final_design.cpu.reg_window\[244\] net947
+ vssd1 vssd1 vccd1 vccd1 _01799_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_21_Right_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07361__B1 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13703__CLK clknet_leaf_63_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09567_ net551 net550 net549 net548 net453 net463 vssd1 vssd1 vccd1 vccd1 _04486_
+ sky130_fd_sc_hd__mux4_1
X_06779_ _01726_ _01727_ _01728_ _01729_ net770 net789 vssd1 vssd1 vccd1 vccd1 _01730_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout821_A net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout442_X net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout919_A net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08518_ net710 _03462_ net724 vssd1 vssd1 vccd1 vccd1 _03469_ sky130_fd_sc_hd__o21a_1
XANTENNA_clkbuf_leaf_18_clk_X clknet_leaf_18_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09498_ _04074_ _04403_ _04416_ _04400_ vssd1 vssd1 vccd1 vccd1 _04417_ sky130_fd_sc_hd__o211a_1
XFILLER_0_66_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11996__B1 net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08310__C1 net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08449_ final_design.cpu.reg_window\[132\] final_design.cpu.reg_window\[164\] net821
+ vssd1 vssd1 vccd1 vccd1 _03400_ sky130_fd_sc_hd__mux2_1
XANTENNA__11323__B net196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout707_X net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13853__CLK clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11460_ net221 net638 vssd1 vssd1 vccd1 vccd1 _06103_ sky130_fd_sc_hd__and2_1
XFILLER_0_68_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11748__A0 net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_5_0_clk_X clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10411_ net250 _05188_ net1030 net1384 vssd1 vssd1 vccd1 vccd1 _00147_ sky130_fd_sc_hd__a2bb2o_1
X_11391_ net661 _03807_ _01491_ vssd1 vssd1 vccd1 vccd1 _06076_ sky130_fd_sc_hd__o21ai_1
XPHY_EDGE_ROW_30_Right_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13130_ clknet_leaf_61_clk _00361_ net1140 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[118\]
+ sky130_fd_sc_hd__dfrtp_1
X_10342_ net1496 net1010 net987 final_design.data_from_mem\[27\] vssd1 vssd1 vccd1
+ vccd1 _00099_ sky130_fd_sc_hd__a22o_1
XANTENNA__08124__S net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13061_ clknet_leaf_49_clk _00292_ net1184 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[49\]
+ sky130_fd_sc_hd__dfrtp_1
X_10273_ final_design.uart.BAUD_counter\[27\] _05133_ vssd1 vssd1 vccd1 vccd1 _05134_
+ sky130_fd_sc_hd__and2_1
X_12012_ _06214_ net292 net402 net2114 vssd1 vssd1 vccd1 vccd1 _00743_ sky130_fd_sc_hd__a22o_1
XANTENNA__07719__A2 _02668_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08916__A1 net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11993__B net242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input48_A mem_adr_start[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07275__S0 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13023__RESET_B net1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11485__S net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13233__CLK clknet_leaf_34_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout470 _03485_ vssd1 vssd1 vccd1 vccd1 net470 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_79_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_35_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout481 net482 vssd1 vssd1 vccd1 vccd1 net481 sky130_fd_sc_hd__buf_2
XANTENNA__12878__Q final_design.data_from_mem\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout492 net493 vssd1 vssd1 vccd1 vccd1 net492 sky130_fd_sc_hd__buf_2
XANTENNA__12476__A1 _06136_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11279__A2 _05977_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13963_ clknet_leaf_53_clk _01194_ net1185 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[951\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_31_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10402__B _05181_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12914_ clknet_leaf_28_clk _00152_ net1193 vssd1 vssd1 vccd1 vccd1 net136 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_31_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13894_ clknet_leaf_52_clk _01125_ net1174 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[882\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_1528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13383__CLK clknet_leaf_58_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09892__A2 net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12845_ clknet_leaf_14_clk _00083_ net1107 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.ready_data\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_914 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1733 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06608__A net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_1777 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11987__B1 net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11727_ net182 net628 vssd1 vssd1 vccd1 vccd1 _06222_ sky130_fd_sc_hd__and2_1
XFILLER_0_72_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_25_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11658_ net581 net423 _06186_ net301 net1441 vssd1 vssd1 vccd1 vccd1 _00461_ sky130_fd_sc_hd__a32o_1
XFILLER_0_71_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11739__A0 net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10609_ _05351_ _05352_ vssd1 vssd1 vccd1 vccd1 _05353_ sky130_fd_sc_hd__nor2_1
XANTENNA__09197__Y _04116_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07407__A1 final_design.data_from_mem\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09638__B net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11589_ net577 net423 _06150_ net304 net2493 vssd1 vssd1 vccd1 vccd1 _00428_ sky130_fd_sc_hd__a32o_1
XFILLER_0_3_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold907 final_design.cpu.reg_window\[505\] vssd1 vssd1 vccd1 vccd1 net2249 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold918 final_design.cpu.reg_window\[824\] vssd1 vssd1 vccd1 vccd1 net2260 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10411__B1 net1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13328_ clknet_leaf_33_clk _00559_ net1238 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[316\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold929 final_design.cpu.reg_window\[599\] vssd1 vssd1 vccd1 vccd1 net2271 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13259_ clknet_leaf_53_clk _00490_ net1187 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[247\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_1873 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07873__S net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07820_ _02734_ _02736_ _02766_ _02767_ vssd1 vssd1 vccd1 vccd1 _02771_ sky130_fd_sc_hd__o22a_1
XANTENNA__11248__X _05951_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09373__B _04046_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07174__A net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07751_ _01626_ _02700_ vssd1 vssd1 vccd1 vccd1 _02702_ sky130_fd_sc_hd__or2_2
XANTENNA__13726__CLK clknet_leaf_11_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06702_ final_design.cpu.reg_window\[601\] final_design.cpu.reg_window\[633\] net930
+ vssd1 vssd1 vccd1 vccd1 _01653_ sky130_fd_sc_hd__mux2_1
XANTENNA__07569__S1 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09660__Y _04579_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07682_ _02629_ _02630_ _02631_ _02632_ net684 net693 vssd1 vssd1 vccd1 vccd1 _02633_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_71_1508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09421_ net497 _04112_ vssd1 vssd1 vccd1 vccd1 _04340_ sky130_fd_sc_hd__nor2_1
X_06633_ final_design.cpu.reg_window\[859\] final_design.cpu.reg_window\[891\] net943
+ vssd1 vssd1 vccd1 vccd1 _01584_ sky130_fd_sc_hd__mux2_1
XANTENNA__08717__B _01690_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09352_ _02673_ net445 net442 _02670_ _04270_ vssd1 vssd1 vccd1 vccd1 _04271_ sky130_fd_sc_hd__o221a_1
XANTENNA__13876__CLK clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08677__A_N net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06564_ _01511_ _01512_ _01513_ _01514_ net777 net794 vssd1 vssd1 vccd1 vccd1 _01515_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__09096__B1 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08303_ final_design.cpu.reg_window\[905\] final_design.cpu.reg_window\[937\] net810
+ vssd1 vssd1 vccd1 vccd1 _03254_ sky130_fd_sc_hd__mux2_1
XANTENNA__11978__B1 net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09283_ _04200_ _04201_ net478 vssd1 vssd1 vccd1 vccd1 _04202_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_79_2902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_1404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06495_ final_design.cpu.reg_window\[734\] final_design.cpu.reg_window\[766\] net933
+ vssd1 vssd1 vccd1 vccd1 _01446_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_79_2913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout235_A _05982_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08234_ _03181_ _03182_ _03183_ _03184_ net678 net698 vssd1 vssd1 vccd1 vccd1 _03185_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_51_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_991 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_30_clk_A clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13106__CLK clknet_leaf_39_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08165_ net716 _03115_ vssd1 vssd1 vccd1 vccd1 _03116_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout402_A _06257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1144_A net1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07116_ _02065_ _02066_ vssd1 vssd1 vccd1 vccd1 _02067_ sky130_fd_sc_hd__nand2_1
XFILLER_0_82_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08096_ final_design.cpu.reg_window\[76\] final_design.cpu.reg_window\[108\] net814
+ vssd1 vssd1 vccd1 vccd1 _03047_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_45_clk_A clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13256__CLK clknet_leaf_41_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07047_ final_design.data_from_mem\[14\] net970 _01997_ vssd1 vssd1 vccd1 vccd1 _01998_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_60_1913 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12155__A0 net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06540__X _01491_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout771_A _01422_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout392_X net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout869_A net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08374__A2 _03321_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08998_ net623 _03932_ vssd1 vssd1 vccd1 vccd1 _03933_ sky130_fd_sc_hd__nor2_1
X_07949_ _02897_ _02899_ vssd1 vssd1 vccd1 vccd1 _02900_ sky130_fd_sc_hd__or2_2
X_10960_ net670 _05674_ _05687_ net966 _05686_ vssd1 vssd1 vccd1 vccd1 _05688_ sky130_fd_sc_hd__o221a_1
XFILLER_0_35_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09619_ _04077_ net319 vssd1 vssd1 vccd1 vccd1 _04538_ sky130_fd_sc_hd__nand2_1
X_10891_ _05621_ vssd1 vssd1 vccd1 vccd1 _05622_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout824_X net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12630_ _06302_ net1401 net980 vssd1 vssd1 vccd1 vccd1 _01317_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_14_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_1452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11969__B1 net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07023__S net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12561_ _06224_ net353 net324 net1886 vssd1 vssd1 vccd1 vccd1 _01265_ sky130_fd_sc_hd__a22o_1
XFILLER_0_19_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11512_ net1685 net216 net521 vssd1 vssd1 vccd1 vccd1 _00381_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12492_ _06152_ net355 net332 net2212 vssd1 vssd1 vccd1 vccd1 _01198_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_43_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14031__CLK clknet_leaf_42_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14231_ net1285 vssd1 vssd1 vccd1 vccd1 gpio_out[9] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_43_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11443_ net673 net638 vssd1 vssd1 vccd1 vccd1 _06094_ sky130_fd_sc_hd__and2_1
XANTENNA__09458__B net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11197__A1 net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14162_ clknet_leaf_18_clk _01336_ net1109 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.data_to_VGA\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_11374_ net436 net581 _06061_ net316 net1623 vssd1 vssd1 vccd1 vccd1 _00302_ sky130_fd_sc_hd__a32o_1
XANTENNA__13204__RESET_B net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13113_ clknet_leaf_52_clk _00344_ net1143 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[101\]
+ sky130_fd_sc_hd__dfrtp_1
X_10325_ net1544 net1009 net986 final_design.data_from_mem\[10\] vssd1 vssd1 vccd1
+ vccd1 _00082_ sky130_fd_sc_hd__a22o_1
X_14093_ clknet_leaf_14_clk _01290_ net1110 vssd1 vssd1 vccd1 vccd1 final_design.reqhand.instruction\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14181__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13044_ clknet_leaf_13_clk _00275_ net1088 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[32\]
+ sky130_fd_sc_hd__dfrtp_1
X_10256_ _05123_ net797 _05122_ vssd1 vssd1 vccd1 vccd1 _00018_ sky130_fd_sc_hd__and3b_1
XANTENNA__13749__CLK clknet_leaf_58_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09905__C _04823_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1210 net1212 vssd1 vssd1 vccd1 vccd1 net1210 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_37_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1221 net1226 vssd1 vssd1 vccd1 vccd1 net1221 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_33_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12104__S net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1232 net1235 vssd1 vssd1 vccd1 vccd1 net1232 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09193__B _03649_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10187_ _05073_ _05074_ _05075_ _05076_ vssd1 vssd1 vccd1 vccd1 _05077_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_33_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1243 net1244 vssd1 vssd1 vccd1 vccd1 net1243 sky130_fd_sc_hd__clkbuf_2
Xclkbuf_leaf_58_clk clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_58_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__09314__A1 net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08117__A2 _03065_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13899__CLK clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13946_ clknet_leaf_63_clk _01177_ net1121 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[934\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_1374 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13877_ clknet_leaf_56_clk _01108_ net1146 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[865\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11244__A net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07971__S1 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12828_ net1363 vssd1 vssd1 vccd1 vccd1 _00269_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__13129__CLK clknet_leaf_36_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1913 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12621__A1 final_design.reqhand.data_from_UART\[7\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_12759_ net954 _06382_ _06394_ _06395_ vssd1 vssd1 vccd1 vccd1 _01353_ sky130_fd_sc_hd__a31o_1
XFILLER_0_45_928 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10294__S net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13279__CLK clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold704 final_design.cpu.reg_window\[400\] vssd1 vssd1 vccd1 vccd1 net2046 sky130_fd_sc_hd__dlygate4sd3_1
Xhold715 final_design.cpu.reg_window\[794\] vssd1 vssd1 vccd1 vccd1 net2057 sky130_fd_sc_hd__dlygate4sd3_1
Xhold726 final_design.cpu.reg_window\[442\] vssd1 vssd1 vccd1 vccd1 net2068 sky130_fd_sc_hd__dlygate4sd3_1
Xhold737 final_design.cpu.reg_window\[438\] vssd1 vssd1 vccd1 vccd1 net2079 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold748 final_design.cpu.reg_window\[729\] vssd1 vssd1 vccd1 vccd1 net2090 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07800__A1 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09970_ _03327_ net446 _04119_ _04066_ _04888_ vssd1 vssd1 vccd1 vccd1 _04889_ sky130_fd_sc_hd__o221a_1
XFILLER_0_60_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold759 final_design.cpu.reg_window\[321\] vssd1 vssd1 vccd1 vccd1 net2101 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08921_ _03757_ _03863_ vssd1 vssd1 vccd1 vccd1 _03864_ sky130_fd_sc_hd__xor2_1
XFILLER_0_21_880 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12998__RESET_B net1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08852_ final_design.CPU_instr_adr\[31\] _03802_ vssd1 vssd1 vccd1 vccd1 _03803_
+ sky130_fd_sc_hd__xor2_1
XANTENNA__07175__Y _02126_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1717 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11360__A1 final_design.data_from_mem\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07803_ final_design.cpu.reg_window\[985\] final_design.cpu.reg_window\[1017\] net853
+ vssd1 vssd1 vccd1 vccd1 _02754_ sky130_fd_sc_hd__mux2_1
X_08783_ _03688_ _03732_ _03687_ vssd1 vssd1 vccd1 vccd1 _03734_ sky130_fd_sc_hd__and3b_1
Xclkbuf_leaf_49_clk clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_49_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout185_A _06060_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07734_ net719 _02684_ vssd1 vssd1 vccd1 vccd1 _02685_ sky130_fd_sc_hd__or2_1
XFILLER_0_27_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07632__A net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07665_ _02612_ _02613_ _02614_ _02615_ net684 net703 vssd1 vssd1 vccd1 vccd1 _02616_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout352_A net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1094_A net1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09404_ _02606_ _04171_ _02576_ vssd1 vssd1 vccd1 vccd1 _04323_ sky130_fd_sc_hd__a21o_1
X_06616_ net885 _01559_ _01565_ _01547_ _01553_ vssd1 vssd1 vccd1 vccd1 _01567_ sky130_fd_sc_hd__a32o_2
XANTENNA__09069__B1 net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07596_ final_design.cpu.reg_window\[477\] final_design.cpu.reg_window\[509\] net870
+ vssd1 vssd1 vccd1 vccd1 _02547_ sky130_fd_sc_hd__mux2_1
XANTENNA__14054__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09335_ _02704_ _04049_ vssd1 vssd1 vccd1 vccd1 _04254_ sky130_fd_sc_hd__nor2_1
X_06547_ _01484_ _01488_ net734 _01494_ vssd1 vssd1 vccd1 vccd1 _01498_ sky130_fd_sc_hd__or4_4
XANTENNA_fanout617_A net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09266_ net72 _04184_ vssd1 vssd1 vccd1 vccd1 _04185_ sky130_fd_sc_hd__or2_2
X_06478_ final_design.cpu.reg_window\[414\] final_design.cpu.reg_window\[446\] net931
+ vssd1 vssd1 vccd1 vccd1 _01429_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08217_ _02097_ net598 vssd1 vssd1 vccd1 vccd1 _03168_ sky130_fd_sc_hd__nand2_1
X_09197_ net497 _04055_ vssd1 vssd1 vccd1 vccd1 _04116_ sky130_fd_sc_hd__nor2_2
XANTENNA_fanout405_X net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08148_ net600 _03096_ _03072_ net540 vssd1 vssd1 vccd1 vccd1 _03099_ sky130_fd_sc_hd__o211a_1
XANTENNA__08044__A1 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout986_A _05167_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09792__A1 net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08079_ _02994_ _02995_ _03025_ _03027_ vssd1 vssd1 vccd1 vccd1 _03030_ sky130_fd_sc_hd__o22a_1
X_10110_ final_design.VGA_data_control.v_count\[2\] final_design.VGA_data_control.v_count\[3\]
+ _05019_ vssd1 vssd1 vccd1 vccd1 _05023_ sky130_fd_sc_hd__and3_1
X_11090_ net963 _05811_ vssd1 vssd1 vccd1 vccd1 _05812_ sky130_fd_sc_hd__nand2_1
XANTENNA__12679__B2 final_design.data_from_mem\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06711__A _01658_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout774_X net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10041_ _04479_ _04532_ _04552_ _04959_ vssd1 vssd1 vccd1 vccd1 _04960_ sky130_fd_sc_hd__and4_1
Xhold20 net131 vssd1 vssd1 vccd1 vccd1 net1362 sky130_fd_sc_hd__dlygate4sd3_1
Xhold31 net104 vssd1 vssd1 vccd1 vccd1 net1373 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold42 net162 vssd1 vssd1 vccd1 vccd1 net1384 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_51_1950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold53 final_design.cpu.reg_window\[28\] vssd1 vssd1 vccd1 vccd1 net1395 sky130_fd_sc_hd__dlygate4sd3_1
Xhold64 final_design.VGA_data_control.data_to_VGA\[11\] vssd1 vssd1 vccd1 vccd1 net1406
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_1238 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold75 final_design.cpu.reg_window\[711\] vssd1 vssd1 vccd1 vccd1 net1417 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11763__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold86 final_design.VGA_data_control.data_to_VGA\[30\] vssd1 vssd1 vccd1 vccd1 net1428
+ sky130_fd_sc_hd__dlygate4sd3_1
X_13800_ clknet_leaf_41_clk _01031_ net1225 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[788\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold97 final_design.VGA_data_control.data_to_VGA\[6\] vssd1 vssd1 vccd1 vccd1 net1439
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_1601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11992_ _06195_ net282 net401 net2108 vssd1 vssd1 vccd1 vccd1 _00724_ sky130_fd_sc_hd__a22o_1
X_10943_ _05604_ _05668_ _05669_ _05670_ vssd1 vssd1 vccd1 vccd1 _05671_ sky130_fd_sc_hd__o211ai_1
X_13731_ clknet_leaf_0_clk _00962_ net1062 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[719\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11654__A2 net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07261__B _01598_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10874_ _05602_ _05605_ vssd1 vssd1 vccd1 vccd1 _05606_ sky130_fd_sc_hd__or2_1
Xclkbuf_3_0_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_3_0_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_42_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13662_ clknet_leaf_11_clk _00893_ net1087 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[650\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_71_1861 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_1356 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12613_ net2182 net998 net984 final_design.data_from_mem\[31\] vssd1 vssd1 vccd1
+ vccd1 _01306_ sky130_fd_sc_hd__a22o_1
X_13593_ clknet_leaf_52_clk _00824_ net1170 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[581\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_45_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12603__B2 final_design.data_from_mem\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13421__CLK clknet_leaf_44_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10614__B1 net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12544_ _06207_ net353 net324 net2053 vssd1 vssd1 vccd1 vccd1 _01248_ sky130_fd_sc_hd__a22o_1
XANTENNA__06592__S net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12891__Q final_design.data_from_mem\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_20_Left_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12475_ _06135_ net344 net330 net1938 vssd1 vssd1 vccd1 vccd1 _01181_ sky130_fd_sc_hd__a22o_1
X_14214_ net1272 vssd1 vssd1 vccd1 vccd1 gpio_oeb[26] sky130_fd_sc_hd__buf_2
X_11426_ net1589 net223 net313 vssd1 vssd1 vccd1 vccd1 _00323_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_1643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_6 _05934_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13571__CLK clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14145_ clknet_leaf_18_clk _01319_ net1114 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.data_to_VGA\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_39_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11357_ net583 net424 _06046_ net316 net1599 vssd1 vssd1 vccd1 vccd1 _00300_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_39_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10393__A2 net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10308_ _05147_ _05159_ _05161_ final_design.VGA_data_control.h_count\[5\] vssd1
+ vssd1 vccd1 vccd1 _05162_ sky130_fd_sc_hd__a31o_1
X_14076_ clknet_leaf_15_clk _01273_ net1095 vssd1 vssd1 vccd1 vccd1 final_design.uart.working_data\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_11288_ net738 _03918_ vssd1 vssd1 vccd1 vccd1 _05986_ sky130_fd_sc_hd__nand2_1
X_13027_ clknet_leaf_0_clk _00258_ net1062 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08338__A2 _03287_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10239_ final_design.uart.BAUD_counter\[13\] final_design.uart.BAUD_counter\[14\]
+ _05109_ vssd1 vssd1 vccd1 vccd1 _05113_ sky130_fd_sc_hd__and3_1
XFILLER_0_20_1226 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11342__A1 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1040 _01394_ vssd1 vssd1 vccd1 vccd1 net1040 sky130_fd_sc_hd__clkbuf_2
Xfanout1051 final_design.VGA_data_control.v_count\[4\] vssd1 vssd1 vccd1 vccd1 net1051
+ sky130_fd_sc_hd__clkbuf_2
Xfanout1062 net1069 vssd1 vssd1 vccd1 vccd1 net1062 sky130_fd_sc_hd__clkbuf_4
Xfanout1073 net1076 vssd1 vssd1 vccd1 vccd1 net1073 sky130_fd_sc_hd__clkbuf_4
Xfanout1084 net1085 vssd1 vssd1 vccd1 vccd1 net1084 sky130_fd_sc_hd__buf_2
Xfanout1095 net1096 vssd1 vssd1 vccd1 vccd1 net1095 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08548__A net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09838__A2 _04435_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14077__CLK clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13929_ clknet_leaf_37_clk _01160_ net1228 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[917\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_18_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07450_ final_design.cpu.reg_window\[64\] final_design.cpu.reg_window\[96\] net895
+ vssd1 vssd1 vccd1 vccd1 _02401_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_1901 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07381_ _02325_ _02330_ vssd1 vssd1 vccd1 vccd1 _02332_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_2_1721 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09120_ net961 _04037_ vssd1 vssd1 vccd1 vccd1 _04039_ sky130_fd_sc_hd__nand2_1
XFILLER_0_17_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07598__S net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_2290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07077__A2 net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12070__A2 net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13914__CLK clknet_leaf_63_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09051_ net622 _03979_ _03977_ net254 vssd1 vssd1 vccd1 vccd1 _03980_ sky130_fd_sc_hd__a211o_1
XPHY_EDGE_ROW_6_Right_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08002_ final_design.cpu.reg_window\[912\] final_design.cpu.reg_window\[944\] net843
+ vssd1 vssd1 vccd1 vccd1 _02953_ sky130_fd_sc_hd__mux2_1
XANTENNA__12358__B1 net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold501 final_design.cpu.reg_window\[468\] vssd1 vssd1 vccd1 vccd1 net1843 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10908__A1 net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10908__B2 net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold512 final_design.cpu.reg_window\[698\] vssd1 vssd1 vccd1 vccd1 net1854 sky130_fd_sc_hd__dlygate4sd3_1
Xhold523 final_design.cpu.reg_window\[131\] vssd1 vssd1 vccd1 vccd1 net1865 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09774__A1 net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold534 final_design.cpu.reg_window\[915\] vssd1 vssd1 vccd1 vccd1 net1876 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09826__B _04744_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold545 final_design.cpu.reg_window\[172\] vssd1 vssd1 vccd1 vccd1 net1887 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold556 final_design.cpu.reg_window\[471\] vssd1 vssd1 vccd1 vccd1 net1898 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11581__A1 net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold567 final_design.cpu.reg_window\[408\] vssd1 vssd1 vccd1 vccd1 net1909 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold578 final_design.cpu.reg_window\[499\] vssd1 vssd1 vccd1 vccd1 net1920 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_55_2072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold589 final_design.cpu.reg_window\[998\] vssd1 vssd1 vccd1 vccd1 net1931 sky130_fd_sc_hd__dlygate4sd3_1
X_09953_ _03487_ net441 vssd1 vssd1 vccd1 vccd1 _04872_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_55_2083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_2094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09526__A1 _04342_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11149__A net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08904_ _01661_ _01662_ _02469_ vssd1 vssd1 vccd1 vccd1 _03849_ sky130_fd_sc_hd__o21ai_1
X_09884_ _04789_ _04791_ _04792_ _04802_ vssd1 vssd1 vccd1 vccd1 _04803_ sky130_fd_sc_hd__and4bb_1
XANTENNA_fanout1107_A net1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11333__B2 net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1201 final_design.CPU_instr_adr\[30\] vssd1 vssd1 vccd1 vccd1 net2543 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1212 final_design.cpu.reg_window\[363\] vssd1 vssd1 vccd1 vccd1 net2554 sky130_fd_sc_hd__dlygate4sd3_1
X_08835_ final_design.CPU_instr_adr\[7\] final_design.CPU_instr_adr\[6\] _03785_ vssd1
+ vssd1 vccd1 vccd1 _03786_ sky130_fd_sc_hd__and3_1
XANTENNA__10988__A _04529_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout188_X net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout567_A net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08766_ _03714_ _03716_ vssd1 vssd1 vccd1 vccd1 _03717_ sky130_fd_sc_hd__and2b_1
XANTENNA__06677__S net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09829__A2 _04744_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_0_220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07717_ net877 _02649_ _02655_ _02661_ _02667_ vssd1 vssd1 vccd1 vccd1 _02668_ sky130_fd_sc_hd__o32a_2
XANTENNA__11155__Y _05869_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08697_ _02028_ _02062_ _01998_ vssd1 vssd1 vccd1 vccd1 _03648_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout355_X net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout734_A net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13444__CLK clknet_leaf_54_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_11_Left_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07935__S1 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07648_ final_design.cpu.reg_window\[540\] final_design.cpu.reg_window\[572\] net867
+ vssd1 vssd1 vccd1 vccd1 _02599_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout901_A net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07579_ final_design.cpu.reg_window\[735\] final_design.cpu.reg_window\[767\] net857
+ vssd1 vssd1 vccd1 vccd1 _02530_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout522_X net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08464__Y _03415_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09318_ _02389_ net456 vssd1 vssd1 vccd1 vccd1 _04237_ sky130_fd_sc_hd__nand2_1
X_10590_ _05311_ _05333_ vssd1 vssd1 vccd1 vccd1 _05335_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_1_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07301__S net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09249_ _02735_ _02768_ _02766_ vssd1 vssd1 vccd1 vccd1 _04168_ sky130_fd_sc_hd__a21o_1
XANTENNA__12349__B1 net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12260_ net586 _06189_ net513 net374 net1643 vssd1 vssd1 vccd1 vccd1 _00976_ sky130_fd_sc_hd__a32o_1
XFILLER_0_27_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11758__S net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11211_ final_design.data_from_mem\[8\] _05914_ _05917_ vssd1 vssd1 vccd1 vccd1 _05918_
+ sky130_fd_sc_hd__a21o_1
XANTENNA__08112__S1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12191_ net2329 net184 net382 vssd1 vssd1 vccd1 vccd1 _00910_ sky130_fd_sc_hd__mux2_1
XANTENNA__10375__A2 net1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07537__A net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11142_ _05855_ _05856_ _05852_ vssd1 vssd1 vccd1 vccd1 _05857_ sky130_fd_sc_hd__a21o_1
XANTENNA__07871__S0 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11073_ _05172_ _05795_ vssd1 vssd1 vccd1 vccd1 _05796_ sky130_fd_sc_hd__nor2_1
XANTENNA__12521__B1 net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input30_A DAT_I[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09752__A _04072_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10024_ _02835_ net442 net439 _02834_ vssd1 vssd1 vccd1 vccd1 _04943_ sky130_fd_sc_hd__o22a_1
XANTENNA__11493__S net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12886__Q final_design.data_from_mem\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10410__B _05181_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11975_ _06177_ net285 net406 net1848 vssd1 vssd1 vccd1 vccd1 _00708_ sky130_fd_sc_hd__a22o_1
XFILLER_0_19_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_1827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13714_ clknet_leaf_38_clk _00945_ net1189 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[702\]
+ sky130_fd_sc_hd__dfrtp_1
X_10926_ _05632_ _05634_ _05652_ _05653_ vssd1 vssd1 vccd1 vccd1 _05655_ sky130_fd_sc_hd__o211a_1
XFILLER_0_67_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13937__CLK clknet_leaf_34_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10857_ net80 net1044 vssd1 vssd1 vccd1 vccd1 _05589_ sky130_fd_sc_hd__nor2_1
X_13645_ clknet_leaf_48_clk _00876_ net1185 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[633\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12588__B1 net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10788_ _05522_ _05523_ vssd1 vssd1 vccd1 vccd1 _05524_ sky130_fd_sc_hd__or2_1
X_13576_ clknet_leaf_35_clk _00807_ net1219 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[564\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_1705 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10451__A1_N net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_59_Right_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11260__B1 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08351__S1 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12527_ _06189_ net358 net328 net2327 vssd1 vssd1 vccd1 vccd1 _01232_ sky130_fd_sc_hd__a22o_1
XFILLER_0_67_1749 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12458_ net2098 net186 net337 vssd1 vssd1 vccd1 vccd1 _01165_ sky130_fd_sc_hd__mux2_1
XANTENNA__12624__Y _06299_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11409_ net673 net429 _06091_ vssd1 vssd1 vccd1 vccd1 _06092_ sky130_fd_sc_hd__and3_4
XFILLER_0_1_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12389_ net1591 net188 net270 vssd1 vssd1 vccd1 vccd1 _01100_ sky130_fd_sc_hd__mux2_1
XANTENNA__10366__A2 net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11563__A1 net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14128_ clknet_leaf_20_clk final_design.vga.v_next_count\[8\] net1158 vssd1 vssd1
+ vccd1 vccd1 final_design.VGA_data_control.v_count\[8\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__13317__CLK clknet_leaf_49_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06950_ _01897_ _01898_ _01899_ _01900_ net773 net791 vssd1 vssd1 vccd1 vccd1 _01901_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_78_1801 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14059_ clknet_leaf_16_clk _00021_ net1092 vssd1 vssd1 vccd1 vccd1 final_design.uart.BAUD_counter\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_68_Right_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12512__B1 net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1845 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06881_ final_design.cpu.reg_window\[83\] final_design.cpu.reg_window\[115\] net912
+ vssd1 vssd1 vccd1 vccd1 _01832_ sky130_fd_sc_hd__mux2_1
XANTENNA__11866__A2 net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13467__CLK clknet_leaf_65_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08620_ _02127_ _03226_ vssd1 vssd1 vccd1 vccd1 _03571_ sky130_fd_sc_hd__and2_1
XFILLER_0_74_1709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1889 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06497__S net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08551_ final_design.cpu.reg_window\[769\] final_design.cpu.reg_window\[801\] net838
+ vssd1 vssd1 vccd1 vccd1 _03502_ sky130_fd_sc_hd__mux2_1
XANTENNA__11618__A2 net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07502_ _01970_ _02001_ _01969_ vssd1 vssd1 vccd1 vccd1 _02453_ sky130_fd_sc_hd__a21o_1
X_08482_ final_design.cpu.reg_window\[3\] final_design.cpu.reg_window\[35\] net820
+ vssd1 vssd1 vccd1 vccd1 _03433_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_63_2352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_2363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07433_ final_design.cpu.reg_window\[641\] final_design.cpu.reg_window\[673\] net914
+ vssd1 vssd1 vccd1 vccd1 _02384_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_82_2997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08590__S1 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_2374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1851 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_77_Right_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07364_ final_design.cpu.reg_window\[963\] final_design.cpu.reg_window\[995\] net904
+ vssd1 vssd1 vccd1 vccd1 _02315_ sky130_fd_sc_hd__mux2_1
X_09103_ _03713_ _03718_ vssd1 vssd1 vccd1 vccd1 _04025_ sky130_fd_sc_hd__xor2_1
XANTENNA__10054__A1 net68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11151__B net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09995__A1 net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07295_ final_design.cpu.reg_window\[133\] final_design.cpu.reg_window\[165\] net921
+ vssd1 vssd1 vccd1 vccd1 _02246_ sky130_fd_sc_hd__mux2_1
XANTENNA__09995__B2 net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout315_A _05851_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1057_A final_design.reqhand.current_client\[3\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09034_ _03789_ _03964_ vssd1 vssd1 vccd1 vccd1 _03965_ sky130_fd_sc_hd__nor2_1
XFILLER_0_14_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_2145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_2156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12942__RESET_B net1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold320 final_design.reqhand.instruction\[14\] vssd1 vssd1 vccd1 vccd1 net1662 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_2167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold331 final_design.cpu.reg_window\[792\] vssd1 vssd1 vccd1 vccd1 net1673 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_53_2009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12263__A net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10357__A2 net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold342 final_design.cpu.reg_window\[241\] vssd1 vssd1 vccd1 vccd1 net1684 sky130_fd_sc_hd__dlygate4sd3_1
Xhold353 final_design.cpu.reg_window\[83\] vssd1 vssd1 vccd1 vccd1 net1695 sky130_fd_sc_hd__dlygate4sd3_1
Xhold364 final_design.cpu.reg_window\[852\] vssd1 vssd1 vccd1 vccd1 net1706 sky130_fd_sc_hd__dlygate4sd3_1
Xhold375 final_design.cpu.reg_window\[461\] vssd1 vssd1 vccd1 vccd1 net1717 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout800 _05090_ vssd1 vssd1 vccd1 vccd1 net800 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_fanout684_A net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold386 final_design.cpu.reg_window\[526\] vssd1 vssd1 vccd1 vccd1 net1728 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_91 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout811 net829 vssd1 vssd1 vccd1 vccd1 net811 sky130_fd_sc_hd__clkbuf_4
Xhold397 final_design.cpu.reg_window\[650\] vssd1 vssd1 vccd1 vccd1 net1739 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08970__A2 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout822 net823 vssd1 vssd1 vccd1 vccd1 net822 sky130_fd_sc_hd__clkbuf_2
X_09936_ _03391_ net446 net441 _03389_ vssd1 vssd1 vccd1 vccd1 _04855_ sky130_fd_sc_hd__o22a_1
Xfanout833 net834 vssd1 vssd1 vccd1 vccd1 net833 sky130_fd_sc_hd__buf_2
XANTENNA__11306__A1 net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout844 net847 vssd1 vssd1 vccd1 vccd1 net844 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_1855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12503__B1 net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout855 net872 vssd1 vssd1 vccd1 vccd1 net855 sky130_fd_sc_hd__clkbuf_4
Xfanout866 net867 vssd1 vssd1 vccd1 vccd1 net866 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07605__S0 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11857__A2 net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09867_ _04125_ _04785_ _04784_ _04777_ vssd1 vssd1 vccd1 vccd1 _04786_ sky130_fd_sc_hd__a211o_1
Xfanout877 net878 vssd1 vssd1 vccd1 vccd1 net877 sky130_fd_sc_hd__buf_4
Xhold1020 final_design.cpu.reg_window\[315\] vssd1 vssd1 vccd1 vccd1 net2362 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout888 net890 vssd1 vssd1 vccd1 vccd1 net888 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_5_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1031 final_design.cpu.reg_window\[809\] vssd1 vssd1 vccd1 vccd1 net2373 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout899 net910 vssd1 vssd1 vccd1 vccd1 net899 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout949_A net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1042 final_design.cpu.reg_window\[613\] vssd1 vssd1 vccd1 vccd1 net2384 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11607__A net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08818_ final_design.CPU_instr_adr\[24\] _01691_ vssd1 vssd1 vccd1 vccd1 _03769_
+ sky130_fd_sc_hd__nor2_1
Xhold1053 final_design.cpu.reg_window\[638\] vssd1 vssd1 vccd1 vccd1 net2395 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10511__A net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1064 final_design.cpu.reg_window\[626\] vssd1 vssd1 vccd1 vccd1 net2406 sky130_fd_sc_hd__dlygate4sd3_1
X_09798_ _04072_ _04714_ _04716_ vssd1 vssd1 vccd1 vccd1 _04717_ sky130_fd_sc_hd__or3b_1
Xhold1075 final_design.cpu.reg_window\[807\] vssd1 vssd1 vccd1 vccd1 net2417 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12834__CLK clknet_leaf_19_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1086 final_design.cpu.reg_window\[672\] vssd1 vssd1 vccd1 vccd1 net2428 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1097 final_design.cpu.reg_window\[541\] vssd1 vssd1 vccd1 vccd1 net2439 sky130_fd_sc_hd__dlygate4sd3_1
X_08749_ final_design.CPU_instr_adr\[6\] _02240_ vssd1 vssd1 vccd1 vccd1 _03700_ sky130_fd_sc_hd__nand2_1
XFILLER_0_68_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_1090 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11760_ net191 net2192 net419 vssd1 vssd1 vccd1 vccd1 _00523_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09683__B1 net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10711_ _05425_ _05429_ _05427_ vssd1 vssd1 vccd1 vccd1 _05450_ sky130_fd_sc_hd__o21ai_1
X_11691_ net216 net626 vssd1 vssd1 vccd1 vccd1 _06204_ sky130_fd_sc_hd__and2_1
XFILLER_0_49_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10642_ _05364_ _05383_ vssd1 vssd1 vccd1 vccd1 _05385_ sky130_fd_sc_hd__and2_2
X_13430_ clknet_leaf_60_clk _00661_ net1138 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[418\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_48_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1214 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10045__B2 _04423_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13361_ clknet_leaf_35_clk _00592_ net1241 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[349\]
+ sky130_fd_sc_hd__dfrtp_1
X_10573_ _05317_ _05318_ vssd1 vssd1 vccd1 vccd1 _05319_ sky130_fd_sc_hd__and2_1
XFILLER_0_1_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_739 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10596__A2 net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12312_ net1592 net206 net364 vssd1 vssd1 vccd1 vccd1 _01026_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13292_ clknet_leaf_46_clk _00523_ net1216 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[280\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input78_A memory_size[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08651__A _01627_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_20_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09738__A1 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12243_ net578 _06173_ net510 net374 net1594 vssd1 vssd1 vccd1 vccd1 _00960_ sky130_fd_sc_hd__a32o_1
XANTENNA__11545__A1 net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12174_ net1739 net217 net380 vssd1 vssd1 vccd1 vccd1 _00893_ sky130_fd_sc_hd__mux2_1
XANTENNA__07844__S0 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11125_ net804 _05839_ vssd1 vssd1 vccd1 vccd1 _05840_ sky130_fd_sc_hd__and2_2
XFILLER_0_60_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11056_ net88 net1045 net89 vssd1 vssd1 vccd1 vccd1 _05779_ sky130_fd_sc_hd__or3b_1
XANTENNA__11848__A2 net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10007_ _03640_ net438 vssd1 vssd1 vccd1 vccd1 _04926_ sky130_fd_sc_hd__nor2_1
XFILLER_0_64_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12112__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10421__A _03192_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11236__B net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11958_ net1933 net404 _06256_ net230 vssd1 vssd1 vccd1 vccd1 _00691_ sky130_fd_sc_hd__a22o_1
XANTENNA__09674__B1 net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06488__B1 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10909_ final_design.CPU_instr_adr\[22\] net1000 vssd1 vssd1 vccd1 vccd1 _05639_
+ sky130_fd_sc_hd__nor2_1
X_11889_ net239 net2120 net273 vssd1 vssd1 vccd1 vccd1 _00631_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14115__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08229__A1 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13628_ clknet_leaf_2_clk _00859_ net1068 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[616\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09426__B1 net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11233__B1 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13559_ clknet_leaf_4_clk _00790_ net1083 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[547\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07876__S net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07080_ _02030_ vssd1 vssd1 vccd1 vccd1 _02031_ sky130_fd_sc_hd__inv_2
XFILLER_0_70_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08561__A net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_71_2621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_71_2632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_2643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07982_ net613 _02929_ _02931_ net545 vssd1 vssd1 vccd1 vccd1 _02933_ sky130_fd_sc_hd__a211oi_2
XANTENNA__12857__CLK clknet_leaf_17_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09721_ _03069_ net444 vssd1 vssd1 vccd1 vccd1 _04640_ sky130_fd_sc_hd__or2_1
X_06933_ _01883_ vssd1 vssd1 vccd1 vccd1 _01884_ sky130_fd_sc_hd__inv_2
XFILLER_0_38_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_1631 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06864_ net885 _01796_ _01802_ _01808_ _01814_ vssd1 vssd1 vccd1 vccd1 _01815_ sky130_fd_sc_hd__o32a_4
X_09652_ net448 _04569_ _04566_ net729 vssd1 vssd1 vccd1 vccd1 _04571_ sky130_fd_sc_hd__o211ai_4
XTAP_TAPCELL_ROW_69_2550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08260__S0 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_2561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_2572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_2414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08603_ net596 _03550_ _03524_ _02419_ vssd1 vssd1 vccd1 vccd1 _03554_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_78_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_65_2425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09583_ net321 _04500_ _04501_ _04494_ vssd1 vssd1 vccd1 vccd1 _04502_ sky130_fd_sc_hd__o31ai_4
XFILLER_0_78_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06795_ final_design.cpu.reg_window\[982\] final_design.cpu.reg_window\[1014\] net919
+ vssd1 vssd1 vccd1 vccd1 _01746_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_65_2436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout265_A net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08534_ net609 _03481_ _03482_ vssd1 vssd1 vccd1 vccd1 _03485_ sky130_fd_sc_hd__a21o_2
XFILLER_0_49_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08465_ _02297_ net596 vssd1 vssd1 vccd1 vccd1 _03416_ sky130_fd_sc_hd__and2_1
XFILLER_0_65_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout432_A _05847_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07140__B2 net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07416_ final_design.cpu.reg_window\[449\] final_design.cpu.reg_window\[481\] net914
+ vssd1 vssd1 vccd1 vccd1 _02367_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09417__A0 _01535_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08396_ final_design.cpu.reg_window\[646\] final_design.cpu.reg_window\[678\] net821
+ vssd1 vssd1 vccd1 vccd1 _03347_ sky130_fd_sc_hd__mux2_1
XANTENNA__12016__A2 net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11224__B1 net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07347_ _02294_ _02297_ vssd1 vssd1 vccd1 vccd1 _02298_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_59_2207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout220_X net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_2218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_59_2229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout318_X net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11775__B2 net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06690__S net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07278_ final_design.cpu.reg_window\[774\] final_design.cpu.reg_window\[806\] net912
+ vssd1 vssd1 vccd1 vccd1 _02229_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09017_ _03790_ _03949_ vssd1 vssd1 vccd1 vccd1 _03950_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout899_A net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1227_X net1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13632__CLK clknet_leaf_11_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold150 final_design.cpu.reg_window\[201\] vssd1 vssd1 vccd1 vccd1 net1492 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09854__X _04773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09196__A2 net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold161 final_design.VGA_data_control.ready_data\[23\] vssd1 vssd1 vccd1 vccd1 net1503
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold172 final_design.VGA_data_control.ready_data\[12\] vssd1 vssd1 vccd1 vccd1 net1514
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout687_X net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold183 final_design.cpu.reg_window\[205\] vssd1 vssd1 vccd1 vccd1 net1525 sky130_fd_sc_hd__dlygate4sd3_1
Xhold194 final_design.cpu.reg_window\[722\] vssd1 vssd1 vccd1 vccd1 net1536 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout630 net631 vssd1 vssd1 vccd1 vccd1 net630 sky130_fd_sc_hd__clkbuf_4
Xfanout641 _05946_ vssd1 vssd1 vccd1 vccd1 net641 sky130_fd_sc_hd__clkbuf_4
X_09919_ net486 _04646_ _04224_ vssd1 vssd1 vccd1 vccd1 _04838_ sky130_fd_sc_hd__a21o_1
Xfanout652 _05143_ vssd1 vssd1 vccd1 vccd1 net652 sky130_fd_sc_hd__buf_4
Xfanout663 _02511_ vssd1 vssd1 vccd1 vccd1 net663 sky130_fd_sc_hd__buf_4
XANTENNA__13782__CLK clknet_leaf_58_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08410__S net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout854_X net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout674 net676 vssd1 vssd1 vccd1 vccd1 net674 sky130_fd_sc_hd__buf_4
Xfanout685 net689 vssd1 vssd1 vccd1 vccd1 net685 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_1696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12930_ clknet_leaf_47_clk _00168_ net1199 vssd1 vssd1 vccd1 vccd1 net153 sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_3_1_0_clk_X clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout696 net698 vssd1 vssd1 vccd1 vccd1 net696 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_77_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06706__A1 net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12861_ clknet_leaf_17_clk _00099_ net1108 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.ready_data\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14138__CLK clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11812_ net229 net2101 net265 vssd1 vssd1 vccd1 vccd1 _00564_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08003__S0 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07550__A net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08554__S1 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11743_ net244 net2076 net416 vssd1 vssd1 vccd1 vccd1 _00506_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12007__A2 net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13162__CLK clknet_leaf_61_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11674_ net428 net566 _06195_ net295 net1666 vssd1 vssd1 vccd1 vccd1 _00468_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_12_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13413_ clknet_leaf_48_clk _00644_ net1182 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[401\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_12_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10625_ net99 final_design.VGA_adr\[7\] vssd1 vssd1 vccd1 vccd1 _05368_ sky130_fd_sc_hd__or2_1
XFILLER_0_68_1833 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10556_ net63 _05301_ vssd1 vssd1 vccd1 vccd1 _05303_ sky130_fd_sc_hd__xnor2_1
X_13344_ clknet_leaf_10_clk _00575_ net1101 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[332\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08631__A1 net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10487_ _05235_ _05236_ vssd1 vssd1 vccd1 vccd1 _05237_ sky130_fd_sc_hd__nand2_1
X_13275_ clknet_leaf_64_clk _00506_ net1074 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[263\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12107__S net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_1432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12226_ net584 _06154_ net512 net378 net2437 vssd1 vssd1 vccd1 vccd1 _00944_ sky130_fd_sc_hd__a32o_1
XFILLER_0_23_1416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12157_ net184 net2393 net386 vssd1 vssd1 vccd1 vccd1 _00878_ sky130_fd_sc_hd__mux2_1
XANTENNA__08934__A2 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06945__A1 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11108_ _05818_ _05828_ vssd1 vssd1 vccd1 vccd1 _05829_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_75_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12088_ net583 _06053_ net514 net394 net2014 vssd1 vssd1 vccd1 vccd1 _00813_ sky130_fd_sc_hd__a32o_1
XANTENNA__13652__RESET_B net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09344__C1 _04097_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11039_ _05761_ _05762_ _05737_ vssd1 vssd1 vccd1 vccd1 _05763_ sky130_fd_sc_hd__a21oi_2
XANTENNA__12494__A2 net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06580_ final_design.cpu.reg_window\[605\] final_design.cpu.reg_window\[637\] net946
+ vssd1 vssd1 vccd1 vccd1 _01531_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13505__CLK clknet_leaf_49_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09662__A3 _04579_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08250_ final_design.cpu.reg_window\[330\] final_design.cpu.reg_window\[362\] net825
+ vssd1 vssd1 vccd1 vccd1 _03201_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_1608 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08870__A1 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07201_ final_design.cpu.reg_window\[649\] final_design.cpu.reg_window\[681\] net888
+ vssd1 vssd1 vccd1 vccd1 _02152_ sky130_fd_sc_hd__mux2_1
X_08181_ net600 net526 _03105_ net542 vssd1 vssd1 vccd1 vccd1 _03132_ sky130_fd_sc_hd__o211a_1
XANTENNA__13655__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_2830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07132_ final_design.cpu.reg_window\[907\] final_design.cpu.reg_window\[939\] net908
+ vssd1 vssd1 vccd1 vccd1 _02083_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_1917 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_2841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_73_2705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07063_ net762 _02013_ net748 vssd1 vssd1 vccd1 vccd1 _02014_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_45_1685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07965_ _02912_ _02913_ _02914_ _02915_ net683 net702 vssd1 vssd1 vccd1 vccd1 _02916_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout382_A net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13035__CLK clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09704_ _04116_ _04310_ _04621_ net496 _04622_ vssd1 vssd1 vccd1 vccd1 _04623_ sky130_fd_sc_hd__a221oi_2
XTAP_TAPCELL_ROW_67_2509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06916_ _01863_ _01864_ _01865_ _01866_ net773 net791 vssd1 vssd1 vccd1 vccd1 _01867_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_78_1461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07036__S1 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07896_ final_design.cpu.reg_window\[215\] final_design.cpu.reg_window\[247\] net849
+ vssd1 vssd1 vccd1 vccd1 _02847_ sky130_fd_sc_hd__mux2_1
XANTENNA__12485__A2 net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_4_clk_A clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09635_ _03031_ _04430_ _02997_ vssd1 vssd1 vccd1 vccd1 _04554_ sky130_fd_sc_hd__o21ai_1
X_06847_ final_design.cpu.reg_window\[20\] final_design.cpu.reg_window\[52\] net948
+ vssd1 vssd1 vccd1 vccd1 _01798_ sky130_fd_sc_hd__mux2_1
XANTENNA__07361__A1 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout268_X net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout647_A net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06778_ final_design.cpu.reg_window\[406\] final_design.cpu.reg_window\[438\] net920
+ vssd1 vssd1 vccd1 vccd1 _01729_ sky130_fd_sc_hd__mux2_1
XANTENNA__06685__S net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09566_ net546 net545 net544 net542 net454 net464 vssd1 vssd1 vccd1 vccd1 _04485_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__13185__CLK clknet_leaf_47_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11445__A0 net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08517_ net718 _03467_ vssd1 vssd1 vccd1 vccd1 _03468_ sky130_fd_sc_hd__or2_1
XFILLER_0_66_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout435_X net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09497_ net474 _04086_ _04411_ _04415_ _04410_ vssd1 vssd1 vccd1 vccd1 _04416_ sky130_fd_sc_hd__o311a_1
XANTENNA__07113__A1 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07113__B2 _02061_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08448_ final_design.cpu.reg_window\[196\] final_design.cpu.reg_window\[228\] net821
+ vssd1 vssd1 vccd1 vccd1 _03399_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_22_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08379_ final_design.cpu.reg_window\[390\] final_design.cpu.reg_window\[422\] net823
+ vssd1 vssd1 vccd1 vccd1 _03330_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_22_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14181__RESET_B net1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06441__C_N net34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10410_ _03352_ _05181_ vssd1 vssd1 vccd1 vccd1 _05188_ sky130_fd_sc_hd__or2_1
X_11390_ net435 net584 _06075_ net316 net2539 vssd1 vssd1 vccd1 vccd1 _00304_ sky130_fd_sc_hd__a32o_1
XFILLER_0_60_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06624__A0 final_design.cpu.reg_window\[411\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10341_ net1479 net1009 net986 final_design.data_from_mem\[26\] vssd1 vssd1 vccd1
+ vccd1 _00098_ sky130_fd_sc_hd__a22o_1
XANTENNA__10420__B2 net246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1438 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13060_ clknet_leaf_54_clk _00291_ net1180 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[48\]
+ sky130_fd_sc_hd__dfrtp_1
X_10272_ _05133_ net797 _05132_ vssd1 vssd1 vccd1 vccd1 _00024_ sky130_fd_sc_hd__and3b_1
XFILLER_0_28_1872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_1774 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_76_Left_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12011_ _06213_ net280 net401 net1920 vssd1 vssd1 vccd1 vccd1 _00742_ sky130_fd_sc_hd__a22o_1
XANTENNA__11766__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1004 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11993__C net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07275__S1 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08140__S net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout460 net461 vssd1 vssd1 vccd1 vccd1 net460 sky130_fd_sc_hd__buf_2
Xfanout471 _03485_ vssd1 vssd1 vccd1 vccd1 net471 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_35_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout482 net483 vssd1 vssd1 vccd1 vccd1 net482 sky130_fd_sc_hd__buf_2
X_13962_ clknet_leaf_60_clk _01193_ net1142 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[950\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout493 _03453_ vssd1 vssd1 vccd1 vccd1 net493 sky130_fd_sc_hd__buf_2
XANTENNA__12476__A2 net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13528__CLK clknet_leaf_65_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12913_ clknet_leaf_28_clk _00151_ net1193 vssd1 vssd1 vccd1 vccd1 net135 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_31_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11684__B1 net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13893_ clknet_leaf_52_clk _01124_ net1183 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[881\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07551__Y _02502_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12228__A2 _06156_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12844_ clknet_leaf_14_clk _00082_ net1106 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.ready_data\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12894__Q final_design.data_from_mem\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1745 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13678__CLK clknet_leaf_44_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1789 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11726_ net582 net423 _06221_ net296 net1595 vssd1 vssd1 vccd1 vccd1 _00494_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_29_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06863__B1 net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11657_ net186 net633 vssd1 vssd1 vccd1 vccd1 _06186_ sky130_fd_sc_hd__and2_1
X_10608_ _05349_ _05350_ _05331_ vssd1 vssd1 vccd1 vccd1 _05352_ sky130_fd_sc_hd__a21boi_1
XANTENNA__07407__A2 net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12400__A2 net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1040 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11588_ net189 net636 vssd1 vssd1 vccd1 vccd1 _06150_ sky130_fd_sc_hd__and2_1
XFILLER_0_40_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13327_ clknet_leaf_42_clk _00558_ net1225 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[315\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold908 final_design.cpu.reg_window\[494\] vssd1 vssd1 vccd1 vccd1 net2250 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10539_ net1405 net1029 net1002 _05286_ vssd1 vssd1 vccd1 vccd1 _00177_ sky130_fd_sc_hd__a22o_1
XFILLER_0_29_1658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold919 final_design.cpu.reg_window\[916\] vssd1 vssd1 vccd1 vccd1 net2261 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13258_ clknet_leaf_60_clk _00489_ net1141 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[246\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_1885 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13058__CLK clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12209_ net560 _06137_ net503 net376 net1598 vssd1 vssd1 vccd1 vccd1 _00927_ sky130_fd_sc_hd__a32o_1
X_13189_ clknet_leaf_50_clk _00420_ net1181 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[177\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07455__A net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07750_ net615 _02698_ _02699_ _01626_ vssd1 vssd1 vccd1 vccd1 _02701_ sky130_fd_sc_hd__a211oi_1
XANTENNA__12467__A2 net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06701_ final_design.cpu.reg_window\[665\] final_design.cpu.reg_window\[697\] net930
+ vssd1 vssd1 vccd1 vccd1 _01652_ sky130_fd_sc_hd__mux2_1
X_07681_ final_design.cpu.reg_window\[542\] final_design.cpu.reg_window\[574\] net853
+ vssd1 vssd1 vccd1 vccd1 _02632_ sky130_fd_sc_hd__mux2_1
XANTENNA__07343__B2 net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11264__X _05965_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06632_ net753 _01576_ net748 vssd1 vssd1 vccd1 vccd1 _01583_ sky130_fd_sc_hd__o21a_1
X_09420_ net487 _04338_ vssd1 vssd1 vccd1 vccd1 _04339_ sky130_fd_sc_hd__nand2_1
XANTENNA__12300__S net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07190__A net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09351_ _02671_ _04094_ vssd1 vssd1 vccd1 vccd1 _04270_ sky130_fd_sc_hd__nand2_1
X_06563_ final_design.cpu.reg_window\[413\] final_design.cpu.reg_window\[445\] net950
+ vssd1 vssd1 vccd1 vccd1 _01514_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08302_ final_design.cpu.reg_window\[969\] final_design.cpu.reg_window\[1001\] net810
+ vssd1 vssd1 vccd1 vccd1 _03253_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09282_ net546 net545 net544 net542 net459 net469 vssd1 vssd1 vccd1 vccd1 _04201_
+ sky130_fd_sc_hd__mux4_1
X_06494_ net753 _01444_ vssd1 vssd1 vccd1 vccd1 _01445_ sky130_fd_sc_hd__or2_2
XFILLER_0_1_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_2903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_79_2914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08233_ final_design.cpu.reg_window\[907\] final_design.cpu.reg_window\[939\] net826
+ vssd1 vssd1 vccd1 vccd1 _03184_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08164_ _03111_ _03112_ _03113_ _03114_ net674 net696 vssd1 vssd1 vccd1 vccd1 _03115_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__09399__A2 net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08225__S net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07115_ _02058_ _02063_ vssd1 vssd1 vccd1 vccd1 _02066_ sky130_fd_sc_hd__nand2_1
XFILLER_0_31_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08095_ _03042_ _03043_ _03044_ _03045_ net675 net697 vssd1 vssd1 vccd1 vccd1 _03046_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_82_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07046_ net1041 net993 net990 final_design.reqhand.instruction\[14\] vssd1 vssd1
+ vccd1 vccd1 _01997_ sky130_fd_sc_hd__a31o_1
XFILLER_0_63_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout597_A net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07031__B1 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08997_ _03738_ _03739_ vssd1 vssd1 vccd1 vccd1 _03932_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout764_A net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout385_X net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09859__A0 net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07948_ net602 _02894_ _02869_ _01750_ vssd1 vssd1 vccd1 vccd1 _02899_ sky130_fd_sc_hd__o211a_1
XFILLER_0_78_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11666__B1 net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout931_A net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07879_ net878 _02811_ _02817_ _02823_ _02829_ vssd1 vssd1 vccd1 vccd1 _02830_ sky130_fd_sc_hd__o32a_4
XANTENNA_fanout552_X net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08467__Y _03418_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11615__A net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09618_ _04059_ net320 vssd1 vssd1 vccd1 vccd1 _04537_ sky130_fd_sc_hd__nand2_1
XANTENNA__13820__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10890_ net49 _05620_ vssd1 vssd1 vccd1 vccd1 _05621_ sky130_fd_sc_hd__xor2_1
XANTENNA__08196__A net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09549_ _04342_ _04460_ _04465_ _04467_ vssd1 vssd1 vccd1 vccd1 _04468_ sky130_fd_sc_hd__o31ai_2
XANTENNA_fanout817_X net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12560_ _06223_ net358 net324 net2357 vssd1 vssd1 vccd1 vccd1 _01264_ sky130_fd_sc_hd__a22o_1
XANTENNA__12091__B1 net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11511_ net1999 net218 net521 vssd1 vssd1 vccd1 vccd1 _00380_ sky130_fd_sc_hd__mux2_1
XANTENNA__13970__CLK clknet_leaf_39_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12491_ _06151_ net355 net332 net2166 vssd1 vssd1 vccd1 vccd1 _01197_ sky130_fd_sc_hd__a22o_1
XFILLER_0_18_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14230_ net1284 vssd1 vssd1 vccd1 vccd1 gpio_out[8] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_43_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11442_ net805 _02359_ net803 vssd1 vssd1 vccd1 vccd1 _06093_ sky130_fd_sc_hd__and3_4
XANTENNA__08135__S net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11197__A2 net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14161_ clknet_leaf_16_clk _01335_ net1096 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.data_to_VGA\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_65_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11373_ net649 net184 vssd1 vssd1 vccd1 vccd1 _06061_ sky130_fd_sc_hd__and2_1
XANTENNA__13200__CLK clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input60_A mem_adr_start[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10324_ net1535 net1009 net986 final_design.data_from_mem\[9\] vssd1 vssd1 vccd1
+ vccd1 _00081_ sky130_fd_sc_hd__a22o_1
X_13112_ clknet_leaf_62_clk _00343_ net1119 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[100\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_46_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14092_ clknet_leaf_20_clk _01289_ net1161 vssd1 vssd1 vccd1 vccd1 final_design.reqhand.instruction\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11496__S net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10255_ final_design.uart.BAUD_counter\[19\] final_design.uart.BAUD_counter\[20\]
+ _05119_ vssd1 vssd1 vccd1 vccd1 _05123_ sky130_fd_sc_hd__and3_1
X_13043_ clknet_leaf_40_clk _00274_ net1210 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08445__S0 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1200 net1201 vssd1 vssd1 vccd1 vccd1 net1200 sky130_fd_sc_hd__clkbuf_4
Xfanout1211 net1212 vssd1 vssd1 vccd1 vccd1 net1211 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_37_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12889__Q final_design.data_from_mem\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13350__CLK clknet_leaf_51_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10186_ final_design.uart.BAUD_counter\[13\] final_design.uart.BAUD_counter\[12\]
+ final_design.uart.BAUD_counter\[15\] final_design.uart.BAUD_counter\[14\] vssd1
+ vssd1 vccd1 vccd1 _05076_ sky130_fd_sc_hd__or4_1
Xfanout1222 net1223 vssd1 vssd1 vccd1 vccd1 net1222 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_33_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1233 net1234 vssd1 vssd1 vccd1 vccd1 net1233 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_33_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1244 net1245 vssd1 vssd1 vccd1 vccd1 net1244 sky130_fd_sc_hd__buf_2
XANTENNA__12918__CLK clknet_leaf_62_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout290 _06228_ vssd1 vssd1 vccd1 vccd1 net290 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07562__X _02513_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13945_ clknet_leaf_54_clk _01176_ net1177 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[933\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_1905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11121__A2 net1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12120__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1140 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13876_ clknet_leaf_8_clk _01107_ net1154 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[864\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09078__A1 _03655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12827_ net1354 vssd1 vssd1 vccd1 vccd1 _00268_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__11244__B _01480_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12779__10 clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 net1320 sky130_fd_sc_hd__inv_2
XANTENNA__12082__B1 _06264_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12758_ _06383_ _06390_ _06391_ net796 final_design.VGA_adr\[6\] vssd1 vssd1 vccd1
+ vccd1 _06395_ sky130_fd_sc_hd__a32o_1
XFILLER_0_70_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07184__S0 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11709_ net200 net627 vssd1 vssd1 vccd1 vccd1 _06213_ sky130_fd_sc_hd__and2_1
XFILLER_0_38_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10575__S net1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12689_ _01401_ _05038_ vssd1 vssd1 vccd1 vccd1 _06332_ sky130_fd_sc_hd__nor2_1
XFILLER_0_71_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12385__A1 _06017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold705 final_design.cpu.reg_window\[1002\] vssd1 vssd1 vccd1 vccd1 net2047 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold716 final_design.cpu.reg_window\[504\] vssd1 vssd1 vccd1 vccd1 net2058 sky130_fd_sc_hd__dlygate4sd3_1
Xhold727 final_design.cpu.reg_window\[343\] vssd1 vssd1 vccd1 vccd1 net2069 sky130_fd_sc_hd__dlygate4sd3_1
Xhold738 final_design.cpu.reg_window\[436\] vssd1 vssd1 vccd1 vccd1 net2080 sky130_fd_sc_hd__dlygate4sd3_1
Xhold749 final_design.cpu.reg_window\[491\] vssd1 vssd1 vccd1 vccd1 net2091 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11259__X _05960_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08920_ final_design.CPU_instr_adr\[22\] _01756_ _03862_ vssd1 vssd1 vccd1 vccd1
+ _03863_ sky130_fd_sc_hd__a21o_1
XFILLER_0_21_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_17_clk_X clknet_leaf_17_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11345__C1 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11896__A0 net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09952__X _04871_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08851_ final_design.CPU_instr_adr\[30\] _03801_ vssd1 vssd1 vccd1 vccd1 _03802_
+ sky130_fd_sc_hd__nand2_1
XANTENNA__11360__A2 net235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07802_ final_design.cpu.reg_window\[793\] final_design.cpu.reg_window\[825\] net851
+ vssd1 vssd1 vccd1 vccd1 _02753_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08782_ _03688_ _03732_ vssd1 vssd1 vccd1 vccd1 _03733_ sky130_fd_sc_hd__nand2b_1
XANTENNA__13843__CLK clknet_leaf_40_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08568__X _03519_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07472__X _02423_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07733_ _02680_ _02681_ _02682_ _02683_ net686 net704 vssd1 vssd1 vccd1 vccd1 _02684_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__11648__B1 net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout178_A _06081_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12030__S net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07664_ final_design.cpu.reg_window\[414\] final_design.cpu.reg_window\[446\] net851
+ vssd1 vssd1 vccd1 vccd1 _02615_ sky130_fd_sc_hd__mux2_1
XANTENNA__10320__B1 net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07124__S net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09403_ _02576_ _02606_ _04171_ vssd1 vssd1 vccd1 vccd1 _04322_ sky130_fd_sc_hd__nand3_1
X_06615_ net884 _01559_ _01565_ _01547_ _01553_ vssd1 vssd1 vccd1 vccd1 _01566_ sky130_fd_sc_hd__a32oi_4
XANTENNA__13993__CLK clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13423__Q final_design.cpu.reg_window\[411\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07595_ _01539_ net605 vssd1 vssd1 vccd1 vccd1 _02546_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout345_A net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1087_A net1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09334_ _04249_ _04251_ vssd1 vssd1 vccd1 vccd1 _04253_ sky130_fd_sc_hd__xnor2_1
X_06546_ _01485_ _01489_ net731 _01495_ vssd1 vssd1 vccd1 vccd1 _01497_ sky130_fd_sc_hd__and4_4
XFILLER_0_36_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12073__B1 net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08277__C1 net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12612__A2 net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10623__A1 net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11820__A0 net219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09265_ net71 _04183_ vssd1 vssd1 vccd1 vccd1 _04184_ sky130_fd_sc_hd__or2_1
X_12778__9 clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 net1319 sky130_fd_sc_hd__inv_2
X_06477_ final_design.cpu.reg_window\[478\] final_design.cpu.reg_window\[510\] net933
+ vssd1 vssd1 vccd1 vccd1 _01428_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_1235 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13223__CLK clknet_leaf_62_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout512_A net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_748 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06922__S0 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11170__A net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08216_ _03103_ _03166_ vssd1 vssd1 vccd1 vccd1 _03167_ sky130_fd_sc_hd__nand2_1
X_09196_ _02545_ net445 _04096_ _04114_ vssd1 vssd1 vccd1 vccd1 _04115_ sky130_fd_sc_hd__o211a_1
XANTENNA__12376__A1 net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11179__A2 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout300_X net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08147_ _02030_ net611 vssd1 vssd1 vccd1 vccd1 _03098_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout1042_X net1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08044__A2 _02991_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07794__S net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09575__A net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09792__A2 _02091_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08078_ _03028_ vssd1 vssd1 vccd1 vccd1 _03029_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_8_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13373__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout881_A net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout979_A net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07029_ _01976_ _01977_ _01978_ _01979_ net765 net780 vssd1 vssd1 vccd1 vccd1 _01980_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_41_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06711__B _01660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10040_ _04637_ _04924_ _04958_ _04574_ vssd1 vssd1 vccd1 vccd1 _04959_ sky130_fd_sc_hd__and4b_1
XANTENNA__11887__A0 _05875_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold10 final_design.cpu.reg_window\[24\] vssd1 vssd1 vccd1 vccd1 net1352 sky130_fd_sc_hd__dlygate4sd3_1
Xhold21 final_design.cpu.reg_window\[26\] vssd1 vssd1 vccd1 vccd1 net1363 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout767_X net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold32 final_design.cpu.reg_window\[9\] vssd1 vssd1 vccd1 vccd1 net1374 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_51_1940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold43 final_design.reqhand.instruction\[16\] vssd1 vssd1 vccd1 vccd1 net1385 sky130_fd_sc_hd__dlygate4sd3_1
Xhold54 net151 vssd1 vssd1 vccd1 vccd1 net1396 sky130_fd_sc_hd__dlygate4sd3_1
Xhold65 final_design.reqhand.instruction\[23\] vssd1 vssd1 vccd1 vccd1 net1407 sky130_fd_sc_hd__dlygate4sd3_1
Xhold76 net145 vssd1 vssd1 vccd1 vccd1 net1418 sky130_fd_sc_hd__dlygate4sd3_1
Xhold87 net106 vssd1 vssd1 vccd1 vccd1 net1429 sky130_fd_sc_hd__dlygate4sd3_1
Xhold98 final_design.VGA_data_control.data_to_VGA\[15\] vssd1 vssd1 vccd1 vccd1 net1440
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout934_X net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11991_ net230 net2464 net400 vssd1 vssd1 vccd1 vccd1 _00723_ sky130_fd_sc_hd__mux2_1
XANTENNA__12300__A1 net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13730_ clknet_leaf_4_clk _00961_ net1079 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[718\]
+ sky130_fd_sc_hd__dfrtp_1
X_10942_ _05646_ _05667_ _05663_ vssd1 vssd1 vccd1 vccd1 _05670_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_39_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13661_ clknet_leaf_2_clk _00892_ net1064 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[649\]
+ sky130_fd_sc_hd__dfrtp_1
X_10873_ _05508_ _05542_ _05603_ _05604_ vssd1 vssd1 vccd1 vccd1 _05605_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_49_1880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1873 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12612_ net1437 net997 net983 final_design.data_from_mem\[30\] vssd1 vssd1 vccd1
+ vccd1 _01305_ sky130_fd_sc_hd__a22o_1
XFILLER_0_6_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12064__B1 net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13592_ clknet_leaf_65_clk _00823_ net1073 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[580\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_45_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08654__A _01566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1879 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11811__A0 net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12543_ _06206_ net344 net322 net1858 vssd1 vssd1 vccd1 vccd1 _01247_ sky130_fd_sc_hd__a22o_1
XFILLER_0_48_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12474_ _06134_ net343 net330 net2390 vssd1 vssd1 vccd1 vccd1 _01180_ sky130_fd_sc_hd__a22o_1
XANTENNA__10408__B _05181_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12367__A1 net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13716__CLK clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14213_ net1271 vssd1 vssd1 vccd1 vccd1 gpio_oeb[25] sky130_fd_sc_hd__buf_2
XFILLER_0_69_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11425_ net1839 net205 net310 vssd1 vssd1 vccd1 vccd1 _00322_ sky130_fd_sc_hd__mux2_1
XANTENNA__10378__B1 net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_7 _05934_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14144_ clknet_leaf_19_clk _01318_ net1157 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.data_to_VGA\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_11356_ net649 net189 vssd1 vssd1 vccd1 vccd1 _06046_ sky130_fd_sc_hd__and2_2
XTAP_TAPCELL_ROW_39_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10307_ _01384_ net1048 _05160_ vssd1 vssd1 vccd1 vccd1 _05161_ sky130_fd_sc_hd__or3b_1
XANTENNA__12115__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14075_ clknet_leaf_14_clk _01272_ net1107 vssd1 vssd1 vccd1 vccd1 final_design.uart.working_data\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11287_ net663 _03912_ net738 vssd1 vssd1 vccd1 vccd1 _05985_ sky130_fd_sc_hd__a21o_1
XANTENNA__13866__CLK clknet_leaf_59_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13026_ clknet_leaf_3_clk _00257_ net1066 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_10238_ final_design.uart.BAUD_counter\[13\] final_design.uart.BAUD_counter\[12\]
+ _05108_ final_design.uart.BAUD_counter\[14\] vssd1 vssd1 vccd1 vccd1 _05112_ sky130_fd_sc_hd__a31o_1
XANTENNA__11878__B1 net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1030 net1036 vssd1 vssd1 vccd1 vccd1 net1030 sky130_fd_sc_hd__buf_4
XFILLER_0_20_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1041 _01393_ vssd1 vssd1 vccd1 vccd1 net1041 sky130_fd_sc_hd__buf_2
X_10169_ final_design.vga.h_current_state\[0\] final_design.vga.h_current_state\[1\]
+ _05044_ vssd1 vssd1 vccd1 vccd1 _05061_ sky130_fd_sc_hd__o21ai_1
Xfanout1052 final_design.uart.receiving vssd1 vssd1 vccd1 vccd1 net1052 sky130_fd_sc_hd__buf_2
Xfanout1063 net1069 vssd1 vssd1 vccd1 vccd1 net1063 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_59_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1074 net1075 vssd1 vssd1 vccd1 vccd1 net1074 sky130_fd_sc_hd__clkbuf_4
Xfanout1085 net1118 vssd1 vssd1 vccd1 vccd1 net1085 sky130_fd_sc_hd__clkbuf_2
XANTENNA__12890__CLK clknet_leaf_18_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1096 net1117 vssd1 vssd1 vccd1 vccd1 net1096 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_16_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13928_ clknet_leaf_41_clk _01159_ net1225 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[916\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07849__A2 _02797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13859_ clknet_leaf_64_clk _01090_ net1075 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[847\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_44_clk_A clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13246__CLK clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06521__A2 final_design.data_from_mem\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1913 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07380_ _02326_ _02330_ vssd1 vssd1 vccd1 vccd1 _02331_ sky130_fd_sc_hd__nand2_1
XANTENNA__06783__S net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1733 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11802__B1 net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09379__B _04097_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_2280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_2291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09050_ _02442_ _03978_ vssd1 vssd1 vccd1 vccd1 _03979_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_2_1777 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_59_clk_A clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13396__CLK clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08001_ final_design.cpu.reg_window\[976\] final_design.cpu.reg_window\[1008\] net843
+ vssd1 vssd1 vccd1 vccd1 _02952_ sky130_fd_sc_hd__mux2_1
XANTENNA__10369__B1 net1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold502 final_design.cpu.reg_window\[839\] vssd1 vssd1 vccd1 vccd1 net1844 sky130_fd_sc_hd__dlygate4sd3_1
Xhold513 final_design.cpu.reg_window\[1017\] vssd1 vssd1 vccd1 vccd1 net1855 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold524 final_design.cpu.reg_window\[905\] vssd1 vssd1 vccd1 vccd1 net1866 sky130_fd_sc_hd__dlygate4sd3_1
Xhold535 final_design.cpu.reg_window\[591\] vssd1 vssd1 vccd1 vccd1 net1877 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkload32_A clknet_leaf_41_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold546 final_design.cpu.reg_window\[44\] vssd1 vssd1 vccd1 vccd1 net1888 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06588__A2 _01537_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold557 final_design.cpu.reg_window\[55\] vssd1 vssd1 vccd1 vccd1 net1899 sky130_fd_sc_hd__dlygate4sd3_1
Xhold568 final_design.cpu.reg_window\[258\] vssd1 vssd1 vccd1 vccd1 net1910 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11581__A2 net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold579 final_design.cpu.reg_window\[730\] vssd1 vssd1 vccd1 vccd1 net1921 sky130_fd_sc_hd__dlygate4sd3_1
X_09952_ net495 _04868_ _04869_ _04870_ vssd1 vssd1 vccd1 vccd1 _04871_ sky130_fd_sc_hd__a22o_2
XTAP_TAPCELL_ROW_55_2073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_55_2084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_2095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07119__S net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08903_ _01661_ _01662_ _02469_ vssd1 vssd1 vccd1 vccd1 _03848_ sky130_fd_sc_hd__or3_1
XANTENNA__11869__B1 net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09883_ _04341_ _04801_ vssd1 vssd1 vccd1 vccd1 _04802_ sky130_fd_sc_hd__or2_1
XANTENNA__11333__A2 net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout295_A _06194_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1202 final_design.VGA_data_control.state\[1\] vssd1 vssd1 vccd1 vccd1 net2544
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08834_ final_design.CPU_instr_adr\[5\] _03784_ vssd1 vssd1 vccd1 vccd1 _03785_ sky130_fd_sc_hd__and2_1
Xhold1213 final_design.reqhand.instruction\[4\] vssd1 vssd1 vccd1 vccd1 net2555 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_57_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1002_A net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10988__B net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14021__CLK clknet_leaf_49_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08765_ final_design.CPU_instr_adr\[1\] _02391_ _02393_ vssd1 vssd1 vccd1 vccd1 _03716_
+ sky130_fd_sc_hd__nand3b_1
XFILLER_0_79_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout462_A net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07716_ net711 _02666_ net877 vssd1 vssd1 vccd1 vccd1 _02667_ sky130_fd_sc_hd__o21ai_1
XANTENNA__12294__B1 net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1600 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08696_ _01487_ _03646_ _02094_ vssd1 vssd1 vccd1 vccd1 _03647_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_73_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout250_X net250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07647_ final_design.cpu.reg_window\[604\] final_design.cpu.reg_window\[636\] net867
+ vssd1 vssd1 vccd1 vccd1 _02598_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout727_A _01493_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout348_X net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14171__CLK clknet_leaf_19_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07578_ final_design.cpu.reg_window\[543\] final_design.cpu.reg_window\[575\] net857
+ vssd1 vssd1 vccd1 vccd1 _02529_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13739__CLK clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12597__B2 final_design.data_from_mem\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09317_ net476 _04235_ vssd1 vssd1 vccd1 vccd1 _04236_ sky130_fd_sc_hd__nor2_1
X_06529_ _01478_ _01479_ vssd1 vssd1 vccd1 vccd1 _01480_ sky130_fd_sc_hd__nand2_2
XANTENNA_fanout515_X net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09248_ _04158_ _04164_ _04166_ _04133_ vssd1 vssd1 vccd1 vccd1 _04167_ sky130_fd_sc_hd__a211o_1
XFILLER_0_35_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09179_ _02502_ net468 net459 vssd1 vssd1 vccd1 vccd1 _04098_ sky130_fd_sc_hd__or3_1
XANTENNA__13889__CLK clknet_leaf_47_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11021__A1 net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11210_ _03620_ _05854_ _05906_ vssd1 vssd1 vccd1 vccd1 _05917_ sky130_fd_sc_hd__and3_2
X_12190_ net1934 net187 net383 vssd1 vssd1 vccd1 vccd1 _00909_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout884_X net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11141_ final_design.reqhand.data_from_UART\[0\] final_design.data_from_mem\[0\]
+ net245 vssd1 vssd1 vccd1 vccd1 _05856_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07871__S1 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13119__CLK clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11072_ _05773_ _05791_ vssd1 vssd1 vccd1 vccd1 _05795_ sky130_fd_sc_hd__and2_1
Xinput100 nrst vssd1 vssd1 vccd1 vccd1 net100 sky130_fd_sc_hd__clkbuf_8
X_10023_ net68 _04940_ vssd1 vssd1 vccd1 vccd1 _04942_ sky130_fd_sc_hd__or2_1
XANTENNA_input23_A DAT_I[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13269__CLK clknet_leaf_56_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12285__B1 net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11974_ _06176_ net287 net406 net2035 vssd1 vssd1 vccd1 vccd1 _00707_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_47_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_47_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13713_ clknet_leaf_35_clk _00944_ net1240 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[701\]
+ sky130_fd_sc_hd__dfrtp_1
X_10925_ _05652_ _05653_ _05632_ _05634_ vssd1 vssd1 vccd1 vccd1 _05654_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_6_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07699__S net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13644_ clknet_leaf_45_clk _00875_ net1213 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[632\]
+ sky130_fd_sc_hd__dfrtp_1
X_10856_ net80 net1044 vssd1 vssd1 vccd1 vccd1 _05588_ sky130_fd_sc_hd__and2_1
XFILLER_0_71_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12588__B2 final_design.data_from_mem\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13575_ clknet_leaf_62_clk _00806_ net1120 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[563\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09199__B net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09453__A1 net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10787_ net43 _05521_ vssd1 vssd1 vccd1 vccd1 _05523_ sky130_fd_sc_hd__nor2_1
XANTENNA__10419__A _03224_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1717 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11260__A1 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12526_ _06188_ net357 net328 net2196 vssd1 vssd1 vccd1 vccd1 _01231_ sky130_fd_sc_hd__a22o_1
XFILLER_0_54_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10853__S net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12457_ net2483 net188 net336 vssd1 vssd1 vccd1 vccd1 _01164_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_10_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11408_ net805 _02359_ net803 vssd1 vssd1 vccd1 vccd1 _06091_ sky130_fd_sc_hd__and3b_1
X_12388_ net1822 net191 net271 vssd1 vssd1 vccd1 vccd1 _01099_ sky130_fd_sc_hd__mux2_1
XANTENNA__06931__A_N net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14127_ clknet_leaf_20_clk final_design.vga.v_next_count\[7\] net1160 vssd1 vssd1
+ vccd1 vccd1 final_design.VGA_data_control.v_count\[7\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_22_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11339_ _06027_ _06029_ _06030_ net590 vssd1 vssd1 vccd1 vccd1 _06031_ sky130_fd_sc_hd__o211a_1
XANTENNA__14044__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14058_ clknet_leaf_16_clk _00020_ net1092 vssd1 vssd1 vccd1 vccd1 final_design.uart.BAUD_counter\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_78_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11315__A2 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13009_ net1340 _00240_ net1234 vssd1 vssd1 vccd1 vccd1 final_design.CPU_instr_adr\[29\]
+ sky130_fd_sc_hd__dfrtp_4
X_06880_ net751 _01830_ vssd1 vssd1 vccd1 vccd1 _01831_ sky130_fd_sc_hd__nor2_1
XFILLER_0_78_1857 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08550_ final_design.cpu.reg_window\[833\] final_design.cpu.reg_window\[865\] net838
+ vssd1 vssd1 vccd1 vccd1 _03501_ sky130_fd_sc_hd__mux2_1
XANTENNA__12276__B1 net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07501_ _02002_ _02450_ _02001_ vssd1 vssd1 vccd1 vccd1 _02452_ sky130_fd_sc_hd__o21a_1
X_08481_ final_design.cpu.reg_window\[67\] final_design.cpu.reg_window\[99\] net824
+ vssd1 vssd1 vccd1 vccd1 _03432_ sky130_fd_sc_hd__mux2_1
XANTENNA__12291__A3 net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_63_2342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11713__A net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_2353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07432_ final_design.cpu.reg_window\[705\] final_design.cpu.reg_window\[737\] net914
+ vssd1 vssd1 vccd1 vccd1 _02383_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_63_2364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_2375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06807__A net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1863 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07402__S net913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07363_ final_design.cpu.reg_window\[771\] final_design.cpu.reg_window\[803\] net917
+ vssd1 vssd1 vccd1 vccd1 _02314_ sky130_fd_sc_hd__mux2_1
XANTENNA__06526__B _01468_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_759 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09102_ _02364_ _02429_ net619 vssd1 vssd1 vccd1 vccd1 _04024_ sky130_fd_sc_hd__a21o_1
XANTENNA__10054__A2 _04940_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11251__A1 final_design.data_from_mem\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07294_ final_design.cpu.reg_window\[197\] final_design.cpu.reg_window\[229\] net919
+ vssd1 vssd1 vccd1 vccd1 _02245_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09033_ final_design.CPU_instr_adr\[11\] _03788_ vssd1 vssd1 vccd1 vccd1 _03964_
+ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout210_A net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout308_A net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07638__A net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_2146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold310 final_design.uart.BAUD_counter\[19\] vssd1 vssd1 vccd1 vccd1 net1652 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12200__B1 net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08404__C1 _02239_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_2157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold321 final_design.cpu.reg_window\[912\] vssd1 vssd1 vccd1 vccd1 net1663 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_2168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold332 final_design.cpu.reg_window\[134\] vssd1 vssd1 vccd1 vccd1 net1674 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07302__S0 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold343 final_design.cpu.reg_window\[138\] vssd1 vssd1 vccd1 vccd1 net1685 sky130_fd_sc_hd__dlygate4sd3_1
Xhold354 final_design.cpu.reg_window\[235\] vssd1 vssd1 vccd1 vccd1 net1696 sky130_fd_sc_hd__dlygate4sd3_1
Xhold365 final_design.cpu.reg_window\[177\] vssd1 vssd1 vccd1 vccd1 net1707 sky130_fd_sc_hd__dlygate4sd3_1
Xhold376 final_design.cpu.reg_window\[982\] vssd1 vssd1 vccd1 vccd1 net1718 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1217_A net1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold387 final_design.cpu.reg_window\[780\] vssd1 vssd1 vccd1 vccd1 net1729 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout801 net802 vssd1 vssd1 vccd1 vccd1 net801 sky130_fd_sc_hd__buf_4
Xhold398 final_design.cpu.reg_window\[752\] vssd1 vssd1 vccd1 vccd1 net1740 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_61_1861 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09935_ net489 _04619_ _04852_ _04853_ _04341_ vssd1 vssd1 vccd1 vccd1 _04854_ sky130_fd_sc_hd__a221o_1
Xfanout812 net815 vssd1 vssd1 vccd1 vccd1 net812 sky130_fd_sc_hd__clkbuf_4
Xfanout823 net824 vssd1 vssd1 vccd1 vccd1 net823 sky130_fd_sc_hd__clkbuf_4
Xfanout834 net842 vssd1 vssd1 vccd1 vccd1 net834 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout677_A net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout845 net847 vssd1 vssd1 vccd1 vccd1 net845 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout298_X net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1282 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout856 net872 vssd1 vssd1 vccd1 vccd1 net856 sky130_fd_sc_hd__buf_2
XANTENNA__13411__CLK clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09866_ _03294_ _03568_ vssd1 vssd1 vccd1 vccd1 _04785_ sky130_fd_sc_hd__xnor2_1
Xfanout867 net872 vssd1 vssd1 vccd1 vccd1 net867 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout1005_X net1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1010 final_design.cpu.reg_window\[375\] vssd1 vssd1 vccd1 vccd1 net2352 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout878 net879 vssd1 vssd1 vccd1 vccd1 net878 sky130_fd_sc_hd__clkbuf_8
XANTENNA__07605__S1 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1021 final_design.cpu.reg_window\[183\] vssd1 vssd1 vccd1 vccd1 net2363 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09380__A0 net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout889 net890 vssd1 vssd1 vccd1 vccd1 net889 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07373__A net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08817_ _03753_ _03763_ _03767_ vssd1 vssd1 vccd1 vccd1 _03768_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_5_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1032 final_design.cpu.reg_window\[501\] vssd1 vssd1 vccd1 vccd1 net2374 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1043 final_design.cpu.reg_window\[931\] vssd1 vssd1 vccd1 vccd1 net2385 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11607__B net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout844_A net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09797_ _03358_ net446 _04242_ _04086_ _04715_ vssd1 vssd1 vccd1 vccd1 _04716_ sky130_fd_sc_hd__o221a_1
Xhold1054 final_design.cpu.reg_window\[106\] vssd1 vssd1 vccd1 vccd1 net2396 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1065 final_design.cpu.reg_window\[300\] vssd1 vssd1 vccd1 vccd1 net2407 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1076 final_design.cpu.reg_window\[812\] vssd1 vssd1 vccd1 vccd1 net2418 sky130_fd_sc_hd__dlygate4sd3_1
X_08748_ _03697_ _03698_ vssd1 vssd1 vccd1 vccd1 _03699_ sky130_fd_sc_hd__nand2b_1
XANTENNA__12267__B1 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1087 final_design.cpu.reg_window\[110\] vssd1 vssd1 vccd1 vccd1 net2429 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1098 final_design.cpu.reg_window\[114\] vssd1 vssd1 vccd1 vccd1 net2440 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_67_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13561__CLK clknet_leaf_54_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1616 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08679_ _03629_ vssd1 vssd1 vccd1 vccd1 _03630_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout632_X net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12282__A3 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10710_ _05447_ _05448_ vssd1 vssd1 vccd1 vccd1 _05449_ sky130_fd_sc_hd__nand2_1
XANTENNA__11623__A net219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12019__B1 net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11690_ net426 net556 _06203_ net294 net1889 vssd1 vssd1 vccd1 vccd1 _00476_ sky130_fd_sc_hd__a32o_1
XANTENNA__06717__A net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10641_ _05347_ _05364_ _05383_ _05362_ vssd1 vssd1 vccd1 vccd1 _05384_ sky130_fd_sc_hd__a211o_1
XFILLER_0_10_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13088__RESET_B net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13360_ clknet_leaf_33_clk _00591_ net1238 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[348\]
+ sky130_fd_sc_hd__dfrtp_1
X_10572_ _05291_ _05294_ _05316_ vssd1 vssd1 vccd1 vccd1 _05318_ sky130_fd_sc_hd__o21ai_1
XANTENNA__11793__A2 net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12311_ net1787 net207 net364 vssd1 vssd1 vccd1 vccd1 _01025_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_1447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11769__S net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13291_ clknet_leaf_38_clk _00522_ net1189 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[279\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12242_ net559 _06172_ net504 net372 net1482 vssd1 vssd1 vccd1 vccd1 _00959_ sky130_fd_sc_hd__a32o_1
XANTENNA__06452__A net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14067__CLK clknet_leaf_15_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11545__A2 net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12173_ net1786 net218 net380 vssd1 vssd1 vccd1 vccd1 _00892_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1901 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07844__S1 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11124_ net672 _02358_ _05838_ vssd1 vssd1 vccd1 vccd1 _05839_ sky130_fd_sc_hd__or3_4
XFILLER_0_60_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13091__CLK clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11055_ _04325_ net248 net669 vssd1 vssd1 vccd1 vccd1 _05778_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12897__Q final_design.data_from_mem\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10006_ _04614_ _04615_ vssd1 vssd1 vccd1 vccd1 _04925_ sky130_fd_sc_hd__nor2_1
XANTENNA__13904__CLK clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10421__B _05190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12258__B1 net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08666__X _03617_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11957_ net427 net555 net630 vssd1 vssd1 vccd1 vccd1 _06256_ sky130_fd_sc_hd__and3_1
XFILLER_0_80_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12273__A3 net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06488__A1 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10908_ net959 _05636_ _05637_ net956 vssd1 vssd1 vccd1 vccd1 _05638_ sky130_fd_sc_hd__o22a_1
XFILLER_0_74_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11888_ net227 net2092 net272 vssd1 vssd1 vccd1 vccd1 _00630_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13627_ clknet_leaf_66_clk _00858_ net1063 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[615\]
+ sky130_fd_sc_hd__dfrtp_1
X_10839_ _05570_ _05571_ vssd1 vssd1 vccd1 vccd1 _05572_ sky130_fd_sc_hd__xor2_1
XFILLER_0_27_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1861 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11233__A1 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13558_ clknet_leaf_61_clk _00789_ net1136 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[546\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_150 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12509_ _06171_ net347 net326 net1577 vssd1 vssd1 vccd1 vccd1 _01214_ sky130_fd_sc_hd__a22o_1
X_13489_ clknet_leaf_35_clk _00720_ net1240 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[477\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_879 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09729__A2 net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_2780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_2622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_2633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13434__CLK clknet_leaf_58_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_2644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07981_ net603 _02929_ _02905_ net545 vssd1 vssd1 vccd1 vccd1 _02932_ sky130_fd_sc_hd__o211a_1
X_09720_ _04627_ _04638_ net449 vssd1 vssd1 vccd1 vccd1 _04639_ sky130_fd_sc_hd__a21o_1
X_06932_ net546 _01881_ vssd1 vssd1 vccd1 vccd1 _01883_ sky130_fd_sc_hd__xor2_1
XANTENNA__12303__S net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13584__CLK clknet_leaf_36_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09651_ net448 _04569_ _04566_ vssd1 vssd1 vccd1 vccd1 _04570_ sky130_fd_sc_hd__o21a_2
XFILLER_0_78_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06863_ net761 _01813_ net886 vssd1 vssd1 vccd1 vccd1 _01814_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_59_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_69_2551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08260__S1 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_2562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07912__B2 net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08602_ net596 _03550_ _03524_ _02419_ vssd1 vssd1 vccd1 vccd1 _03553_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_69_2573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12249__B1 net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_2415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09582_ _03582_ _04499_ _03134_ vssd1 vssd1 vccd1 vccd1 _04501_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_65_2426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06794_ final_design.cpu.reg_window\[790\] final_design.cpu.reg_window\[822\] net918
+ vssd1 vssd1 vccd1 vccd1 _01745_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_65_2437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08533_ net609 _03481_ _03482_ vssd1 vssd1 vccd1 vccd1 _03484_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_52_1805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09665__A1 net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08468__A2 _03415_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09665__B2 net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout258_A net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08464_ _03402_ _03403_ _03414_ net875 vssd1 vssd1 vccd1 vccd1 _03415_ sky130_fd_sc_hd__a22oi_4
XFILLER_0_72_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07415_ final_design.cpu.reg_window\[257\] final_design.cpu.reg_window\[289\] net922
+ vssd1 vssd1 vccd1 vccd1 _02366_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09417__A1 _01566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08395_ final_design.cpu.reg_window\[710\] final_design.cpu.reg_window\[742\] net820
+ vssd1 vssd1 vccd1 vccd1 _03346_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout425_A net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1167_A net100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11224__A1 net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10027__A2 net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12421__B1 net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07346_ net744 net666 net724 _01496_ _02296_ vssd1 vssd1 vccd1 vccd1 _02297_ sky130_fd_sc_hd__o221a_1
XANTENNA__09848__A net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_2208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_2219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_1579 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11775__A2 net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07277_ final_design.cpu.reg_window\[838\] final_design.cpu.reg_window\[870\] net912
+ vssd1 vssd1 vccd1 vccd1 _02228_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout213_X net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09016_ final_design.CPU_instr_adr\[12\] _03789_ final_design.CPU_instr_adr\[13\]
+ vssd1 vssd1 vccd1 vccd1 _03949_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_41_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout794_A net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold140 final_design.cpu.reg_window\[716\] vssd1 vssd1 vccd1 vccd1 net1482 sky130_fd_sc_hd__dlygate4sd3_1
Xhold151 final_design.cpu.reg_window\[222\] vssd1 vssd1 vccd1 vccd1 net1493 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold162 final_design.VGA_data_control.ready_data\[18\] vssd1 vssd1 vccd1 vccd1 net1504
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold173 final_design.cpu.reg_window\[728\] vssd1 vssd1 vccd1 vccd1 net1515 sky130_fd_sc_hd__dlygate4sd3_1
Xhold184 final_design.VGA_data_control.ready_data\[4\] vssd1 vssd1 vccd1 vccd1 net1526
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold195 final_design.cpu.reg_window\[706\] vssd1 vssd1 vccd1 vccd1 net1537 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout961_A _04036_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13927__CLK clknet_leaf_62_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout582_X net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout620 _02507_ vssd1 vssd1 vccd1 vccd1 net620 sky130_fd_sc_hd__buf_2
Xfanout631 _06157_ vssd1 vssd1 vccd1 vccd1 net631 sky130_fd_sc_hd__buf_4
Xfanout642 _05946_ vssd1 vssd1 vccd1 vccd1 net642 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07374__Y _02325_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09918_ net484 _04407_ _04835_ _04219_ vssd1 vssd1 vccd1 vccd1 _04837_ sky130_fd_sc_hd__o211ai_1
XANTENNA__12488__B1 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout653 net654 vssd1 vssd1 vccd1 vccd1 net653 sky130_fd_sc_hd__clkbuf_4
Xfanout675 net676 vssd1 vssd1 vccd1 vccd1 net675 sky130_fd_sc_hd__buf_4
Xfanout686 net688 vssd1 vssd1 vccd1 vccd1 net686 sky130_fd_sc_hd__buf_4
X_09849_ _04751_ _04767_ vssd1 vssd1 vccd1 vccd1 _04768_ sky130_fd_sc_hd__xnor2_1
Xfanout697 net698 vssd1 vssd1 vccd1 vccd1 net697 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout847_X net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12951__CLK clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12860_ clknet_leaf_18_clk _00098_ net1106 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.ready_data\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11811_ net231 net2279 net264 vssd1 vssd1 vccd1 vccd1 _00563_ sky130_fd_sc_hd__mux2_1
XANTENNA__08003__S1 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12255__A3 net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11742_ net238 net2263 net416 vssd1 vssd1 vccd1 vccd1 _00505_ sky130_fd_sc_hd__mux2_1
XANTENNA__13307__CLK clknet_leaf_65_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11673_ net228 net627 vssd1 vssd1 vccd1 vccd1 _06195_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_12_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_1801 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07977__S net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13412_ clknet_leaf_52_clk _00643_ net1174 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[400\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10018__A2 _03635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input90_A memory_size[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10624_ _04745_ net247 net668 vssd1 vssd1 vccd1 vccd1 _05367_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_12_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12412__B1 net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06881__S net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1845 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13343_ clknet_leaf_7_clk _00574_ net1145 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[331\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10555_ net63 _05301_ vssd1 vssd1 vccd1 vccd1 _05302_ sky130_fd_sc_hd__and2_1
XFILLER_0_52_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13457__CLK clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08631__A2 _03160_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1889 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13274_ clknet_leaf_58_clk _00505_ net1132 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[262\]
+ sky130_fd_sc_hd__dfrtp_1
X_10486_ net90 final_design.VGA_adr\[0\] vssd1 vssd1 vccd1 vccd1 _05236_ sky130_fd_sc_hd__or2_1
XFILLER_0_59_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12225_ net584 _06153_ net512 net378 net1803 vssd1 vssd1 vccd1 vccd1 _00943_ sky130_fd_sc_hd__a32o_1
XFILLER_0_20_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12156_ net187 net2208 net386 vssd1 vssd1 vccd1 vccd1 _00877_ sky130_fd_sc_hd__mux2_1
X_11107_ net60 _05827_ vssd1 vssd1 vccd1 vccd1 _05828_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12479__B1 net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12123__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12087_ net578 _06046_ net510 net394 net1596 vssd1 vssd1 vccd1 vccd1 _00812_ sky130_fd_sc_hd__a32o_1
XANTENNA__09344__B1 net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11038_ net88 net1045 vssd1 vssd1 vccd1 vccd1 _05762_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_1805 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_1849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09647__A1 _04046_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12989_ net1320 _00220_ net1166 vssd1 vssd1 vccd1 vccd1 final_design.CPU_instr_adr\[9\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_59_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07200_ final_design.cpu.reg_window\[713\] final_design.cpu.reg_window\[745\] net889
+ vssd1 vssd1 vccd1 vccd1 _02151_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12403__B1 net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08180_ _01967_ net612 vssd1 vssd1 vccd1 vccd1 _03131_ sky130_fd_sc_hd__nor2_1
XFILLER_0_12_1877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_2820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07131_ final_design.cpu.reg_window\[971\] final_design.cpu.reg_window\[1003\] net915
+ vssd1 vssd1 vccd1 vccd1 _02082_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_77_2831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_2842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08622__A2 _03257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07062_ _02009_ _02010_ _02011_ _02012_ net772 net795 vssd1 vssd1 vccd1 vccd1 _02013_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_73_2706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1219 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11390__B1 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12974__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12033__S net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07964_ final_design.cpu.reg_window\[145\] final_design.cpu.reg_window\[177\] net848
+ vssd1 vssd1 vccd1 vccd1 _02915_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09703_ net491 _04578_ _04579_ _04620_ _04341_ vssd1 vssd1 vccd1 vccd1 _04622_ sky130_fd_sc_hd__a311oi_1
XFILLER_0_78_1440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06915_ final_design.cpu.reg_window\[146\] final_design.cpu.reg_window\[178\] net920
+ vssd1 vssd1 vccd1 vccd1 _01866_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07895_ final_design.cpu.reg_window\[23\] final_design.cpu.reg_window\[55\] net849
+ vssd1 vssd1 vccd1 vccd1 _02846_ sky130_fd_sc_hd__mux2_1
XANTENNA__08689__A2 _03549_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09886__A1 net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout375_A _06272_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09886__B2 net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09634_ _02997_ _03031_ _04430_ vssd1 vssd1 vccd1 vccd1 _04553_ sky130_fd_sc_hd__or3_1
X_06846_ final_design.cpu.reg_window\[84\] final_design.cpu.reg_window\[116\] net948
+ vssd1 vssd1 vccd1 vccd1 _01797_ sky130_fd_sc_hd__mux2_1
XANTENNA__11444__Y _06095_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09565_ _03134_ _04087_ _04483_ vssd1 vssd1 vccd1 vccd1 _04484_ sky130_fd_sc_hd__a21oi_1
X_06777_ final_design.cpu.reg_window\[470\] final_design.cpu.reg_window\[502\] net920
+ vssd1 vssd1 vccd1 vccd1 _01728_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout542_A net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12237__A3 net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08516_ _03463_ _03464_ _03465_ _03466_ net679 net699 vssd1 vssd1 vccd1 vccd1 _03467_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_65_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09496_ net478 _04086_ _04412_ _04414_ _04269_ vssd1 vssd1 vccd1 vccd1 _04415_ sky130_fd_sc_hd__o311a_1
XANTENNA__07113__A2 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11996__A2 net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08447_ final_design.cpu.reg_window\[4\] final_design.cpu.reg_window\[36\] net821
+ vssd1 vssd1 vccd1 vccd1 _03398_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_1911 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout330_X net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout428_X net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07797__S net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08378_ final_design.cpu.reg_window\[454\] final_design.cpu.reg_window\[486\] net823
+ vssd1 vssd1 vccd1 vccd1 _03329_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_22_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06554__X _01505_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07329_ _02276_ _02277_ _02278_ _02279_ net767 net787 vssd1 vssd1 vccd1 vccd1 _02280_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__09297__B net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10340_ net1628 net1009 net986 final_design.data_from_mem\[25\] vssd1 vssd1 vccd1
+ vccd1 _00097_ sky130_fd_sc_hd__a22o_1
X_10271_ final_design.uart.BAUD_counter\[25\] final_design.uart.BAUD_counter\[26\]
+ _05129_ vssd1 vssd1 vccd1 vccd1 _05133_ sky130_fd_sc_hd__and3_1
XFILLER_0_44_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12010_ _06212_ net283 net402 net2147 vssd1 vssd1 vccd1 vccd1 _00741_ sky130_fd_sc_hd__a22o_1
XANTENNA__09574__B1 net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout964_X net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11348__A net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14105__CLK clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout450 _04069_ vssd1 vssd1 vccd1 vccd1 net450 sky130_fd_sc_hd__buf_4
Xfanout461 _03519_ vssd1 vssd1 vccd1 vccd1 net461 sky130_fd_sc_hd__buf_2
Xfanout472 net474 vssd1 vssd1 vccd1 vccd1 net472 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_35_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13961_ clknet_leaf_37_clk _01192_ net1235 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[949\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout483 net488 vssd1 vssd1 vccd1 vccd1 net483 sky130_fd_sc_hd__clkbuf_2
Xfanout494 net495 vssd1 vssd1 vccd1 vccd1 net494 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_31_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12912_ clknet_leaf_61_clk _00150_ net1136 vssd1 vssd1 vccd1 vccd1 net165 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_31_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11684__A1 net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13892_ clknet_leaf_52_clk _01123_ net1174 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[880\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_31_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07561__A net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12843_ clknet_leaf_15_clk _00081_ net1107 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.ready_data\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12228__A3 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11987__A2 net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11725_ net184 net628 vssd1 vssd1 vccd1 vccd1 _06221_ sky130_fd_sc_hd__and2_1
XFILLER_0_51_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_29_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09488__A net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06863__A1 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06464__X _01415_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11656_ net434 net577 _06185_ net300 net1520 vssd1 vssd1 vccd1 vccd1 _00460_ sky130_fd_sc_hd__a32o_1
XANTENNA__06905__A net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12847__CLK clknet_leaf_18_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10607_ _05331_ _05349_ _05350_ vssd1 vssd1 vccd1 vccd1 _05351_ sky130_fd_sc_hd__and3b_1
XFILLER_0_68_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12118__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11587_ net436 net582 _06149_ net304 net1633 vssd1 vssd1 vccd1 vccd1 _00427_ sky130_fd_sc_hd__a32o_1
XANTENNA__10427__A _03160_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06615__A1 net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13326_ clknet_leaf_43_clk _00557_ net1223 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[314\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10538_ _05268_ _05285_ vssd1 vssd1 vccd1 vccd1 _05286_ sky130_fd_sc_hd__xnor2_1
Xhold909 final_design.cpu.reg_window\[97\] vssd1 vssd1 vccd1 vccd1 net2251 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13257_ clknet_leaf_36_clk _00488_ net1229 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[245\]
+ sky130_fd_sc_hd__dfrtp_1
X_10469_ net36 _05220_ vssd1 vssd1 vccd1 vccd1 _05221_ sky130_fd_sc_hd__and2_1
XFILLER_0_20_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12208_ net565 _06136_ net505 net377 net1670 vssd1 vssd1 vccd1 vccd1 _00926_ sky130_fd_sc_hd__a32o_1
XFILLER_0_81_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13188_ clknet_leaf_54_clk _00419_ net1180 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[176\]
+ sky130_fd_sc_hd__dfrtp_1
X_12139_ net218 net2378 net384 vssd1 vssd1 vccd1 vccd1 _00860_ sky130_fd_sc_hd__mux2_1
XANTENNA__07455__B _02405_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07591__A2 _02540_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06700_ final_design.cpu.reg_window\[729\] final_design.cpu.reg_window\[761\] net930
+ vssd1 vssd1 vccd1 vccd1 _01651_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07680_ final_design.cpu.reg_window\[606\] final_design.cpu.reg_window\[638\] net851
+ vssd1 vssd1 vccd1 vccd1 _02631_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06631_ net761 _01581_ vssd1 vssd1 vccd1 vccd1 _01582_ sky130_fd_sc_hd__or2_1
XANTENNA__11705__B net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12219__A3 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13622__CLK clknet_leaf_62_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09350_ net494 _04268_ _04231_ vssd1 vssd1 vccd1 vccd1 _04269_ sky130_fd_sc_hd__a21o_1
X_06562_ final_design.cpu.reg_window\[477\] final_design.cpu.reg_window\[509\] net949
+ vssd1 vssd1 vccd1 vccd1 _01513_ sky130_fd_sc_hd__mux2_1
X_08301_ final_design.cpu.reg_window\[777\] final_design.cpu.reg_window\[809\] net810
+ vssd1 vssd1 vccd1 vccd1 _03252_ sky130_fd_sc_hd__mux2_1
XANTENNA__11978__A2 net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09281_ net551 net550 net549 net548 net458 net469 vssd1 vssd1 vccd1 vccd1 _04200_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_16_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_1764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06493_ _01440_ _01441_ _01442_ _01443_ net774 net792 vssd1 vssd1 vccd1 vccd1 _01444_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_74_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08573__Y _03524_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_2904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_79_2915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11721__A net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08232_ final_design.cpu.reg_window\[971\] final_design.cpu.reg_window\[1003\] net835
+ vssd1 vssd1 vccd1 vccd1 _03183_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13772__CLK clknet_leaf_46_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08163_ final_design.cpu.reg_window\[143\] final_design.cpu.reg_window\[175\] net807
+ vssd1 vssd1 vccd1 vccd1 _03114_ sky130_fd_sc_hd__mux2_1
XANTENNA__12028__S net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10938__B1 net1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07114_ _02059_ _02064_ vssd1 vssd1 vccd1 vccd1 _02065_ sky130_fd_sc_hd__nand2_1
XFILLER_0_71_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08094_ final_design.cpu.reg_window\[396\] final_design.cpu.reg_window\[428\] net817
+ vssd1 vssd1 vccd1 vccd1 _03045_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07045_ net882 _01988_ _01994_ _01981_ _01982_ vssd1 vssd1 vccd1 vccd1 _01996_ sky130_fd_sc_hd__a32o_4
XFILLER_0_42_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14128__CLK clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1032_A net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09020__A2 net1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout492_A net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11363__B1 net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07031__A1 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10072__A net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08996_ net255 _03930_ net1016 vssd1 vssd1 vccd1 vccd1 _03931_ sky130_fd_sc_hd__a21oi_1
X_07947_ _01750_ _02896_ vssd1 vssd1 vccd1 vccd1 _02898_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout280_X net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09859__A1 net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout378_X net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout757_A net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11666__A1 net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07878_ net719 _02828_ net877 vssd1 vssd1 vccd1 vccd1 _02829_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_39_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07381__A _02325_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07965__S0 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09617_ _04066_ _04108_ _04117_ vssd1 vssd1 vccd1 vccd1 _04536_ sky130_fd_sc_hd__o21ai_1
XANTENNA__11615__B net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06829_ final_design.cpu.reg_window\[597\] final_design.cpu.reg_window\[629\] net940
+ vssd1 vssd1 vccd1 vccd1 _01780_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout924_A net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout545_X net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11418__A1 net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09548_ net319 _04373_ _04376_ net320 _04466_ vssd1 vssd1 vccd1 vccd1 _04467_ sky130_fd_sc_hd__a221o_1
XFILLER_0_6_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11969__A2 net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09479_ _04396_ _04397_ net475 vssd1 vssd1 vccd1 vccd1 _04398_ sky130_fd_sc_hd__mux2_2
XANTENNA_fanout712_X net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11631__A net209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11510_ net1973 net220 net521 vssd1 vssd1 vccd1 vccd1 _00379_ sky130_fd_sc_hd__mux2_1
X_12490_ _06150_ net352 net332 net2025 vssd1 vssd1 vccd1 vccd1 _01196_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_43_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11441_ net2349 net177 net312 vssd1 vssd1 vccd1 vccd1 _00338_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_43_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08598__A1 net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14160_ clknet_leaf_19_clk _01334_ net1110 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.data_to_VGA\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09795__B1 _04348_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11372_ net589 _06058_ _06059_ vssd1 vssd1 vccd1 vccd1 _06060_ sky130_fd_sc_hd__and3_2
X_13111_ clknet_leaf_6_clk _00342_ net1128 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[99\]
+ sky130_fd_sc_hd__dfrtp_1
X_10323_ net1650 net1009 net986 final_design.data_from_mem\[8\] vssd1 vssd1 vccd1
+ vccd1 _00080_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14091_ clknet_leaf_19_clk _01288_ net1161 vssd1 vssd1 vccd1 vccd1 final_design.reqhand.instruction\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_46_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09547__B1 _04116_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input53_A mem_adr_start[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13042_ clknet_leaf_39_clk _00273_ net1209 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_10254_ final_design.uart.BAUD_counter\[19\] final_design.uart.BAUD_counter\[18\]
+ _05118_ final_design.uart.BAUD_counter\[20\] vssd1 vssd1 vccd1 vccd1 _05122_ sky130_fd_sc_hd__a31o_1
XANTENNA__08445__S1 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11354__B1 _05143_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1201 net1204 vssd1 vssd1 vccd1 vccd1 net1201 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_37_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1212 net1227 vssd1 vssd1 vccd1 vccd1 net1212 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_37_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10185_ final_design.uart.BAUD_counter\[9\] final_design.uart.BAUD_counter\[8\] final_design.uart.BAUD_counter\[11\]
+ final_design.uart.BAUD_counter\[10\] vssd1 vssd1 vccd1 vccd1 _05075_ sky130_fd_sc_hd__or4b_1
Xfanout1223 net1226 vssd1 vssd1 vccd1 vccd1 net1223 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_33_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11087__A1_N net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1870 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1234 net1235 vssd1 vssd1 vccd1 vccd1 net1234 sky130_fd_sc_hd__clkbuf_4
Xfanout1245 net100 vssd1 vssd1 vccd1 vccd1 net1245 sky130_fd_sc_hd__buf_4
Xfanout280 net281 vssd1 vssd1 vccd1 vccd1 net280 sky130_fd_sc_hd__clkbuf_4
Xfanout291 net293 vssd1 vssd1 vccd1 vccd1 net291 sky130_fd_sc_hd__clkbuf_4
XANTENNA__13645__CLK clknet_leaf_48_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13944_ clknet_leaf_64_clk _01175_ net1074 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[932\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_1917 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13875_ clknet_leaf_36_clk _01106_ net1210 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[863\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_1152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12826_ net1352 vssd1 vssd1 vccd1 vccd1 _00267_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_57_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13795__CLK clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12757_ _06392_ _06393_ vssd1 vssd1 vccd1 vccd1 _06394_ sky130_fd_sc_hd__or2_1
XANTENNA__12196__X _06271_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08825__A2 _01570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07184__S1 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11708_ net572 net424 _06212_ net297 net1900 vssd1 vssd1 vccd1 vccd1 _00485_ sky130_fd_sc_hd__a32o_1
XANTENNA__06836__A1 final_design.data_from_mem\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12688_ _06331_ net1390 net981 vssd1 vssd1 vccd1 vccd1 _01346_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11639_ net204 net633 vssd1 vssd1 vccd1 vccd1 _06177_ sky130_fd_sc_hd__and2_1
XANTENNA__13025__CLK clknet_leaf_47_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12794__25 clknet_leaf_31_clk vssd1 vssd1 vccd1 vccd1 net1335 sky130_fd_sc_hd__inv_2
XFILLER_0_68_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_3_clk_A clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold706 final_design.reqhand.data_from_UART\[1\] vssd1 vssd1 vccd1 vccd1 net2048
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11593__B1 net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold717 final_design.cpu.reg_window\[592\] vssd1 vssd1 vccd1 vccd1 net2059 sky130_fd_sc_hd__dlygate4sd3_1
X_13309_ clknet_leaf_2_clk _00540_ net1078 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[297\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold728 final_design.cpu.reg_window\[390\] vssd1 vssd1 vccd1 vccd1 net2070 sky130_fd_sc_hd__dlygate4sd3_1
Xhold739 final_design.cpu.reg_window\[928\] vssd1 vssd1 vccd1 vccd1 net2081 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09538__A0 net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13175__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11345__B1 _06035_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08850_ final_design.CPU_instr_adr\[29\] _03800_ vssd1 vssd1 vccd1 vccd1 _03801_
+ sky130_fd_sc_hd__and2_1
X_07801_ final_design.cpu.reg_window\[857\] final_design.cpu.reg_window\[889\] net853
+ vssd1 vssd1 vccd1 vccd1 _02752_ sky130_fd_sc_hd__mux2_1
X_08781_ _03692_ _03694_ _03729_ _03690_ _03689_ vssd1 vssd1 vccd1 vccd1 _03732_ sky130_fd_sc_hd__a311o_1
XFILLER_0_58_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07732_ final_design.cpu.reg_window\[154\] final_design.cpu.reg_window\[186\] net861
+ vssd1 vssd1 vccd1 vccd1 _02683_ sky130_fd_sc_hd__mux2_1
XANTENNA__11648__A1 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12311__S net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07913__B _02863_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09710__B1 net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07663_ final_design.cpu.reg_window\[478\] final_design.cpu.reg_window\[510\] net853
+ vssd1 vssd1 vccd1 vccd1 _02614_ sky130_fd_sc_hd__mux2_1
X_09402_ _04051_ _04291_ _04292_ _04320_ vssd1 vssd1 vccd1 vccd1 _04321_ sky130_fd_sc_hd__o31a_1
X_06614_ net763 _01564_ vssd1 vssd1 vccd1 vccd1 _01565_ sky130_fd_sc_hd__or2_1
XFILLER_0_18_1861 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07594_ _02543_ _02544_ vssd1 vssd1 vccd1 vccd1 _02545_ sky130_fd_sc_hd__or2_4
XANTENNA__09069__A2 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09333_ _04251_ vssd1 vssd1 vccd1 vccd1 _04252_ sky130_fd_sc_hd__inv_2
X_06545_ _01489_ net731 _01495_ vssd1 vssd1 vccd1 vccd1 _01496_ sky130_fd_sc_hd__and3_1
XANTENNA__12936__RESET_B net1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout240_A _05890_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08744__B net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout338_A net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09264_ net69 _04182_ net70 vssd1 vssd1 vccd1 vccd1 _04183_ sky130_fd_sc_hd__a21o_1
XFILLER_0_1_1414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06476_ final_design.data_from_mem\[18\] net969 _01425_ vssd1 vssd1 vccd1 vccd1 _01427_
+ sky130_fd_sc_hd__o21ai_4
XFILLER_0_69_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06922__S1 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08215_ _03132_ _03133_ _03162_ _03163_ vssd1 vssd1 vccd1 vccd1 _03166_ sky130_fd_sc_hd__o22a_1
X_09195_ _02543_ net442 _04113_ net527 vssd1 vssd1 vccd1 vccd1 _04114_ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout505_A net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08146_ net599 _03096_ vssd1 vssd1 vccd1 vccd1 _03097_ sky130_fd_sc_hd__or2_1
XANTENNA__13518__CLK clknet_leaf_43_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06686__S0 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08077_ _03025_ _03027_ vssd1 vssd1 vccd1 vccd1 _03028_ sky130_fd_sc_hd__nor2_1
XANTENNA__09792__A3 net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1035_X net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07028_ final_design.cpu.reg_window\[14\] final_design.cpu.reg_window\[46\] net893
+ vssd1 vssd1 vccd1 vccd1 _01979_ sky130_fd_sc_hd__mux2_1
XANTENNA__07376__A final_design.data_from_mem\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11336__B1 net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout495_X net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout874_A net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13668__CLK clknet_leaf_54_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold11 final_design.cpu.reg_window\[30\] vssd1 vssd1 vccd1 vccd1 net1353 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09591__A net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold22 final_design.cpu.reg_window\[23\] vssd1 vssd1 vccd1 vccd1 net1364 sky130_fd_sc_hd__dlygate4sd3_1
Xhold33 final_design.cpu.reg_window\[7\] vssd1 vssd1 vccd1 vccd1 net1375 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_51_1941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08979_ net625 _03914_ _03915_ vssd1 vssd1 vccd1 vccd1 _03916_ sky130_fd_sc_hd__a21o_1
Xhold44 final_design.cpu.reg_window\[1\] vssd1 vssd1 vccd1 vccd1 net1386 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_51_1952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout662_X net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold55 net115 vssd1 vssd1 vccd1 vccd1 net1397 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_51_1963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold66 net134 vssd1 vssd1 vccd1 vccd1 net1408 sky130_fd_sc_hd__dlygate4sd3_1
Xhold77 final_design.VGA_data_control.data_to_VGA\[3\] vssd1 vssd1 vccd1 vccd1 net1419
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold88 net163 vssd1 vssd1 vccd1 vccd1 net1430 sky130_fd_sc_hd__dlygate4sd3_1
X_11990_ net673 _06118_ _06193_ vssd1 vssd1 vccd1 vccd1 _06257_ sky130_fd_sc_hd__or3_4
Xhold99 final_design.cpu.reg_window\[218\] vssd1 vssd1 vccd1 vccd1 net1441 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10941_ _05662_ _05643_ vssd1 vssd1 vccd1 vccd1 _05669_ sky130_fd_sc_hd__nand2b_1
XANTENNA_fanout927_X net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06439__B net34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13660_ clknet_leaf_3_clk _00891_ net1065 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[648\]
+ sky130_fd_sc_hd__dfrtp_1
X_10872_ _05560_ _05578_ _05603_ _05563_ _05580_ vssd1 vssd1 vccd1 vccd1 _05604_ sky130_fd_sc_hd__o221a_1
XFILLER_0_71_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_1870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_1881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12611_ net1472 net999 net985 final_design.data_from_mem\[29\] vssd1 vssd1 vccd1
+ vccd1 _01304_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_26_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1885 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13048__CLK clknet_leaf_62_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13591_ clknet_leaf_4_clk _00822_ net1084 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[579\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_45_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08363__S0 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12542_ _06205_ net347 net323 net2222 vssd1 vssd1 vccd1 vccd1 _01246_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_41_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12473_ _06133_ net344 net330 net2172 vssd1 vssd1 vccd1 vccd1 _01179_ sky130_fd_sc_hd__a22o_1
XFILLER_0_81_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14212_ net1270 vssd1 vssd1 vccd1 vccd1 gpio_oeb[24] sky130_fd_sc_hd__buf_2
XANTENNA__13198__CLK clknet_leaf_45_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11424_ net2085 net208 net310 vssd1 vssd1 vccd1 vccd1 _00321_ sky130_fd_sc_hd__mux2_1
XANTENNA__09766__A net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10378__B2 final_design.data_from_mem\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11575__B1 net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_8 _06228_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14143_ clknet_leaf_19_clk _01317_ net1157 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.data_to_VGA\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_39_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11355_ _06041_ _06043_ _06044_ net589 vssd1 vssd1 vccd1 vccd1 _06045_ sky130_fd_sc_hd__o211a_1
XANTENNA__10705__A _04632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_1066 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10306_ final_design.VGA_data_control.data_to_VGA\[27\] final_design.VGA_data_control.data_to_VGA\[26\]
+ final_design.VGA_data_control.data_to_VGA\[25\] final_design.VGA_data_control.data_to_VGA\[24\]
+ net1050 net1049 vssd1 vssd1 vccd1 vccd1 _05160_ sky130_fd_sc_hd__mux4_1
XFILLER_0_21_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14074_ clknet_leaf_14_clk _01271_ net1107 vssd1 vssd1 vccd1 vccd1 final_design.uart.working_data\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_11286_ final_design.data_from_mem\[17\] net235 net233 vssd1 vssd1 vccd1 vccd1 _05984_
+ sky130_fd_sc_hd__a21o_2
XANTENNA__14180__Q final_design.VGA_adr\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13025_ clknet_leaf_47_clk _00256_ net1198 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_10237_ net1505 _05109_ _05111_ vssd1 vssd1 vccd1 vccd1 _00010_ sky130_fd_sc_hd__a21oi_1
Xfanout1020 _06298_ vssd1 vssd1 vccd1 vccd1 net1020 sky130_fd_sc_hd__clkbuf_2
Xfanout1031 net1036 vssd1 vssd1 vccd1 vccd1 net1031 sky130_fd_sc_hd__clkbuf_2
X_14193__1310 vssd1 vssd1 vccd1 vccd1 net1310 _14193__1310/LO sky130_fd_sc_hd__conb_1
Xfanout1042 _01371_ vssd1 vssd1 vccd1 vccd1 net1042 sky130_fd_sc_hd__clkbuf_8
XANTENNA__09940__B1 _04046_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10168_ _05041_ _05060_ vssd1 vssd1 vccd1 vccd1 final_design.vga.h_next_count\[8\]
+ sky130_fd_sc_hd__nor2_1
Xfanout1053 net1056 vssd1 vssd1 vccd1 vccd1 net1053 sky130_fd_sc_hd__clkbuf_4
Xfanout1064 net1069 vssd1 vssd1 vccd1 vccd1 net1064 sky130_fd_sc_hd__clkbuf_4
Xfanout1075 net1076 vssd1 vssd1 vccd1 vccd1 net1075 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08829__B _02504_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1086 net1117 vssd1 vssd1 vccd1 vccd1 net1086 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12131__S net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1097 net1098 vssd1 vssd1 vccd1 vccd1 net1097 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10440__A _02830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10099_ _05011_ _05014_ vssd1 vssd1 vccd1 vccd1 _05015_ sky130_fd_sc_hd__or2_1
XFILLER_0_76_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07929__S0 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13927_ clknet_leaf_62_clk _01158_ net1124 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[915\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_77_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06601__S0 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13858_ clknet_leaf_4_clk _01089_ net1083 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[846\]
+ sky130_fd_sc_hd__dfrtp_1
X_12809_ net1375 vssd1 vssd1 vccd1 vccd1 _00250_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_50_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09456__C1 net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13789_ clknet_leaf_1_clk _01020_ net1078 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[777\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08056__S net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_2281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_1745 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_2292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_1789 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08000_ final_design.cpu.reg_window\[784\] final_design.cpu.reg_window\[816\] net843
+ vssd1 vssd1 vccd1 vccd1 _02951_ sky130_fd_sc_hd__mux2_1
XANTENNA__12358__A2 net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10369__B2 final_design.data_from_mem\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold503 final_design.cpu.reg_window\[854\] vssd1 vssd1 vccd1 vccd1 net1845 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07234__A1 net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold514 final_design.cpu.reg_window\[237\] vssd1 vssd1 vccd1 vccd1 net1856 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12306__S net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold525 final_design.cpu.reg_window\[748\] vssd1 vssd1 vccd1 vccd1 net1867 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10615__A net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold536 final_design.cpu.reg_window\[188\] vssd1 vssd1 vccd1 vccd1 net1878 sky130_fd_sc_hd__dlygate4sd3_1
Xhold547 final_design.cpu.reg_window\[233\] vssd1 vssd1 vccd1 vccd1 net1889 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13810__CLK clknet_leaf_44_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07785__A2 _02731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold558 final_design.cpu.reg_window\[242\] vssd1 vssd1 vccd1 vccd1 net1900 sky130_fd_sc_hd__dlygate4sd3_1
X_09951_ _04091_ _04436_ _04446_ net494 vssd1 vssd1 vccd1 vccd1 _04870_ sky130_fd_sc_hd__a31oi_2
XFILLER_0_60_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold569 final_design.uart.BAUD_counter\[28\] vssd1 vssd1 vccd1 vccd1 net1911 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_55_2074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_2085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkload25_A clknet_leaf_25_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08902_ _03771_ _03846_ vssd1 vssd1 vccd1 vccd1 _03847_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_55_2096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09882_ net483 _04733_ _04799_ _04800_ vssd1 vssd1 vccd1 vccd1 _04801_ sky130_fd_sc_hd__o22a_1
XANTENNA__11149__C _05862_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08833_ final_design.CPU_instr_adr\[4\] final_design.CPU_instr_adr\[3\] net1018 vssd1
+ vssd1 vccd1 vccd1 _03784_ sky130_fd_sc_hd__and3_1
XANTENNA__07924__A net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1203 final_design.cpu.reg_window\[52\] vssd1 vssd1 vccd1 vccd1 net2545 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1214 final_design.cpu.reg_window\[420\] vssd1 vssd1 vccd1 vccd1 net2556 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout190_A _06038_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13960__CLK clknet_leaf_41_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout288_A net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12041__S net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08764_ final_design.CPU_instr_adr\[0\] _02425_ vssd1 vssd1 vccd1 vccd1 _03715_ sky130_fd_sc_hd__and2_1
XANTENNA__07135__S net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07715_ _02662_ _02663_ _02664_ _02665_ net686 net704 vssd1 vssd1 vccd1 vccd1 _02666_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_0_211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12294__A1 net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08695_ _01998_ _02028_ vssd1 vssd1 vccd1 vccd1 _03646_ sky130_fd_sc_hd__nand2_2
XFILLER_0_75_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1612 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1197_A net1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07646_ final_design.cpu.reg_window\[668\] final_design.cpu.reg_window\[700\] net866
+ vssd1 vssd1 vccd1 vccd1 _02597_ sky130_fd_sc_hd__mux2_1
XANTENNA__10349__X _05170_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07577_ final_design.cpu.reg_window\[607\] final_design.cpu.reg_window\[639\] net857
+ vssd1 vssd1 vccd1 vccd1 _02528_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout622_A _02506_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10057__B1 _04954_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09316_ net532 net530 net529 _02325_ net456 net465 vssd1 vssd1 vccd1 vccd1 _04235_
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_48_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06528_ net1041 net993 net990 _01378_ vssd1 vssd1 vccd1 vccd1 _01479_ sky130_fd_sc_hd__a31o_1
XANTENNA__11254__C1 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1211 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13340__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1244 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09247_ _02673_ _02705_ _02738_ _02770_ vssd1 vssd1 vccd1 vccd1 _04166_ sky130_fd_sc_hd__or4_1
X_06459_ net1053 net1037 vssd1 vssd1 vccd1 vccd1 _01412_ sky130_fd_sc_hd__or2_1
XFILLER_0_7_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout410_X net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1891 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12908__CLK clknet_leaf_61_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout508_X net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12349__A2 net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09178_ net489 _03629_ net659 vssd1 vssd1 vccd1 vccd1 _04097_ sky130_fd_sc_hd__or3_4
XANTENNA__11557__B1 net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08129_ final_design.cpu.reg_window\[205\] final_design.cpu.reg_window\[237\] net850
+ vssd1 vssd1 vccd1 vccd1 _03080_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_63_clk_X clknet_leaf_63_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13490__CLK clknet_leaf_39_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11140_ net645 _05854_ vssd1 vssd1 vccd1 vccd1 _05855_ sky130_fd_sc_hd__and2_2
XFILLER_0_43_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11309__B1 net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout877_X net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11071_ _05757_ _05775_ _05792_ vssd1 vssd1 vccd1 vccd1 _05794_ sky130_fd_sc_hd__or3_1
X_10022_ net68 _04940_ vssd1 vssd1 vccd1 vccd1 _04941_ sky130_fd_sc_hd__nand2_1
XANTENNA__12521__A2 net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10532__A1 net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10532__B2 net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11356__A net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06831__S0 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input16_A DAT_I[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11973_ _06175_ net276 net404 net1586 vssd1 vssd1 vccd1 vccd1 _00706_ sky130_fd_sc_hd__a22o_1
XANTENNA__12285__A1 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_47_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10924_ net82 net1046 net83 vssd1 vssd1 vccd1 vccd1 _05653_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_47_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13712_ clknet_leaf_36_clk _00943_ net1237 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[700\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_47_1829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08665__A _01999_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10855_ _05549_ _05570_ vssd1 vssd1 vccd1 vccd1 _05587_ sky130_fd_sc_hd__nor2_1
X_13643_ clknet_leaf_52_clk _00874_ net1183 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[631\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_16_clk_X clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12588__A2 net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11245__C1 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13574_ clknet_leaf_51_clk _00805_ net1169 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[562\]
+ sky130_fd_sc_hd__dfrtp_1
X_10786_ net43 _05521_ vssd1 vssd1 vccd1 vccd1 _05522_ sky130_fd_sc_hd__and2_1
XANTENNA__09453__A2 _04342_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10419__B _05190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12525_ _06187_ net355 net328 net1730 vssd1 vssd1 vccd1 vccd1 _01230_ sky130_fd_sc_hd__a22o_1
XFILLER_0_32_1699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08661__B1 _02542_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13833__CLK clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12456_ net1875 net191 net337 vssd1 vssd1 vccd1 vccd1 _01163_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_10_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12771__2_A clknet_leaf_25_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11407_ net437 net579 _06090_ net316 net1722 vssd1 vssd1 vccd1 vccd1 _00306_ sky130_fd_sc_hd__a32o_1
X_12387_ net1725 net193 net270 vssd1 vssd1 vccd1 vccd1 _01098_ sky130_fd_sc_hd__mux2_1
XANTENNA__12126__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14126_ clknet_leaf_20_clk final_design.vga.v_next_count\[6\] net1160 vssd1 vssd1
+ vccd1 vccd1 final_design.VGA_data_control.v_count\[6\] sky130_fd_sc_hd__dfrtp_2
X_11338_ _04546_ _04549_ net652 vssd1 vssd1 vccd1 vccd1 _06030_ sky130_fd_sc_hd__a21o_1
XFILLER_0_61_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13983__CLK clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14057_ clknet_leaf_16_clk _00019_ net1091 vssd1 vssd1 vccd1 vccd1 final_design.uart.BAUD_counter\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_11269_ net738 _03930_ vssd1 vssd1 vccd1 vccd1 _05969_ sky130_fd_sc_hd__nand2_1
X_13008_ net1339 _00239_ net1234 vssd1 vssd1 vccd1 vccd1 final_design.CPU_instr_adr\[28\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__12512__A2 net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11720__B1 net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13213__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12276__A1 net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07500_ _02002_ _02450_ vssd1 vssd1 vccd1 vccd1 _02451_ sky130_fd_sc_hd__nor2_1
X_08480_ _03427_ _03428_ _03429_ _03430_ net677 net699 vssd1 vssd1 vccd1 vccd1 _03431_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__06647__X _01598_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_2490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13363__CLK clknet_leaf_40_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire211_X net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_2343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12028__A1 net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07431_ net752 _02381_ vssd1 vssd1 vccd1 vccd1 _02382_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_63_2354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11272__Y _05972_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11713__B net196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_2988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_2365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1875 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07362_ final_design.cpu.reg_window\[835\] final_design.cpu.reg_window\[867\] net912
+ vssd1 vssd1 vccd1 vccd1 _02313_ sky130_fd_sc_hd__mux2_1
XANTENNA__11787__B1 net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09101_ final_design.CPU_instr_adr\[3\] _04023_ net1037 vssd1 vssd1 vccd1 vccd1 _00214_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07293_ final_design.cpu.reg_window\[5\] final_design.cpu.reg_window\[37\] net921
+ vssd1 vssd1 vccd1 vccd1 _02244_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09032_ _03960_ _03962_ net620 vssd1 vssd1 vccd1 vccd1 _03963_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11539__A0 net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold300 final_design.cpu.reg_window\[725\] vssd1 vssd1 vccd1 vccd1 net1642 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_2147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold311 final_design.cpu.reg_window\[162\] vssd1 vssd1 vccd1 vccd1 net1653 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12036__S net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_2158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout203_A _05989_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold322 final_design.cpu.reg_window\[742\] vssd1 vssd1 vccd1 vccd1 net1664 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_2169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold333 final_design.cpu.reg_window\[859\] vssd1 vssd1 vccd1 vccd1 net1675 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07302__S1 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold344 final_design.cpu.reg_window\[182\] vssd1 vssd1 vccd1 vccd1 net1686 sky130_fd_sc_hd__dlygate4sd3_1
Xhold355 final_design.cpu.reg_window\[255\] vssd1 vssd1 vccd1 vccd1 net1697 sky130_fd_sc_hd__dlygate4sd3_1
Xhold366 final_design.cpu.reg_window\[908\] vssd1 vssd1 vccd1 vccd1 net1708 sky130_fd_sc_hd__dlygate4sd3_1
Xhold377 final_design.cpu.reg_window\[530\] vssd1 vssd1 vccd1 vccd1 net1719 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout802 _04039_ vssd1 vssd1 vccd1 vccd1 net802 sky130_fd_sc_hd__buf_4
Xhold388 final_design.cpu.reg_window\[987\] vssd1 vssd1 vccd1 vccd1 net1730 sky130_fd_sc_hd__dlygate4sd3_1
Xhold399 final_design.cpu.reg_window\[231\] vssd1 vssd1 vccd1 vccd1 net1741 sky130_fd_sc_hd__dlygate4sd3_1
X_09934_ net470 _04732_ net482 vssd1 vssd1 vccd1 vccd1 _04853_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout1112_A net1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout813 net815 vssd1 vssd1 vccd1 vccd1 net813 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_61_1873 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout824 net829 vssd1 vssd1 vccd1 vccd1 net824 sky130_fd_sc_hd__buf_2
XANTENNA__09345__S net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout835 net842 vssd1 vssd1 vccd1 vccd1 net835 sky130_fd_sc_hd__clkbuf_4
Xfanout846 net847 vssd1 vssd1 vccd1 vccd1 net846 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12503__A2 net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09904__B1 net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input8_A DAT_I[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout857 net860 vssd1 vssd1 vccd1 vccd1 net857 sky130_fd_sc_hd__clkbuf_4
X_09865_ _04781_ _04783_ net497 vssd1 vssd1 vccd1 vccd1 _04784_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_42_1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1000 final_design.cpu.reg_window\[60\] vssd1 vssd1 vccd1 vccd1 net2342 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_1879 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout572_A net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout868 net871 vssd1 vssd1 vccd1 vccd1 net868 sky130_fd_sc_hd__clkbuf_4
Xhold1011 net154 vssd1 vssd1 vccd1 vccd1 net2353 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout879 _01687_ vssd1 vssd1 vccd1 vccd1 net879 sky130_fd_sc_hd__buf_4
XANTENNA__09380__A1 net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1022 final_design.cpu.reg_window\[907\] vssd1 vssd1 vccd1 vccd1 net2364 sky130_fd_sc_hd__dlygate4sd3_1
X_08816_ _03759_ _03761_ _03764_ _03766_ vssd1 vssd1 vccd1 vccd1 _03767_ sky130_fd_sc_hd__a31o_1
Xhold1033 final_design.cpu.reg_window\[433\] vssd1 vssd1 vccd1 vccd1 net2375 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06813__S0 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11607__C net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1044 final_design.cpu.reg_window\[414\] vssd1 vssd1 vccd1 vccd1 net2386 sky130_fd_sc_hd__dlygate4sd3_1
X_09796_ _03357_ net441 net438 _03356_ vssd1 vssd1 vccd1 vccd1 _04715_ sky130_fd_sc_hd__o22a_1
XFILLER_0_38_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1055 final_design.cpu.reg_window\[295\] vssd1 vssd1 vccd1 vccd1 net2397 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1066 final_design.cpu.reg_window\[614\] vssd1 vssd1 vccd1 vccd1 net2408 sky130_fd_sc_hd__dlygate4sd3_1
X_08747_ net666 _01598_ final_design.CPU_instr_adr\[7\] vssd1 vssd1 vccd1 vccd1 _03698_
+ sky130_fd_sc_hd__a21o_1
XANTENNA__13706__CLK clknet_leaf_60_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1077 final_design.cpu.reg_window\[564\] vssd1 vssd1 vccd1 vccd1 net2419 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12951__RESET_B net1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1088 final_design.cpu.reg_window\[945\] vssd1 vssd1 vccd1 vccd1 net2430 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout360_X net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1099 final_design.uart.BAUD_counter\[7\] vssd1 vssd1 vccd1 vccd1 net2441 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14175__RESET_B net1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout837_A net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08678_ _03617_ net594 vssd1 vssd1 vccd1 vccd1 _03629_ sky130_fd_sc_hd__or2_2
XFILLER_0_16_1628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09683__A2 _04087_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11623__B net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07629_ final_design.cpu.reg_window\[476\] final_design.cpu.reg_window\[508\] net858
+ vssd1 vssd1 vccd1 vccd1 _02580_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout625_X net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13856__CLK clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10640_ net67 _05382_ vssd1 vssd1 vccd1 vccd1 _05383_ sky130_fd_sc_hd__xor2_1
XANTENNA__11778__B1 net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10571_ _05291_ _05294_ _05316_ vssd1 vssd1 vccd1 vccd1 _05317_ sky130_fd_sc_hd__or3_1
XANTENNA__11192__A_N final_design.reqhand.data_from_UART\[6\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_12310_ net2112 net210 net367 vssd1 vssd1 vccd1 vccd1 _01024_ sky130_fd_sc_hd__mux2_1
X_13290_ clknet_leaf_59_clk _00521_ net1170 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[278\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12880__CLK clknet_leaf_18_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12241_ net568 _06171_ net507 net373 net1489 vssd1 vssd1 vccd1 vccd1 _00958_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_20_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_903 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06452__B net1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07749__A2 _02698_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12172_ net1793 net221 net380 vssd1 vssd1 vccd1 vccd1 _00891_ sky130_fd_sc_hd__mux2_1
XANTENNA__11950__B1 net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11123_ net805 _02392_ vssd1 vssd1 vccd1 vccd1 _05838_ sky130_fd_sc_hd__or2_2
XANTENNA_clkbuf_leaf_43_clk_A clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1913 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07564__A _02504_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11054_ _05776_ _05777_ net1452 net1034 vssd1 vssd1 vccd1 vccd1 _00201_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__06709__B1 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11702__B1 net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10005_ _04703_ _04885_ _04906_ _04923_ vssd1 vssd1 vccd1 vccd1 _04924_ sky130_fd_sc_hd__and4_1
XFILLER_0_64_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13386__CLK clknet_leaf_51_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_58_clk_A clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11956_ net568 _06118_ _06158_ vssd1 vssd1 vccd1 vccd1 _06255_ sky130_fd_sc_hd__or3_4
XANTENNA__06467__X _01418_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10907_ final_design.CPU_instr_adr\[22\] _03879_ net1059 vssd1 vssd1 vccd1 vccd1
+ _05637_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_17_Left_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08882__B1 net1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11887_ _05875_ net2280 net273 vssd1 vssd1 vccd1 vccd1 _00629_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10838_ _05549_ _05551_ vssd1 vssd1 vccd1 vccd1 _05571_ sky130_fd_sc_hd__nand2_1
XFILLER_0_67_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13626_ clknet_leaf_64_clk _00857_ net1075 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[614\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_13_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09426__A2 net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10769_ _05497_ _05503_ _05504_ vssd1 vssd1 vccd1 vccd1 _05505_ sky130_fd_sc_hd__or3_1
XFILLER_0_3_1873 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13557_ clknet_leaf_57_clk _00788_ net1133 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[545\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12508_ _06170_ net344 net326 net1572 vssd1 vssd1 vccd1 vccd1 _01213_ sky130_fd_sc_hd__a22o_1
X_13488_ clknet_leaf_36_clk _00719_ net1236 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[476\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12439_ net1815 net244 net334 vssd1 vssd1 vccd1 vccd1 _01146_ sky130_fd_sc_hd__mux2_1
XANTENNA__10165__A _05058_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_75_2770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_2781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07296__S0 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_2623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_2000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_2634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_71_2645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11941__B1 net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14109_ clknet_leaf_24_clk _01306_ net1163 vssd1 vssd1 vccd1 vccd1 final_design.reqhand.instruction\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14161__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07980_ _01909_ net613 vssd1 vssd1 vccd1 vccd1 _02931_ sky130_fd_sc_hd__nor2_1
XFILLER_0_38_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06931_ net546 _01881_ vssd1 vssd1 vccd1 vccd1 _01882_ sky130_fd_sc_hd__and2b_1
XANTENNA__13729__CLK clknet_leaf_47_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09362__A1 _04158_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09650_ _04567_ _04568_ vssd1 vssd1 vccd1 vccd1 _04569_ sky130_fd_sc_hd__or2_1
X_06862_ _01809_ _01810_ _01811_ _01812_ net776 net783 vssd1 vssd1 vccd1 vccd1 _01813_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_78_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_2552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08601_ net614 _03550_ _02423_ vssd1 vssd1 vccd1 vccd1 _03552_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_69_2563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12249__A1 net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09581_ _03134_ _03582_ _04499_ vssd1 vssd1 vccd1 vccd1 _04500_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_69_2574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06793_ final_design.cpu.reg_window\[854\] final_design.cpu.reg_window\[886\] net918
+ vssd1 vssd1 vccd1 vccd1 _01744_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_65_2416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_2427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_2438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13879__CLK clknet_leaf_58_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08532_ _02361_ net609 vssd1 vssd1 vccd1 vccd1 _03483_ sky130_fd_sc_hd__or2_1
XFILLER_0_78_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_1374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08463_ _03408_ _03413_ net707 vssd1 vssd1 vccd1 vccd1 _03414_ sky130_fd_sc_hd__mux2_1
XANTENNA__11443__B net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07414_ final_design.cpu.reg_window\[321\] final_design.cpu.reg_window\[353\] net922
+ vssd1 vssd1 vccd1 vccd1 _02365_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_50 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08394_ _03341_ _03342_ _03343_ _03344_ net679 net699 vssd1 vssd1 vccd1 vccd1 _03345_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__13109__CLK clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09417__A2 _01596_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07345_ _01484_ _02295_ vssd1 vssd1 vccd1 vccd1 _02296_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout320_A _04073_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_2209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_30_clk clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_30_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout418_A net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1062_A net1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09200__Y _04119_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07276_ net759 _02226_ net745 vssd1 vssd1 vccd1 vccd1 _02227_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_72_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09015_ net623 _03947_ _03946_ net255 vssd1 vssd1 vccd1 vccd1 _03948_ sky130_fd_sc_hd__a211o_1
XANTENNA__13259__CLK clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout206_X net206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12185__B1 _06270_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08928__A1 net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold130 final_design.reqhand.instruction\[29\] vssd1 vssd1 vccd1 vccd1 net1472 sky130_fd_sc_hd__dlygate4sd3_1
Xhold141 final_design.VGA_data_control.ready_data\[6\] vssd1 vssd1 vccd1 vccd1 net1483
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold152 final_design.VGA_data_control.ready_data\[22\] vssd1 vssd1 vccd1 vccd1 net1494
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10735__A1 net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10735__B2 _04042_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold163 final_design.uart.BAUD_counter\[13\] vssd1 vssd1 vccd1 vccd1 net1505 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11932__B1 net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout787_A net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold174 net153 vssd1 vssd1 vccd1 vccd1 net1516 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold185 final_design.VGA_data_control.data_to_VGA\[19\] vssd1 vssd1 vccd1 vccd1 net1527
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1115_X net1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold196 final_design.cpu.reg_window\[219\] vssd1 vssd1 vccd1 vccd1 net1538 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout610 net612 vssd1 vssd1 vccd1 vccd1 net610 sky130_fd_sc_hd__buf_2
Xfanout621 _02507_ vssd1 vssd1 vccd1 vccd1 net621 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11408__A_N net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09917_ net485 _04407_ _04835_ vssd1 vssd1 vccd1 vccd1 _04836_ sky130_fd_sc_hd__o21ai_2
Xfanout632 net633 vssd1 vssd1 vccd1 vccd1 net632 sky130_fd_sc_hd__buf_4
Xfanout643 net644 vssd1 vssd1 vccd1 vccd1 net643 sky130_fd_sc_hd__buf_2
XANTENNA_fanout954_A _05039_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout654 net655 vssd1 vssd1 vccd1 vccd1 net654 sky130_fd_sc_hd__buf_2
Xfanout665 _01503_ vssd1 vssd1 vccd1 vccd1 net665 sky130_fd_sc_hd__clkbuf_8
XANTENNA__10499__B1 net1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout676 net690 vssd1 vssd1 vccd1 vccd1 net676 sky130_fd_sc_hd__buf_4
X_09848_ net726 _04763_ _04765_ vssd1 vssd1 vccd1 vccd1 _04767_ sky130_fd_sc_hd__or3_1
Xfanout687 net688 vssd1 vssd1 vccd1 vccd1 net687 sky130_fd_sc_hd__buf_4
Xfanout698 net701 vssd1 vssd1 vccd1 vccd1 net698 sky130_fd_sc_hd__buf_4
XFILLER_0_77_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09779_ net75 _04186_ vssd1 vssd1 vccd1 vccd1 _04698_ sky130_fd_sc_hd__nand2_1
XANTENNA__10432__A_N net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11810_ _06091_ net281 vssd1 vssd1 vccd1 vccd1 _06237_ sky130_fd_sc_hd__nand2_1
XFILLER_0_55_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07323__S net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11999__B1 net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11741_ net224 net2477 net417 vssd1 vssd1 vccd1 vccd1 _00504_ sky130_fd_sc_hd__mux2_1
X_11672_ net232 net2299 net294 vssd1 vssd1 vccd1 vccd1 _00467_ sky130_fd_sc_hd__mux2_1
XANTENNA__14034__CLK clknet_leaf_39_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10623_ net1002 _05365_ _05366_ net1031 net1362 vssd1 vssd1 vccd1 vccd1 _00181_ sky130_fd_sc_hd__a32o_1
X_13411_ clknet_leaf_1_clk _00642_ net1072 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[399\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_12_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10018__A3 _04053_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_12_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_21_clk clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_21_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__08662__B _02029_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13342_ clknet_leaf_9_clk _00573_ net1103 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[330\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input83_A memory_size[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10554_ net668 _05287_ _05300_ net964 _05299_ vssd1 vssd1 vccd1 vccd1 _05301_ sky130_fd_sc_hd__o221a_1
XFILLER_0_68_1857 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13273_ clknet_leaf_55_clk _00504_ net1148 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[261\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14184__CLK clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10485_ net90 final_design.VGA_adr\[0\] vssd1 vssd1 vccd1 vccd1 _05235_ sky130_fd_sc_hd__nand2_1
XFILLER_0_49_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12224_ net585 _06152_ net512 net378 net1736 vssd1 vssd1 vccd1 vccd1 _00942_ sky130_fd_sc_hd__a32o_1
XANTENNA__07846__X _02797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11923__B1 net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09592__A1 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11368__X _06056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12155_ net188 net2305 net386 vssd1 vssd1 vccd1 vccd1 _00876_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11106_ _05819_ _05826_ vssd1 vssd1 vccd1 vccd1 _05827_ sky130_fd_sc_hd__nand2_1
X_12086_ net583 _06039_ net514 net395 net1937 vssd1 vssd1 vccd1 vccd1 _00811_ sky130_fd_sc_hd__a32o_1
XANTENNA__10432__B _02961_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11037_ net88 net1045 vssd1 vssd1 vccd1 vccd1 _05761_ sky130_fd_sc_hd__or2_1
XFILLER_0_75_1817 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12988_ net1319 _00219_ net1165 vssd1 vssd1 vccd1 vccd1 final_design.CPU_instr_adr\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06638__A net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07202__S0 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11939_ _06140_ net276 net408 net2298 vssd1 vssd1 vccd1 vccd1 _00674_ sky130_fd_sc_hd__a22o_1
XANTENNA__12651__B2 final_design.data_from_mem\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10594__S net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13609_ clknet_leaf_37_clk _00840_ net1228 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[597\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13401__CLK clknet_leaf_56_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_12_clk clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_12_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__08572__B net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07130_ final_design.cpu.reg_window\[779\] final_design.cpu.reg_window\[811\] net908
+ vssd1 vssd1 vccd1 vccd1 _02081_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_77_2821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1889 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_2832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_2843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07061_ final_design.cpu.reg_window\[141\] final_design.cpu.reg_window\[173\] net930
+ vssd1 vssd1 vccd1 vccd1 _02012_ sky130_fd_sc_hd__mux2_1
XFILLER_0_40_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_2707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07269__S0 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10717__A1 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13551__CLK clknet_leaf_39_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11278__X _05977_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09583__A1 net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12314__S net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11390__A1 net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire543_X net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07963_ final_design.cpu.reg_window\[209\] final_design.cpu.reg_window\[241\] net848
+ vssd1 vssd1 vccd1 vccd1 _02914_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06914_ final_design.cpu.reg_window\[210\] final_design.cpu.reg_window\[242\] net924
+ vssd1 vssd1 vccd1 vccd1 _01865_ sky130_fd_sc_hd__mux2_1
X_09702_ _04092_ _04312_ _04298_ vssd1 vssd1 vccd1 vccd1 _04621_ sky130_fd_sc_hd__o21ai_1
X_07894_ final_design.cpu.reg_window\[87\] final_design.cpu.reg_window\[119\] net849
+ vssd1 vssd1 vccd1 vccd1 _02845_ sky130_fd_sc_hd__mux2_1
XANTENNA__07346__B1 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09886__A2 _04793_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09633_ _04550_ _04551_ vssd1 vssd1 vccd1 vccd1 _04552_ sky130_fd_sc_hd__xor2_1
X_06845_ net754 _01795_ vssd1 vssd1 vccd1 vccd1 _01796_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout270_A net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout368_A net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09564_ _03132_ net443 net440 _03133_ vssd1 vssd1 vccd1 vccd1 _04483_ sky130_fd_sc_hd__a2bb2o_1
X_06776_ final_design.cpu.reg_window\[278\] final_design.cpu.reg_window\[310\] net920
+ vssd1 vssd1 vccd1 vccd1 _01727_ sky130_fd_sc_hd__mux2_1
XANTENNA__06548__A net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14057__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08515_ final_design.cpu.reg_window\[130\] final_design.cpu.reg_window\[162\] net837
+ vssd1 vssd1 vccd1 vccd1 _03466_ sky130_fd_sc_hd__mux2_1
X_09495_ _02607_ net443 net439 _02606_ _04413_ vssd1 vssd1 vccd1 vccd1 _04414_ sky130_fd_sc_hd__o221a_1
XFILLER_0_78_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout535_A net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08310__A2 _03257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08446_ final_design.cpu.reg_window\[68\] final_design.cpu.reg_window\[100\] net822
+ vssd1 vssd1 vccd1 vccd1 _03397_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_1923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08377_ _02240_ net597 vssd1 vssd1 vccd1 vccd1 _03328_ sky130_fd_sc_hd__nand2_1
XFILLER_0_50_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13081__CLK clknet_leaf_59_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout702_A _01752_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout323_X net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_983 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07328_ final_design.cpu.reg_window\[132\] final_design.cpu.reg_window\[164\] net902
+ vssd1 vssd1 vccd1 vccd1 _02279_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_22_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08074__A1 net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07259_ _02204_ _02209_ net749 vssd1 vssd1 vccd1 vccd1 _02210_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10270_ final_design.uart.BAUD_counter\[25\] final_design.uart.BAUD_counter\[24\]
+ _05128_ final_design.uart.BAUD_counter\[26\] vssd1 vssd1 vccd1 vccd1 _05132_ sky130_fd_sc_hd__a31o_1
XANTENNA__11905__A0 net197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout692_X net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10092__X _05008_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11629__A net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout440 _04094_ vssd1 vssd1 vccd1 vccd1 net440 sky130_fd_sc_hd__buf_4
XANTENNA_fanout957_X net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout451 _04069_ vssd1 vssd1 vccd1 vccd1 net451 sky130_fd_sc_hd__buf_1
Xfanout462 net463 vssd1 vssd1 vccd1 vccd1 net462 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_35_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13960_ clknet_leaf_41_clk _01191_ net1224 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[948\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout473 net474 vssd1 vssd1 vccd1 vccd1 net473 sky130_fd_sc_hd__buf_2
Xfanout484 net488 vssd1 vssd1 vccd1 vccd1 net484 sky130_fd_sc_hd__buf_2
Xfanout495 _03419_ vssd1 vssd1 vccd1 vccd1 net495 sky130_fd_sc_hd__buf_4
XANTENNA__12330__B1 net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12911_ clknet_leaf_61_clk _00149_ net1137 vssd1 vssd1 vccd1 vccd1 net164 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_31_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13891_ clknet_leaf_64_clk _01122_ net1075 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[879\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11684__A2 net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11364__A net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12842_ clknet_leaf_15_clk _00080_ net1094 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.ready_data\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06458__A net1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12633__B2 final_design.data_from_mem\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13424__CLK clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11724_ net581 net423 _06220_ net297 net1904 vssd1 vssd1 vccd1 vccd1 _00493_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_29_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08673__A _01999_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11655_ net189 net632 vssd1 vssd1 vccd1 vccd1 _06185_ sky130_fd_sc_hd__and2_1
XANTENNA__09488__B _04406_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12397__B1 net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10606_ net98 final_design.VGA_adr\[6\] vssd1 vssd1 vccd1 vccd1 _05350_ sky130_fd_sc_hd__or2_1
X_11586_ net190 net636 vssd1 vssd1 vccd1 vccd1 _06149_ sky130_fd_sc_hd__and2_1
XANTENNA__13574__CLK clknet_leaf_51_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10427__B _05190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14183__Q final_design.VGA_adr\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13001__RESET_B net1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10537_ _05283_ _05284_ vssd1 vssd1 vccd1 vccd1 _05285_ sky130_fd_sc_hd__nand2_1
X_13325_ clknet_leaf_44_clk _00556_ net1204 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[313\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07812__B2 net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10468_ net668 _05216_ _05219_ vssd1 vssd1 vccd1 vccd1 _05220_ sky130_fd_sc_hd__o21a_1
X_13256_ clknet_leaf_41_clk _00487_ net1220 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[244\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12207_ net560 _06135_ net503 net376 net1660 vssd1 vssd1 vccd1 vccd1 _00925_ sky130_fd_sc_hd__a32o_1
XANTENNA__12134__S net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13187_ clknet_leaf_0_clk _00418_ net1061 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[175\]
+ sky130_fd_sc_hd__dfrtp_1
X_10399_ net250 _05182_ net1027 net1408 vssd1 vssd1 vccd1 vccd1 _00141_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_23_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12138_ net220 net2466 net384 vssd1 vssd1 vccd1 vccd1 _00859_ sky130_fd_sc_hd__mux2_1
X_12069_ net558 _05911_ net502 net392 net2220 vssd1 vssd1 vccd1 vccd1 _00794_ sky130_fd_sc_hd__a32o_1
XFILLER_0_79_1761 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_1_clk clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_1_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_75_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07423__S0 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07879__A1 net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1024 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06630_ _01577_ _01578_ _01579_ _01580_ net775 net793 vssd1 vssd1 vccd1 vccd1 _01581_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__06551__A1 final_design.data_from_mem\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06561_ final_design.cpu.reg_window\[285\] final_design.cpu.reg_window\[317\] net950
+ vssd1 vssd1 vccd1 vccd1 _01512_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1721 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08300_ final_design.cpu.reg_window\[841\] final_design.cpu.reg_window\[873\] net820
+ vssd1 vssd1 vccd1 vccd1 _03251_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_16_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09280_ _02641_ _04172_ vssd1 vssd1 vccd1 vccd1 _04199_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_16_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06492_ final_design.cpu.reg_window\[926\] final_design.cpu.reg_window\[958\] net935
+ vssd1 vssd1 vccd1 vccd1 _01443_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_16_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08231_ final_design.cpu.reg_window\[779\] final_design.cpu.reg_window\[811\] net826
+ vssd1 vssd1 vccd1 vccd1 _03182_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_79_2905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11721__B net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13917__CLK clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_2916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12309__S net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08162_ final_design.cpu.reg_window\[207\] final_design.cpu.reg_window\[239\] net807
+ vssd1 vssd1 vccd1 vccd1 _03113_ sky130_fd_sc_hd__mux2_1
XANTENNA__10938__A1 net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07113_ net743 net667 _01851_ _02061_ _01821_ vssd1 vssd1 vccd1 vccd1 _02064_ sky130_fd_sc_hd__o221ai_4
X_08093_ final_design.cpu.reg_window\[460\] final_design.cpu.reg_window\[492\] net817
+ vssd1 vssd1 vccd1 vccd1 _03044_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12941__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07044_ net882 _01988_ _01994_ _01981_ _01982_ vssd1 vssd1 vccd1 vccd1 _01995_ sky130_fd_sc_hd__a32oi_4
XFILLER_0_62_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_284 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12044__S net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12560__B1 net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08995_ final_design.CPU_instr_adr\[15\] _03791_ vssd1 vssd1 vccd1 vccd1 _03930_
+ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout485_A net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07946_ net613 _02894_ _02895_ _01750_ vssd1 vssd1 vccd1 vccd1 _02897_ sky130_fd_sc_hd__a211oi_1
XANTENNA__09859__A2 net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11666__A2 net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07877_ _02824_ _02825_ _02826_ _02827_ net687 net694 vssd1 vssd1 vccd1 vccd1 _02828_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout273_X net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout652_A _05143_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13447__CLK clknet_leaf_63_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07965__S1 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09616_ _02867_ _04094_ vssd1 vssd1 vccd1 vccd1 _04535_ sky130_fd_sc_hd__nand2_1
X_06828_ final_design.cpu.reg_window\[661\] final_design.cpu.reg_window\[693\] net938
+ vssd1 vssd1 vccd1 vccd1 _01779_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_1889 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06759_ net756 _01709_ vssd1 vssd1 vccd1 vccd1 _01710_ sky130_fd_sc_hd__or2_1
X_09547_ net481 _04377_ _04116_ vssd1 vssd1 vccd1 vccd1 _04466_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout440_X net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout538_X net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout917_A net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09492__A0 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09478_ net465 _03639_ vssd1 vssd1 vccd1 vccd1 _04397_ sky130_fd_sc_hd__or2_1
XANTENNA__13597__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11631__B net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08429_ final_design.cpu.reg_window\[581\] final_design.cpu.reg_window\[613\] net840
+ vssd1 vssd1 vccd1 vccd1 _03380_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout705_X net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1106 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload0 clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 clkload0/X sky130_fd_sc_hd__clkbuf_8
X_11440_ net1712 net179 net313 vssd1 vssd1 vccd1 vccd1 _00337_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_43_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10929__A1 net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1805 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11371_ _04280_ _04285_ _05143_ vssd1 vssd1 vccd1 vccd1 _06059_ sky130_fd_sc_hd__a21o_1
XFILLER_0_65_1849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13110_ clknet_leaf_61_clk _00341_ net1136 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[98\]
+ sky130_fd_sc_hd__dfrtp_1
X_10322_ net1521 net1011 net988 final_design.data_from_mem\[7\] vssd1 vssd1 vccd1
+ vccd1 _00079_ sky130_fd_sc_hd__a22o_1
X_14090_ clknet_leaf_25_clk _01287_ net1156 vssd1 vssd1 vccd1 vccd1 final_design.reqhand.instruction\[12\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__08432__S net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06741__A _01686_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13041_ clknet_leaf_34_clk _00272_ net1243 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_10253_ net1652 _05119_ _05121_ vssd1 vssd1 vccd1 vccd1 _00016_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12551__B1 net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input46_A mem_adr_start[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10184_ final_design.uart.BAUD_counter\[1\] final_design.uart.BAUD_counter\[7\] final_design.uart.BAUD_counter\[6\]
+ final_design.uart.BAUD_counter\[0\] vssd1 vssd1 vccd1 vccd1 _05074_ sky130_fd_sc_hd__or4b_1
Xfanout1202 net1204 vssd1 vssd1 vccd1 vccd1 net1202 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_37_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1213 net1214 vssd1 vssd1 vccd1 vccd1 net1213 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_37_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1224 net1226 vssd1 vssd1 vccd1 vccd1 net1224 sky130_fd_sc_hd__clkbuf_4
Xfanout1235 net1245 vssd1 vssd1 vccd1 vccd1 net1235 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_41_1882 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_1901 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout270 net271 vssd1 vssd1 vccd1 vccd1 net270 sky130_fd_sc_hd__buf_6
Xfanout281 net284 vssd1 vssd1 vccd1 vccd1 net281 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_57_1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout292 net293 vssd1 vssd1 vccd1 vccd1 net292 sky130_fd_sc_hd__clkbuf_4
X_13943_ clknet_leaf_6_clk _01174_ net1128 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[931\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13874_ clknet_leaf_44_clk _01105_ net1208 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[862\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12825_ net1364 vssd1 vssd1 vccd1 vccd1 _00266_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_70_1522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12606__B2 final_design.data_from_mem\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09483__A0 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12756_ _06351_ _06385_ _06344_ vssd1 vssd1 vccd1 vccd1 _06393_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_35_1686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12082__A2 net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06475__X _01426_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11707_ net201 net629 vssd1 vssd1 vccd1 vccd1 _06212_ sky130_fd_sc_hd__and2_1
X_12687_ final_design.VGA_data_control.ready_data\[31\] net1021 net977 final_design.data_from_mem\[31\]
+ vssd1 vssd1 vccd1 vccd1 _06331_ sky130_fd_sc_hd__a22o_1
XANTENNA__10438__A _02991_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11638_ net432 net572 _06176_ net301 net1913 vssd1 vssd1 vccd1 vccd1 _00451_ sky130_fd_sc_hd__a32o_1
XFILLER_0_21_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11569_ net556 net420 _06140_ net302 net1969 vssd1 vssd1 vccd1 vccd1 _00418_ sky130_fd_sc_hd__a32o_1
XANTENNA__11593__A1 net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold707 final_design.cpu.reg_window\[378\] vssd1 vssd1 vccd1 vccd1 net2049 sky130_fd_sc_hd__dlygate4sd3_1
X_13308_ clknet_leaf_4_clk _00539_ net1083 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[296\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold718 final_design.cpu.reg_window\[330\] vssd1 vssd1 vccd1 vccd1 net2060 sky130_fd_sc_hd__dlygate4sd3_1
Xhold729 final_design.cpu.reg_window\[334\] vssd1 vssd1 vccd1 vccd1 net2071 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09538__A1 net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11269__A net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13239_ clknet_leaf_6_clk _00470_ net1082 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[227\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12542__B1 net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11345__B2 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07800_ net713 _02744_ net723 vssd1 vssd1 vccd1 vccd1 _02751_ sky130_fd_sc_hd__o21a_1
X_08780_ _03690_ _03730_ vssd1 vssd1 vccd1 vccd1 _03731_ sky130_fd_sc_hd__nor2_1
XFILLER_0_46_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07731_ final_design.cpu.reg_window\[218\] final_design.cpu.reg_window\[250\] net865
+ vssd1 vssd1 vccd1 vccd1 _02682_ sky130_fd_sc_hd__mux2_1
XANTENNA__11648__A2 net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07662_ final_design.cpu.reg_window\[286\] final_design.cpu.reg_window\[318\] net873
+ vssd1 vssd1 vccd1 vccd1 _02613_ sky130_fd_sc_hd__mux2_1
X_09401_ net261 _04311_ _04313_ _04319_ vssd1 vssd1 vccd1 vccd1 _04320_ sky130_fd_sc_hd__and4_1
X_06613_ _01560_ _01561_ _01562_ _01563_ net776 net783 vssd1 vssd1 vccd1 vccd1 _01564_
+ sky130_fd_sc_hd__mux4_1
X_07593_ net617 _02540_ _02541_ net527 vssd1 vssd1 vccd1 vccd1 _02544_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_75_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09332_ _04196_ _04250_ vssd1 vssd1 vccd1 vccd1 _04251_ sky130_fd_sc_hd__and2_1
XANTENNA__08277__A1 net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06544_ _01463_ _01474_ _01480_ _01482_ vssd1 vssd1 vccd1 vccd1 _01495_ sky130_fd_sc_hd__or4_4
XANTENNA__09474__A0 net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06826__A net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12073__A2 net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08744__C _01537_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09263_ net99 _04181_ vssd1 vssd1 vccd1 vccd1 _04182_ sky130_fd_sc_hd__or2_2
XANTENNA__09202__A net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06475_ final_design.data_from_mem\[18\] net969 _01425_ vssd1 vssd1 vccd1 vccd1 _01426_
+ sky130_fd_sc_hd__o21a_4
XANTENNA__12039__S net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout233_A _05983_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06545__B net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08214_ _03164_ vssd1 vssd1 vccd1 vccd1 _03165_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_1448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09194_ net594 _04111_ vssd1 vssd1 vccd1 vccd1 _04113_ sky130_fd_sc_hd__nand2_2
XFILLER_0_12_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08145_ net878 _03095_ _03084_ _03083_ vssd1 vssd1 vccd1 vccd1 _03096_ sky130_fd_sc_hd__o2bb2a_4
XANTENNA__09777__A1 _04046_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout400_A net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1142_A net1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08252__S net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08076_ net602 _03022_ _02998_ net547 vssd1 vssd1 vccd1 vccd1 _03027_ sky130_fd_sc_hd__o211a_1
XANTENNA__06686__S1 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09529__A1 net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07027_ final_design.cpu.reg_window\[78\] final_design.cpu.reg_window\[110\] net894
+ vssd1 vssd1 vccd1 vccd1 _01978_ sky130_fd_sc_hd__mux2_1
XANTENNA__07376__B net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11336__A1 final_design.data_from_mem\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12533__B1 net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout390_X net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout867_A net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout488_X net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold12 final_design.cpu.reg_window\[25\] vssd1 vssd1 vccd1 vccd1 net1354 sky130_fd_sc_hd__dlygate4sd3_1
Xhold23 final_design.cpu.reg_window\[22\] vssd1 vssd1 vccd1 vccd1 net1365 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_51_1942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold34 net120 vssd1 vssd1 vccd1 vccd1 net1376 sky130_fd_sc_hd__dlygate4sd3_1
X_08978_ net621 _03912_ net258 vssd1 vssd1 vccd1 vccd1 _03915_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_51_1953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold45 final_design.reqhand.instruction\[9\] vssd1 vssd1 vccd1 vccd1 net1387 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07392__A net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold56 final_design.uart.working_data\[1\] vssd1 vssd1 vccd1 vccd1 net1398 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12837__CLK clknet_leaf_19_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11185__Y _05895_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold67 final_design.reqhand.instruction\[18\] vssd1 vssd1 vccd1 vccd1 net1409 sky130_fd_sc_hd__dlygate4sd3_1
Xhold78 final_design.VGA_data_control.data_to_VGA\[23\] vssd1 vssd1 vccd1 vccd1 net1420
+ sky130_fd_sc_hd__dlygate4sd3_1
X_07929_ _02876_ _02877_ _02878_ _02879_ net680 net700 vssd1 vssd1 vccd1 vccd1 _02880_
+ sky130_fd_sc_hd__mux4_1
Xhold89 final_design.VGA_data_control.data_to_VGA\[24\] vssd1 vssd1 vccd1 vccd1 net1431
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout655_X net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09162__C1 _02423_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10940_ _05602_ _05622_ _05667_ vssd1 vssd1 vccd1 vccd1 _05668_ sky130_fd_sc_hd__or3_1
X_10871_ _05562_ _05578_ _05579_ vssd1 vssd1 vccd1 vccd1 _05603_ sky130_fd_sc_hd__or3_1
XFILLER_0_6_1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_1871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12610_ net1442 net999 net985 final_design.data_from_mem\[28\] vssd1 vssd1 vccd1
+ vccd1 _01303_ sky130_fd_sc_hd__a22o_1
XANTENNA_input100_A nrst vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12064__A2 net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13590_ clknet_leaf_62_clk _00821_ net1124 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[578\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_26_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_45_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11272__B1 _05843_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08363__S1 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12541_ _06204_ net345 net322 net2047 vssd1 vssd1 vccd1 vccd1 _01245_ sky130_fd_sc_hd__a22o_1
X_12472_ _06254_ net498 net330 net2078 vssd1 vssd1 vccd1 vccd1 _01178_ sky130_fd_sc_hd__a22o_1
XFILLER_0_30_1583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14211_ net1269 vssd1 vssd1 vccd1 vccd1 gpio_oeb[23] sky130_fd_sc_hd__buf_2
XANTENNA__09768__A1 net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11423_ net2024 net209 net312 vssd1 vssd1 vccd1 vccd1 _00320_ sky130_fd_sc_hd__mux2_1
XANTENNA__09768__B2 net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10378__A2 net1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11575__A1 net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_9 _06257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14142_ clknet_leaf_19_clk _01316_ net1111 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.data_to_VGA\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_65_1657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11354_ _04381_ _04384_ _05143_ vssd1 vssd1 vccd1 vccd1 _06044_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_39_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10705__B net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10305_ final_design.VGA_data_control.h_count\[3\] net1048 _05158_ vssd1 vssd1 vccd1
+ vccd1 _05159_ sky130_fd_sc_hd__or3b_1
XFILLER_0_21_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11285_ final_design.data_from_mem\[16\] _02062_ _02509_ _05912_ _05917_ vssd1 vssd1
+ vccd1 vccd1 _05983_ sky130_fd_sc_hd__a41o_1
X_14073_ clknet_leaf_13_clk _01270_ net1099 vssd1 vssd1 vccd1 vccd1 final_design.uart.working_data\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13612__CLK clknet_leaf_45_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12524__B1 net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10236_ final_design.uart.BAUD_counter\[13\] _05109_ net799 vssd1 vssd1 vccd1 vccd1
+ _05111_ sky130_fd_sc_hd__o21ai_1
X_13024_ clknet_leaf_12_clk _00255_ net1090 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11878__A2 net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1010 _05166_ vssd1 vssd1 vccd1 vccd1 net1010 sky130_fd_sc_hd__clkbuf_2
Xfanout1021 _06298_ vssd1 vssd1 vccd1 vccd1 net1021 sky130_fd_sc_hd__clkbuf_4
Xfanout1032 net1036 vssd1 vssd1 vccd1 vccd1 net1032 sky130_fd_sc_hd__buf_2
X_10167_ _05040_ _05057_ _05060_ vssd1 vssd1 vccd1 vccd1 final_design.vga.h_next_count\[7\]
+ sky130_fd_sc_hd__and3_1
Xfanout1043 final_design.VGA_adr\[10\] vssd1 vssd1 vccd1 vccd1 net1043 sky130_fd_sc_hd__buf_2
Xfanout1054 net1056 vssd1 vssd1 vccd1 vccd1 net1054 sky130_fd_sc_hd__clkbuf_2
Xfanout1065 net1069 vssd1 vssd1 vccd1 vccd1 net1065 sky130_fd_sc_hd__buf_2
Xfanout1076 net1118 vssd1 vssd1 vccd1 vccd1 net1076 sky130_fd_sc_hd__buf_2
X_10098_ net1049 _05012_ net1048 final_design.VGA_data_control.h_count\[3\] vssd1
+ vssd1 vccd1 vccd1 _05014_ sky130_fd_sc_hd__a211o_1
XANTENNA__13762__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1087 net1117 vssd1 vssd1 vccd1 vccd1 net1087 sky130_fd_sc_hd__buf_2
Xfanout1098 net1105 vssd1 vssd1 vccd1 vccd1 net1098 sky130_fd_sc_hd__clkbuf_2
XANTENNA__10440__B net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13926_ clknet_leaf_51_clk _01157_ net1174 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[914\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07929__S1 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_18_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13857_ clknet_leaf_48_clk _01088_ net1202 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[845\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_18_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06601__S1 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14118__CLK clknet_leaf_17_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12808_ net1380 vssd1 vssd1 vccd1 vccd1 _00249_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_69_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13788_ clknet_leaf_4_clk _01019_ net1079 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[776\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_31_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12739_ _05058_ _06366_ _06376_ vssd1 vssd1 vccd1 vccd1 _06379_ sky130_fd_sc_hd__and3_1
XANTENNA__11802__A2 net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_0_clk_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_2282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_2293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13142__CLK clknet_leaf_60_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10369__A2 net1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold504 final_design.cpu.reg_window\[658\] vssd1 vssd1 vccd1 vccd1 net1846 sky130_fd_sc_hd__dlygate4sd3_1
Xhold515 final_design.cpu.reg_window\[761\] vssd1 vssd1 vccd1 vccd1 net1857 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_1877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07865__S0 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold526 final_design.cpu.reg_window\[896\] vssd1 vssd1 vccd1 vccd1 net1868 sky130_fd_sc_hd__dlygate4sd3_1
Xhold537 final_design.cpu.reg_window\[81\] vssd1 vssd1 vccd1 vccd1 net1879 sky130_fd_sc_hd__dlygate4sd3_1
Xhold548 final_design.cpu.reg_window\[429\] vssd1 vssd1 vccd1 vccd1 net1890 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13292__CLK clknet_leaf_46_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09950_ _04438_ _04112_ _04436_ vssd1 vssd1 vccd1 vccd1 _04869_ sky130_fd_sc_hd__or3b_1
Xhold559 final_design.cpu.reg_window\[220\] vssd1 vssd1 vccd1 vccd1 net1901 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11318__A1 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12515__B1 net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_2075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08901_ _03665_ _03667_ vssd1 vssd1 vccd1 vccd1 _03846_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_55_2086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_2097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09881_ net470 _04797_ _04798_ net490 vssd1 vssd1 vccd1 vccd1 _04800_ sky130_fd_sc_hd__a31o_1
XANTENNA__11869__A2 net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07617__S0 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload18_A clknet_leaf_18_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11286__X _05984_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08832_ net624 _02508_ net256 _03782_ vssd1 vssd1 vccd1 vccd1 _03783_ sky130_fd_sc_hd__a211o_1
XANTENNA__12322__S net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1204 final_design.data_from_mem\[7\] vssd1 vssd1 vccd1 vccd1 net2546 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07942__B1 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11446__B net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08763_ _02391_ _02393_ final_design.CPU_instr_adr\[1\] vssd1 vssd1 vccd1 vccd1 _03714_
+ sky130_fd_sc_hd__a21boi_1
XANTENNA__08101__A net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout183_A _06067_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09144__C1 _02422_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1241 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07714_ final_design.cpu.reg_window\[923\] final_design.cpu.reg_window\[955\] net865
+ vssd1 vssd1 vccd1 vccd1 _02665_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_0_212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08694_ _02772_ _03296_ _03593_ _03644_ vssd1 vssd1 vccd1 vccd1 _03645_ sky130_fd_sc_hd__and4_2
XTAP_TAPCELL_ROW_0_223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13104__RESET_B net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07645_ final_design.cpu.reg_window\[732\] final_design.cpu.reg_window\[764\] net866
+ vssd1 vssd1 vccd1 vccd1 _02596_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout350_A _06277_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11462__A net219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout448_A net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07576_ net720 _02526_ vssd1 vssd1 vccd1 vccd1 _02527_ sky130_fd_sc_hd__nor2_1
XANTENNA__07151__S net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10057__A1 net68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06527_ _01379_ net1040 net994 net991 vssd1 vssd1 vccd1 vccd1 _01478_ sky130_fd_sc_hd__or4_1
X_09315_ _04232_ _04233_ net477 vssd1 vssd1 vccd1 vccd1 _04234_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06458_ net1057 _01393_ vssd1 vssd1 vccd1 vccd1 _01411_ sky130_fd_sc_hd__nand2_1
X_09246_ _04158_ _04164_ _04133_ vssd1 vssd1 vccd1 vccd1 _04165_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_69_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1256 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09177_ _02544_ net440 vssd1 vssd1 vccd1 vccd1 _04096_ sky130_fd_sc_hd__nand2_1
XFILLER_0_1_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout403_X net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13635__CLK clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1145_X net1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08128_ final_design.cpu.reg_window\[13\] final_design.cpu.reg_window\[45\] net850
+ vssd1 vssd1 vccd1 vccd1 _03079_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_1917 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_1376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08059_ net714 _03003_ net723 vssd1 vssd1 vccd1 vccd1 _03010_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_47_1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12506__B1 net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11070_ _05773_ _05776_ _05791_ vssd1 vssd1 vccd1 vccd1 _05793_ sky130_fd_sc_hd__or3_1
XANTENNA__11908__Y _06248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout772_X net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13785__CLK clknet_leaf_55_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10021_ _04936_ _04937_ _04938_ net726 vssd1 vssd1 vccd1 vccd1 _04940_ sky130_fd_sc_hd__a211o_2
XANTENNA__06736__A1 final_design.data_from_mem\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07326__S net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06831__S1 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13015__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11972_ _06174_ net278 net404 net1554 vssd1 vssd1 vccd1 vccd1 _00705_ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_2_clk_A clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13711_ clknet_leaf_40_clk _00942_ net1219 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[699\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_47_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10923_ _05650_ _05651_ _05631_ vssd1 vssd1 vccd1 vccd1 _05652_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_47_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_19_Right_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06595__S0 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11372__A net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13642_ clknet_leaf_50_clk _00873_ net1168 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[630\]
+ sky130_fd_sc_hd__dfrtp_1
X_10854_ net78 _05548_ _05551_ vssd1 vssd1 vccd1 vccd1 _05586_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_71_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12898__RESET_B net1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13165__CLK clknet_leaf_48_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10048__A1 _04529_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09989__A1 _04370_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11245__B1 _05946_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13573_ clknet_leaf_50_clk _00804_ net1172 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[561\]
+ sky130_fd_sc_hd__dfrtp_1
X_10785_ net669 _05509_ _05518_ net962 _05520_ vssd1 vssd1 vccd1 vccd1 _05521_ sky130_fd_sc_hd__o221a_1
XFILLER_0_66_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09453__A3 _04368_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12524_ _06186_ net355 net328 net1757 vssd1 vssd1 vccd1 vccd1 _01229_ sky130_fd_sc_hd__a22o_1
XANTENNA__08661__A1 _02545_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12455_ net1814 net193 net336 vssd1 vssd1 vccd1 vccd1 _01162_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_10_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07297__A net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11406_ net649 net177 vssd1 vssd1 vccd1 vccd1 _06090_ sky130_fd_sc_hd__and2_1
XFILLER_0_1_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12386_ net1845 net194 net269 vssd1 vssd1 vccd1 vccd1 _01097_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_28_Right_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14125_ clknet_leaf_21_clk final_design.vga.v_next_count\[5\] net1160 vssd1 vssd1
+ vccd1 vccd1 final_design.VGA_data_control.v_count\[5\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_1_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11337_ _01722_ net642 _06028_ net644 net656 vssd1 vssd1 vccd1 vccd1 _06029_ sky130_fd_sc_hd__a221o_1
XFILLER_0_65_1498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14056_ clknet_leaf_16_clk _00018_ net1091 vssd1 vssd1 vccd1 vccd1 final_design.uart.BAUD_counter\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_11268_ net660 _03932_ net732 vssd1 vssd1 vccd1 vccd1 _05968_ sky130_fd_sc_hd__o21ai_1
X_13007_ net1338 _00238_ net1234 vssd1 vssd1 vccd1 vccd1 final_design.CPU_instr_adr\[27\]
+ sky130_fd_sc_hd__dfrtp_2
X_10219_ final_design.uart.BAUD_counter\[6\] _05098_ _05100_ net799 vssd1 vssd1 vccd1
+ vccd1 _00034_ sky130_fd_sc_hd__o211a_1
XANTENNA__12142__S net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11199_ net660 _03992_ vssd1 vssd1 vccd1 vccd1 _05907_ sky130_fd_sc_hd__nor2_1
XANTENNA__11720__A1 net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_37_Right_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09677__B1 net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13508__CLK clknet_leaf_54_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09304__X _04223_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13909_ clknet_leaf_57_clk _01140_ net1144 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[897\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10597__S net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_2480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07430_ _02377_ _02378_ _02379_ _02380_ net769 net790 vssd1 vssd1 vccd1 vccd1 _02381_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__11282__A net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_2344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_2355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11713__C net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_2366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14090__CLK clknet_leaf_25_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07361_ net751 _02305_ net746 vssd1 vssd1 vccd1 vccd1 _02312_ sky130_fd_sc_hd__o21a_1
XFILLER_0_45_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1887 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09100_ _04021_ _04022_ net254 vssd1 vssd1 vccd1 vccd1 _04023_ sky130_fd_sc_hd__mux2_1
XANTENNA__11787__B2 _05959_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07292_ final_design.cpu.reg_window\[69\] final_design.cpu.reg_window\[101\] net920
+ vssd1 vssd1 vccd1 vccd1 _02243_ sky130_fd_sc_hd__mux2_1
XANTENNA__08591__A net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09031_ _03731_ _03961_ vssd1 vssd1 vccd1 vccd1 _03962_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_26_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12317__S net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_46_Right_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09601__B1 net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold301 final_design.cpu.reg_window\[733\] vssd1 vssd1 vccd1 vccd1 net1643 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_2148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold312 final_design.cpu.reg_window\[848\] vssd1 vssd1 vccd1 vccd1 net1654 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_2159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold323 final_design.cpu.reg_window\[899\] vssd1 vssd1 vccd1 vccd1 net1665 sky130_fd_sc_hd__dlygate4sd3_1
Xhold334 final_design.cpu.reg_window\[529\] vssd1 vssd1 vccd1 vccd1 net1676 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_15_Left_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold345 final_design.cpu.reg_window\[161\] vssd1 vssd1 vccd1 vccd1 net1687 sky130_fd_sc_hd__dlygate4sd3_1
Xhold356 final_design.cpu.reg_window\[178\] vssd1 vssd1 vccd1 vccd1 net1698 sky130_fd_sc_hd__dlygate4sd3_1
Xhold367 final_design.cpu.reg_window\[228\] vssd1 vssd1 vccd1 vccd1 net1709 sky130_fd_sc_hd__dlygate4sd3_1
Xhold378 final_design.cpu.reg_window\[571\] vssd1 vssd1 vccd1 vccd1 net1720 sky130_fd_sc_hd__dlygate4sd3_1
Xhold389 final_design.cpu.reg_window\[249\] vssd1 vssd1 vccd1 vccd1 net1731 sky130_fd_sc_hd__dlygate4sd3_1
X_09933_ net475 _04795_ vssd1 vssd1 vccd1 vccd1 _04852_ sky130_fd_sc_hd__or2_1
Xfanout803 _02392_ vssd1 vssd1 vccd1 vccd1 net803 sky130_fd_sc_hd__clkbuf_2
Xfanout814 net815 vssd1 vssd1 vccd1 vccd1 net814 sky130_fd_sc_hd__clkbuf_4
XANTENNA__13038__CLK clknet_leaf_45_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout825 net828 vssd1 vssd1 vccd1 vccd1 net825 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_0_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout398_A net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1885 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout836 net842 vssd1 vssd1 vccd1 vccd1 net836 sky130_fd_sc_hd__buf_2
XANTENNA__12052__S net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout847 net873 vssd1 vssd1 vccd1 vccd1 net847 sky130_fd_sc_hd__clkbuf_2
X_09864_ _04112_ _04782_ vssd1 vssd1 vccd1 vccd1 _04783_ sky130_fd_sc_hd__or2_1
Xfanout858 net860 vssd1 vssd1 vccd1 vccd1 net858 sky130_fd_sc_hd__clkbuf_4
Xhold1001 final_design.cpu.reg_window\[816\] vssd1 vssd1 vccd1 vccd1 net2343 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1105_A net1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout869 net871 vssd1 vssd1 vccd1 vccd1 net869 sky130_fd_sc_hd__clkbuf_2
Xhold1012 final_design.cpu.reg_window\[160\] vssd1 vssd1 vccd1 vccd1 net2354 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11176__B net251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08815_ final_design.CPU_instr_adr\[22\] _01756_ _03755_ _03756_ vssd1 vssd1 vccd1
+ vccd1 _03766_ sky130_fd_sc_hd__a31o_1
XANTENNA__09380__A2 net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1023 final_design.cpu.reg_window\[126\] vssd1 vssd1 vccd1 vccd1 net2365 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1034 final_design.cpu.reg_window\[312\] vssd1 vssd1 vccd1 vccd1 net2376 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06813__S1 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09795_ _04340_ _04709_ _04713_ _04348_ _04708_ vssd1 vssd1 vccd1 vccd1 _04714_ sky130_fd_sc_hd__a32o_1
XANTENNA__11891__S net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout565_A net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1045 final_design.cpu.reg_window\[508\] vssd1 vssd1 vccd1 vccd1 net2387 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_55_Right_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1056 final_design.cpu.reg_window\[736\] vssd1 vssd1 vccd1 vccd1 net2398 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_77_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1067 final_design.cpu.reg_window\[823\] vssd1 vssd1 vccd1 vccd1 net2409 sky130_fd_sc_hd__dlygate4sd3_1
X_08746_ final_design.CPU_instr_adr\[7\] net666 _01598_ vssd1 vssd1 vccd1 vccd1 _03697_
+ sky130_fd_sc_hd__and3_1
Xhold1078 final_design.cpu.reg_window\[622\] vssd1 vssd1 vccd1 vccd1 net2420 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09668__B1 _04586_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13188__CLK clknet_leaf_54_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1089 final_design.cpu.reg_window\[364\] vssd1 vssd1 vccd1 vccd1 net2431 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout353_X net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08677_ net594 _03617_ vssd1 vssd1 vccd1 vccd1 _03628_ sky130_fd_sc_hd__nand2b_2
XANTENNA_fanout732_A _01491_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12019__A2 net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07628_ final_design.cpu.reg_window\[284\] final_design.cpu.reg_window\[316\] net866
+ vssd1 vssd1 vccd1 vccd1 _02579_ sky130_fd_sc_hd__mux2_1
XANTENNA__08891__A1 net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_864 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12778__9_A clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09515__S0 net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout520_X net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_514 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07559_ _02094_ _02509_ vssd1 vssd1 vccd1 vccd1 _02510_ sky130_fd_sc_hd__or2_2
XFILLER_0_64_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout618_X net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10570_ _05314_ _05315_ vssd1 vssd1 vccd1 vccd1 _05316_ sky130_fd_sc_hd__and2_1
XFILLER_0_75_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09840__B1 net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_64_Right_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09229_ _03638_ _04146_ _03637_ vssd1 vssd1 vccd1 vccd1 _04148_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_20_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12240_ net561 _06170_ net503 net372 net1498 vssd1 vssd1 vccd1 vccd1 _00957_ sky130_fd_sc_hd__a32o_1
XFILLER_0_66_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12171_ net1540 net244 net380 vssd1 vssd1 vccd1 vccd1 _00890_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11122_ _01372_ _04993_ net1036 _05837_ wb_manage.BUSY_O vssd1 vssd1 vccd1 vccd1
+ _00212_ sky130_fd_sc_hd__o32a_1
XFILLER_0_40_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold890 final_design.cpu.reg_window\[572\] vssd1 vssd1 vccd1 vccd1 net2232 sky130_fd_sc_hd__dlygate4sd3_1
X_11053_ _05757_ _05775_ _05172_ vssd1 vssd1 vccd1 vccd1 _05777_ sky130_fd_sc_hd__a21o_1
XANTENNA__08254__S0 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06709__A1 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_73_Right_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10004_ _04918_ _04921_ vssd1 vssd1 vccd1 vccd1 _04923_ sky130_fd_sc_hd__xnor2_1
XANTENNA__11466__A0 net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11955_ _06156_ net288 net411 net2159 vssd1 vssd1 vccd1 vccd1 _00690_ sky130_fd_sc_hd__a22o_1
XFILLER_0_34_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10906_ _05634_ _05635_ vssd1 vssd1 vccd1 vccd1 _05636_ sky130_fd_sc_hd__nor2_1
XFILLER_0_80_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08882__A1 _03655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13800__CLK clknet_leaf_41_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11886_ net229 net2138 net273 vssd1 vssd1 vccd1 vccd1 _00628_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13625_ clknet_leaf_54_clk _00856_ net1177 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[613\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10837_ net78 _05548_ _05569_ vssd1 vssd1 vccd1 vccd1 _05570_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_82_Right_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_1464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13556_ clknet_leaf_10_clk _00787_ net1102 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[544\]
+ sky130_fd_sc_hd__dfrtp_1
X_10768_ _05496_ _05477_ vssd1 vssd1 vccd1 vccd1 _05504_ sky130_fd_sc_hd__and2b_1
XANTENNA__12430__A2 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1885 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09300__A net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12507_ _06169_ net342 net326 net1543 vssd1 vssd1 vccd1 vccd1 _01212_ sky130_fd_sc_hd__a22o_1
XANTENNA__13950__CLK clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10441__B2 net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12137__S net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10446__A _02863_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13487_ clknet_leaf_42_clk _00718_ net1222 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[475\]
+ sky130_fd_sc_hd__dfrtp_1
X_10699_ _05402_ _05421_ vssd1 vssd1 vccd1 vccd1 _05439_ sky130_fd_sc_hd__or2_1
X_12438_ net1645 net238 net335 vssd1 vssd1 vccd1 vccd1 _01145_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_75_2760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_2771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_2782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07296__S1 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12369_ net1761 net225 net269 vssd1 vssd1 vccd1 vccd1 _01080_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_71_2624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_2001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_2635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14108_ clknet_leaf_25_clk _01305_ net1151 vssd1 vssd1 vccd1 vccd1 final_design.reqhand.instruction\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_71_2646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14039_ clknet_leaf_15_clk _00031_ net1094 vssd1 vssd1 vccd1 vccd1 final_design.uart.BAUD_counter\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06930_ net742 _01498_ net664 net756 _01821_ vssd1 vssd1 vccd1 vccd1 _01881_ sky130_fd_sc_hd__o221ai_4
XFILLER_0_59_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13330__CLK clknet_leaf_38_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06861_ final_design.cpu.reg_window\[532\] final_design.cpu.reg_window\[564\] net947
+ vssd1 vssd1 vccd1 vccd1 _01812_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_1891 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08600_ net614 _03550_ _02423_ vssd1 vssd1 vccd1 vccd1 _03551_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_69_2553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_2564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06792_ net760 _01742_ vssd1 vssd1 vccd1 vccd1 _01743_ sky130_fd_sc_hd__nor2_1
X_09580_ _03164_ _04498_ vssd1 vssd1 vccd1 vccd1 _04499_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_69_2575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_2417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_2428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_1905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08531_ _02361_ net595 vssd1 vssd1 vccd1 vccd1 _03482_ sky130_fd_sc_hd__and2_2
XTAP_TAPCELL_ROW_65_2439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_62_clk_X clknet_leaf_62_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13480__CLK clknet_leaf_41_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08462_ _03409_ _03410_ _03411_ _03412_ net677 net691 vssd1 vssd1 vccd1 vccd1 _03413_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__08873__A1 net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07413_ _02362_ _02363_ vssd1 vssd1 vccd1 vccd1 _02364_ sky130_fd_sc_hd__or2_1
X_08393_ final_design.cpu.reg_window\[902\] final_design.cpu.reg_window\[934\] net821
+ vssd1 vssd1 vccd1 vccd1 _03344_ sky130_fd_sc_hd__mux2_1
XANTENNA__09417__A3 _01626_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07344_ final_design.data_from_mem\[11\] final_design.reqhand.instruction\[11\] net970
+ vssd1 vssd1 vccd1 vccd1 _02295_ sky130_fd_sc_hd__mux2_4
XFILLER_0_45_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12421__A2 net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08752__C _01659_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07275_ _02222_ _02223_ _02224_ _02225_ net767 net781 vssd1 vssd1 vccd1 vccd1 _02226_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__12047__S net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout313_A _06092_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1055_A net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06873__A_N net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09014_ _02448_ _03945_ vssd1 vssd1 vccd1 vccd1 _03947_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_5_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08389__B1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11886__S net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold120 final_design.VGA_data_control.ready_data\[28\] vssd1 vssd1 vccd1 vccd1 net1462
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold131 net158 vssd1 vssd1 vccd1 vccd1 net1473 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold142 final_design.cpu.reg_window\[198\] vssd1 vssd1 vccd1 vccd1 net1484 sky130_fd_sc_hd__dlygate4sd3_1
Xhold153 final_design.VGA_data_control.data_to_VGA\[25\] vssd1 vssd1 vccd1 vccd1 net1495
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09356__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10291__S0 net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold164 final_design.cpu.reg_window\[212\] vssd1 vssd1 vccd1 vccd1 net1506 sky130_fd_sc_hd__dlygate4sd3_1
Xhold175 final_design.VGA_data_control.ready_data\[24\] vssd1 vssd1 vccd1 vccd1 net1517
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout682_A net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold186 final_design.reqhand.instruction\[11\] vssd1 vssd1 vccd1 vccd1 net1528 sky130_fd_sc_hd__dlygate4sd3_1
Xhold197 net125 vssd1 vssd1 vccd1 vccd1 net1539 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout600 net601 vssd1 vssd1 vccd1 vccd1 net600 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__09338__C1 _01453_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout611 net612 vssd1 vssd1 vccd1 vccd1 net611 sky130_fd_sc_hd__clkbuf_4
X_09916_ net485 _04646_ vssd1 vssd1 vccd1 vccd1 _04835_ sky130_fd_sc_hd__nand2_1
Xfanout622 _02506_ vssd1 vssd1 vccd1 vccd1 net622 sky130_fd_sc_hd__clkbuf_4
Xfanout633 _06157_ vssd1 vssd1 vccd1 vccd1 net633 sky130_fd_sc_hd__buf_4
Xfanout644 net645 vssd1 vssd1 vccd1 vccd1 net644 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12488__A2 net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_15_clk_X clknet_leaf_15_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_6_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout655 _05142_ vssd1 vssd1 vccd1 vccd1 net655 sky130_fd_sc_hd__buf_2
XANTENNA__10499__A1 net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout666 net667 vssd1 vssd1 vccd1 vccd1 net666 sky130_fd_sc_hd__buf_2
XANTENNA__10499__B2 net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout677 net690 vssd1 vssd1 vccd1 vccd1 net677 sky130_fd_sc_hd__buf_4
XANTENNA__11696__B1 net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09847_ _04763_ _04765_ vssd1 vssd1 vccd1 vccd1 _04766_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout470_X net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout688 net689 vssd1 vssd1 vccd1 vccd1 net688 sky130_fd_sc_hd__clkbuf_4
Xfanout699 net701 vssd1 vssd1 vccd1 vccd1 net699 sky130_fd_sc_hd__buf_4
XANTENNA_fanout947_A net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11160__A2 net251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout568_X net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13823__CLK clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09778_ net729 _04681_ _04696_ vssd1 vssd1 vccd1 vccd1 _04697_ sky130_fd_sc_hd__and3_1
X_08729_ final_design.CPU_instr_adr\[15\] _01967_ vssd1 vssd1 vccd1 vccd1 _03680_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_69_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11740_ net240 net2115 net416 vssd1 vssd1 vccd1 vccd1 _00503_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13973__CLK clknet_leaf_57_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout902_X net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11671_ net671 _05848_ _06193_ vssd1 vssd1 vccd1 vccd1 _06194_ sky130_fd_sc_hd__or3_4
XANTENNA__12746__A _05058_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13410_ clknet_leaf_11_clk _00641_ net1098 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[398\]
+ sky130_fd_sc_hd__dfrtp_1
X_10622_ _05347_ _05364_ vssd1 vssd1 vccd1 vccd1 _05366_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_12_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09813__A0 net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12412__A2 net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09120__A net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11620__B1 net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13341_ clknet_leaf_5_clk _00572_ net1081 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[329\]
+ sky130_fd_sc_hd__dfrtp_1
X_10553_ net1053 _05295_ net1001 final_design.CPU_instr_adr\[5\] vssd1 vssd1 vccd1
+ vccd1 _05300_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__13203__CLK clknet_leaf_40_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06722__S0 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input76_A memory_size[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13272_ clknet_leaf_63_clk _00503_ net1121 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[260\]
+ sky130_fd_sc_hd__dfrtp_1
X_10484_ _04880_ net250 _04990_ vssd1 vssd1 vccd1 vccd1 _05234_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_27_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12176__A1 net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12223_ net581 _06151_ net514 net379 net1854 vssd1 vssd1 vccd1 vccd1 _00941_ sky130_fd_sc_hd__a32o_1
XFILLER_0_62_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12154_ net190 net2234 net387 vssd1 vssd1 vccd1 vccd1 _00875_ sky130_fd_sc_hd__mux2_1
XANTENNA__13353__CLK clknet_leaf_36_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11105_ net802 _05823_ _05825_ net963 vssd1 vssd1 vccd1 vccd1 _05826_ sky130_fd_sc_hd__o22a_1
XANTENNA__12784__15_A clknet_leaf_28_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12085_ net575 _06032_ net509 net395 net1961 vssd1 vssd1 vccd1 vccd1 _00810_ sky130_fd_sc_hd__a32o_1
XANTENNA__12479__A2 net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08227__S0 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input31_X net31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11036_ _05722_ _05739_ _05759_ vssd1 vssd1 vccd1 vccd1 _05760_ sky130_fd_sc_hd__a21o_1
XANTENNA__11384__X _06070_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1829 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11544__B net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12987_ net1318 _00218_ net1165 vssd1 vssd1 vccd1 vccd1 final_design.CPU_instr_adr\[7\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__07107__A1 net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11938_ _06139_ net278 net408 net2307 vssd1 vssd1 vccd1 vccd1 _00673_ sky130_fd_sc_hd__a22o_1
XANTENNA__07202__S1 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08855__B2 net1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11869_ _06109_ net292 net519 net2054 vssd1 vssd1 vccd1 vccd1 _00615_ sky130_fd_sc_hd__a22o_1
XFILLER_0_28_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13608_ clknet_leaf_40_clk _00839_ net1219 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[596\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12403__A2 net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13539_ clknet_leaf_0_clk _00770_ net1061 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[527\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07815__C1 _01657_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_2822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10176__A net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_2833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_2844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12094__C net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07060_ final_design.cpu.reg_window\[205\] final_design.cpu.reg_window\[237\] net930
+ vssd1 vssd1 vccd1 vccd1 _02011_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_2708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07269__S1 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11719__B net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07962_ final_design.cpu.reg_window\[17\] final_design.cpu.reg_window\[49\] net850
+ vssd1 vssd1 vccd1 vccd1 _02913_ sky130_fd_sc_hd__mux2_1
XANTENNA__13846__CLK clknet_leaf_59_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09701_ net485 _04619_ vssd1 vssd1 vccd1 vccd1 _04620_ sky130_fd_sc_hd__and2_1
X_06913_ final_design.cpu.reg_window\[18\] final_design.cpu.reg_window\[50\] net924
+ vssd1 vssd1 vccd1 vccd1 _01864_ sky130_fd_sc_hd__mux2_1
XANTENNA_wire536_X net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11678__B1 net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14211__1269 vssd1 vssd1 vccd1 vccd1 _14211__1269/HI net1269 sky130_fd_sc_hd__conb_1
XFILLER_0_4_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07893_ _02840_ _02841_ _02842_ _02843_ net683 net702 vssd1 vssd1 vccd1 vccd1 _02844_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__07346__A1 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09632_ net83 _04191_ vssd1 vssd1 vccd1 vccd1 _04551_ sky130_fd_sc_hd__xor2_2
X_06844_ _01791_ _01792_ _01793_ _01794_ net776 net794 vssd1 vssd1 vccd1 vccd1 _01795_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_74_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_1328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12870__CLK clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09563_ _04481_ vssd1 vssd1 vccd1 vccd1 _04482_ sky130_fd_sc_hd__inv_2
XANTENNA__13996__CLK clknet_leaf_46_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11454__B net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06775_ final_design.cpu.reg_window\[342\] final_design.cpu.reg_window\[374\] net920
+ vssd1 vssd1 vccd1 vccd1 _01726_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout263_A _04071_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06548__B net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08514_ final_design.cpu.reg_window\[194\] final_design.cpu.reg_window\[226\] net832
+ vssd1 vssd1 vccd1 vccd1 _03465_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09699__X _04618_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09494_ _02608_ _04087_ vssd1 vssd1 vccd1 vccd1 _04413_ sky130_fd_sc_hd__nand2_1
XFILLER_0_77_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08445_ _03392_ _03393_ _03394_ _03395_ net677 net698 vssd1 vssd1 vccd1 vccd1 _03396_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__11850__B1 net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout430_A net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13226__CLK clknet_leaf_60_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_42_clk_A clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout528_A _02356_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08376_ _03324_ _03325_ vssd1 vssd1 vccd1 vccd1 _03327_ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_22_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10405__B2 net246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07327_ final_design.cpu.reg_window\[196\] final_design.cpu.reg_window\[228\] net902
+ vssd1 vssd1 vccd1 vccd1 _02278_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_22_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08074__A2 _03022_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_36_Left_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout316_X net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1058_X net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06704__S0 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07258_ _02205_ _02206_ _02207_ _02208_ net764 net780 vssd1 vssd1 vccd1 vccd1 _02209_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_clkbuf_leaf_57_clk_A clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13376__CLK clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout897_A net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07189_ _02136_ _02137_ _02138_ _02139_ net764 net780 vssd1 vssd1 vccd1 vccd1 _02140_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_44_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08457__S0 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11629__B net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1176 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout685_X net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout430 net431 vssd1 vssd1 vccd1 vccd1 net430 sky130_fd_sc_hd__buf_4
Xfanout441 net444 vssd1 vssd1 vccd1 vccd1 net441 sky130_fd_sc_hd__clkbuf_4
Xfanout452 net455 vssd1 vssd1 vccd1 vccd1 net452 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09814__S net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout463 net464 vssd1 vssd1 vccd1 vccd1 net463 sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_45_Left_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_35_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout474 _03485_ vssd1 vssd1 vccd1 vccd1 net474 sky130_fd_sc_hd__buf_2
Xfanout485 net488 vssd1 vssd1 vccd1 vccd1 net485 sky130_fd_sc_hd__buf_2
X_12910_ clknet_leaf_61_clk _00148_ net1136 vssd1 vssd1 vccd1 vccd1 net163 sky130_fd_sc_hd__dfrtp_1
XANTENNA__11645__A net197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout496 net497 vssd1 vssd1 vccd1 vccd1 net496 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_31_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13890_ clknet_leaf_4_clk _01121_ net1083 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[878\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_31_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07334__S net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14001__CLK clknet_leaf_34_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11364__B net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12841_ clknet_leaf_19_clk _00079_ net1110 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.ready_data\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07196__S0 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11723_ net186 net629 vssd1 vssd1 vccd1 vccd1 _06220_ sky130_fd_sc_hd__and2_1
XFILLER_0_35_1879 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06943__S0 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14151__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09121__Y _04040_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11654_ net582 net423 _06184_ net300 net1563 vssd1 vssd1 vccd1 vccd1 _00459_ sky130_fd_sc_hd__a32o_1
XPHY_EDGE_ROW_54_Left_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13719__CLK clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12397__A1 net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10605_ net98 final_design.VGA_adr\[6\] vssd1 vssd1 vccd1 vccd1 _05349_ sky130_fd_sc_hd__nand2_1
XFILLER_0_52_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1833 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11585_ net432 net576 _06148_ net305 net2363 vssd1 vssd1 vccd1 vccd1 _00426_ sky130_fd_sc_hd__a32o_1
XFILLER_0_51_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13324_ clknet_leaf_46_clk _00555_ net1215 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[312\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_1877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10536_ net62 _05282_ vssd1 vssd1 vccd1 vccd1 _05284_ sky130_fd_sc_hd__or2_1
XFILLER_0_68_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13255_ clknet_leaf_62_clk _00486_ net1120 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[243\]
+ sky130_fd_sc_hd__dfrtp_1
X_10467_ net801 _05217_ _05218_ net961 vssd1 vssd1 vccd1 vccd1 _05219_ sky130_fd_sc_hd__o22a_1
XANTENNA__10724__A net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13869__CLK clknet_leaf_39_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12206_ net556 _06134_ net502 net376 net1558 vssd1 vssd1 vccd1 vccd1 _00924_ sky130_fd_sc_hd__a32o_1
XFILLER_0_62_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09565__A2 _04087_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13186_ clknet_leaf_11_clk _00417_ net1086 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[174\]
+ sky130_fd_sc_hd__dfrtp_1
X_10398_ net525 _05181_ vssd1 vssd1 vccd1 vccd1 _05182_ sky130_fd_sc_hd__or2_1
X_12137_ net243 net2072 net384 vssd1 vssd1 vccd1 vccd1 _00858_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_63_Left_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09724__S net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12893__CLK clknet_leaf_17_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12068_ net563 _05905_ net505 net392 net1943 vssd1 vssd1 vccd1 vccd1 _00793_ sky130_fd_sc_hd__a32o_1
XFILLER_0_79_1773 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11019_ _01359_ _03837_ net1059 vssd1 vssd1 vccd1 vccd1 _05744_ sky130_fd_sc_hd__mux2_1
XANTENNA__12150__S net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06649__A _01596_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07423__S1 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07244__S net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13249__CLK clknet_leaf_49_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06551__A2 net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12085__B1 net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06560_ final_design.cpu.reg_window\[349\] final_design.cpu.reg_window\[381\] net949
+ vssd1 vssd1 vccd1 vccd1 _01511_ sky130_fd_sc_hd__mux2_1
XANTENNA__11832__A0 _06017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06491_ final_design.cpu.reg_window\[990\] final_design.cpu.reg_window\[1022\] net933
+ vssd1 vssd1 vccd1 vccd1 _01442_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_16_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_72_Left_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_16_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08230_ final_design.cpu.reg_window\[843\] final_design.cpu.reg_window\[875\] net826
+ vssd1 vssd1 vccd1 vccd1 _03181_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_79_2906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13399__CLK clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_2917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08161_ final_design.cpu.reg_window\[15\] final_design.cpu.reg_window\[47\] net807
+ vssd1 vssd1 vccd1 vccd1 _03112_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09695__A net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07112_ net743 _01498_ _01851_ _02061_ _01821_ vssd1 vssd1 vccd1 vccd1 _02063_ sky130_fd_sc_hd__o221a_1
XFILLER_0_42_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08092_ final_design.cpu.reg_window\[268\] final_design.cpu.reg_window\[300\] net828
+ vssd1 vssd1 vccd1 vccd1 _03043_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload40 clknet_leaf_31_clk vssd1 vssd1 vccd1 vccd1 clkload40/Y sky130_fd_sc_hd__clkinv_4
X_07043_ net758 _01993_ vssd1 vssd1 vccd1 vccd1 _01994_ sky130_fd_sc_hd__or2_1
XFILLER_0_67_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12325__S net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11899__A0 net207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_81_Left_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11363__A2 _05143_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09961__C1 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08994_ _03925_ _03929_ final_design.CPU_instr_adr\[16\] net1016 vssd1 vssd1 vccd1
+ vccd1 _00227_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_23_1772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14024__CLK clknet_leaf_41_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07945_ net602 _02894_ _02869_ vssd1 vssd1 vccd1 vccd1 _02896_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout380_A net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12312__A1 net206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09206__Y _04125_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07876_ final_design.cpu.reg_window\[532\] final_design.cpu.reg_window\[564\] net867
+ vssd1 vssd1 vccd1 vccd1 _02827_ sky130_fd_sc_hd__mux2_1
XANTENNA__07154__S net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09615_ _03418_ _04533_ _04231_ vssd1 vssd1 vccd1 vccd1 _04534_ sky130_fd_sc_hd__o21ba_1
X_06827_ final_design.cpu.reg_window\[725\] final_design.cpu.reg_window\[757\] net938
+ vssd1 vssd1 vccd1 vccd1 _01778_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout266_X net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14174__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12076__B1 net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09546_ net490 _04368_ vssd1 vssd1 vccd1 vccd1 _04465_ sky130_fd_sc_hd__and2_1
X_06758_ _01705_ _01706_ _01707_ _01708_ net779 net795 vssd1 vssd1 vccd1 vccd1 _01709_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__11823__A0 net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09477_ net529 _02325_ net528 _02389_ net456 net465 vssd1 vssd1 vccd1 vccd1 _04396_
+ sky130_fd_sc_hd__mux4_1
X_06689_ final_design.cpu.reg_window\[217\] final_design.cpu.reg_window\[249\] net935
+ vssd1 vssd1 vccd1 vccd1 _01640_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout433_X net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12091__A3 net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08428_ final_design.cpu.reg_window\[645\] final_design.cpu.reg_window\[677\] net840
+ vssd1 vssd1 vccd1 vccd1 _03379_ sky130_fd_sc_hd__mux2_1
XANTENNA__12379__A1 net206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_24_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload1 clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 clkload1/X sky130_fd_sc_hd__clkbuf_8
X_08359_ final_design.cpu.reg_window\[839\] final_design.cpu.reg_window\[871\] net819
+ vssd1 vssd1 vccd1 vccd1 _03310_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1817 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11370_ net657 _06055_ _06057_ vssd1 vssd1 vccd1 vccd1 _06058_ sky130_fd_sc_hd__or3_1
XFILLER_0_46_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10321_ net1483 net1011 net988 final_design.data_from_mem\[6\] vssd1 vssd1 vccd1
+ vccd1 _00078_ sky130_fd_sc_hd__a22o_1
XFILLER_0_46_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06741__B _01690_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11339__C1 net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13040_ clknet_leaf_33_clk _00271_ net1238 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_10252_ final_design.uart.BAUD_counter\[19\] _05119_ net798 vssd1 vssd1 vccd1 vccd1
+ _05121_ sky130_fd_sc_hd__o21ai_1
XANTENNA__12000__B1 net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10183_ final_design.uart.BAUD_counter\[3\] final_design.uart.BAUD_counter\[2\] final_design.uart.BAUD_counter\[5\]
+ final_design.uart.BAUD_counter\[4\] vssd1 vssd1 vccd1 vccd1 _05073_ sky130_fd_sc_hd__or4b_1
XTAP_TAPCELL_ROW_37_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1203 net1204 vssd1 vssd1 vccd1 vccd1 net1203 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_37_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1214 net1227 vssd1 vssd1 vccd1 vccd1 net1214 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_37_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1225 net1226 vssd1 vssd1 vccd1 vccd1 net1225 sky130_fd_sc_hd__buf_2
Xfanout1236 net1244 vssd1 vssd1 vccd1 vccd1 net1236 sky130_fd_sc_hd__clkbuf_4
XANTENNA_input39_A mem_adr_start[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout271 _06278_ vssd1 vssd1 vccd1 vccd1 net271 sky130_fd_sc_hd__buf_6
XFILLER_0_76_1913 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_3_Left_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout282 net284 vssd1 vssd1 vccd1 vccd1 net282 sky130_fd_sc_hd__clkbuf_4
X_13942_ clknet_leaf_59_clk _01173_ net1126 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[930\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout293 _06228_ vssd1 vssd1 vccd1 vccd1 net293 sky130_fd_sc_hd__buf_2
XANTENNA__07064__S net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13873_ clknet_leaf_34_clk _01104_ net1243 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[861\]
+ sky130_fd_sc_hd__dfrtp_1
X_12824_ net1365 vssd1 vssd1 vccd1 vccd1 _00265_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__12067__B1 net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13541__CLK clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10617__A1 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1198 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11814__A0 net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12755_ _06344_ _06351_ _06385_ vssd1 vssd1 vccd1 vccd1 _06392_ sky130_fd_sc_hd__and3_1
XANTENNA__10617__B2 net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09483__A1 net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06916__S0 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11706_ net433 net574 _06211_ net297 net1684 vssd1 vssd1 vccd1 vccd1 _00484_ sky130_fd_sc_hd__a32o_1
XFILLER_0_38_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11290__A1 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12686_ _06330_ net1428 net980 vssd1 vssd1 vccd1 vccd1 _01345_ sky130_fd_sc_hd__mux2_1
XANTENNA__10438__B net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_910 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11637_ net222 net633 vssd1 vssd1 vccd1 vccd1 _06176_ sky130_fd_sc_hd__and2_1
X_14210__1268 vssd1 vssd1 vccd1 vccd1 _14210__1268/HI net1268 sky130_fd_sc_hd__conb_1
XFILLER_0_80_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13691__CLK clknet_leaf_65_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11568_ net205 net634 vssd1 vssd1 vccd1 vccd1 _06140_ sky130_fd_sc_hd__and2_1
XANTENNA__06932__A net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07341__S0 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold708 final_design.cpu.reg_window\[269\] vssd1 vssd1 vccd1 vccd1 net2050 sky130_fd_sc_hd__dlygate4sd3_1
X_13307_ clknet_leaf_65_clk _00538_ net1070 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[295\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11593__A2 net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10519_ _05249_ _05264_ _05263_ vssd1 vssd1 vccd1 vccd1 _05267_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_64_1338 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold719 final_design.cpu.reg_window\[245\] vssd1 vssd1 vccd1 vccd1 net2061 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12145__S net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10454__A _02668_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11499_ net804 _05842_ vssd1 vssd1 vccd1 vccd1 _06118_ sky130_fd_sc_hd__or2_1
XANTENNA__14047__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13238_ clknet_leaf_60_clk _00469_ net1137 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[226\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09538__A2 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11345__A2 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13169_ clknet_leaf_34_clk _00400_ net1242 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[157\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10553__B1 net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1901 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09454__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10460__Y _05214_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14081__RESET_B net1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13071__CLK clknet_leaf_42_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07730_ final_design.cpu.reg_window\[26\] final_design.cpu.reg_window\[58\] net862
+ vssd1 vssd1 vccd1 vccd1 _02681_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07661_ final_design.cpu.reg_window\[350\] final_design.cpu.reg_window\[382\] net853
+ vssd1 vssd1 vccd1 vccd1 _02612_ sky130_fd_sc_hd__mux2_1
X_09400_ net496 _04298_ _04301_ _04074_ _04318_ vssd1 vssd1 vccd1 vccd1 _04319_ sky130_fd_sc_hd__o221a_1
X_06612_ final_design.cpu.reg_window\[540\] final_design.cpu.reg_window\[572\] net947
+ vssd1 vssd1 vccd1 vccd1 _01563_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07592_ net603 _02540_ _02515_ net527 vssd1 vssd1 vccd1 vccd1 _02543_ sky130_fd_sc_hd__o211a_1
XANTENNA__07702__S net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09331_ net89 _04195_ net91 vssd1 vssd1 vccd1 vccd1 _04250_ sky130_fd_sc_hd__o21ai_1
XANTENNA__11291__Y _05989_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11805__B1 net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06543_ _01474_ _01482_ _01481_ _01464_ vssd1 vssd1 vccd1 vccd1 _01494_ sky130_fd_sc_hd__and4bb_1
XANTENNA__09474__A1 net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08277__A2 _03224_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09262_ net98 _04180_ vssd1 vssd1 vccd1 vccd1 _04181_ sky130_fd_sc_hd__and2_1
X_06474_ final_design.reqhand.instruction\[18\] net971 vssd1 vssd1 vccd1 vccd1 _01425_
+ sky130_fd_sc_hd__or2_1
XANTENNA__10348__B net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08213_ _03162_ _03163_ vssd1 vssd1 vccd1 vccd1 _03164_ sky130_fd_sc_hd__nor2_2
X_09193_ _03617_ _03649_ vssd1 vssd1 vccd1 vccd1 _04112_ sky130_fd_sc_hd__or2_2
X_12785__16 clknet_leaf_28_clk vssd1 vssd1 vccd1 vccd1 net1326 sky130_fd_sc_hd__inv_2
XFILLER_0_15_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout226_A net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08144_ _03089_ _03094_ net720 vssd1 vssd1 vccd1 vccd1 _03095_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12055__S net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08075_ net547 _03024_ vssd1 vssd1 vccd1 vccd1 _03026_ sky130_fd_sc_hd__nand2b_1
XANTENNA_fanout1135_A net1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07026_ final_design.cpu.reg_window\[142\] final_design.cpu.reg_window\[174\] net893
+ vssd1 vssd1 vccd1 vccd1 _01977_ sky130_fd_sc_hd__mux2_1
XANTENNA__11894__S net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11336__A2 net235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13414__CLK clknet_leaf_51_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1867 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold13 net107 vssd1 vssd1 vccd1 vccd1 net1355 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_1179 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold24 final_design.cpu.reg_window\[10\] vssd1 vssd1 vccd1 vccd1 net1366 sky130_fd_sc_hd__dlygate4sd3_1
X_08977_ _02456_ _03913_ vssd1 vssd1 vccd1 vccd1 _03914_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_23_1580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout383_X net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout762_A net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold35 final_design.cpu.reg_window\[29\] vssd1 vssd1 vccd1 vccd1 net1377 sky130_fd_sc_hd__dlygate4sd3_1
Xhold46 final_design.VGA_data_control.data_to_VGA\[26\] vssd1 vssd1 vccd1 vccd1 net1388
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_51_1954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07928_ final_design.cpu.reg_window\[150\] final_design.cpu.reg_window\[182\] net837
+ vssd1 vssd1 vccd1 vccd1 _02879_ sky130_fd_sc_hd__mux2_1
Xhold57 final_design.reqhand.instruction\[22\] vssd1 vssd1 vccd1 vccd1 net1399 sky130_fd_sc_hd__dlygate4sd3_1
Xhold68 net129 vssd1 vssd1 vccd1 vccd1 net1410 sky130_fd_sc_hd__dlygate4sd3_1
Xhold79 final_design.VGA_data_control.data_to_VGA\[14\] vssd1 vssd1 vccd1 vccd1 net1421
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09162__B1 _01658_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13564__CLK clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07859_ _02806_ _02807_ _02808_ _02809_ net687 net705 vssd1 vssd1 vccd1 vccd1 _02810_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout550_X net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout648_X net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10870_ _05600_ _05601_ vssd1 vssd1 vccd1 vccd1 _05602_ sky130_fd_sc_hd__or2_1
XFILLER_0_78_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_1872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09529_ net494 _04439_ _04447_ _04231_ vssd1 vssd1 vccd1 vccd1 _04448_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_49_1883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11272__A1 _04509_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12540_ _06203_ net342 net322 net2150 vssd1 vssd1 vccd1 vccd1 _01244_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_45_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_1297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12471_ _06131_ net346 net331 net1945 vssd1 vssd1 vccd1 vccd1 _01177_ sky130_fd_sc_hd__a22o_1
X_14210_ net1268 vssd1 vssd1 vccd1 vccd1 gpio_oeb[22] sky130_fd_sc_hd__buf_2
XFILLER_0_69_1761 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11422_ net1912 net212 net310 vssd1 vssd1 vccd1 vccd1 _00319_ sky130_fd_sc_hd__mux2_1
XANTENNA__12221__B1 net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08443__S net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06752__A net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11575__A2 net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14141_ clknet_leaf_19_clk _01315_ net1157 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.data_to_VGA\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_62_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11353_ _01660_ net641 _06042_ net643 net656 vssd1 vssd1 vccd1 vccd1 _06043_ sky130_fd_sc_hd__a221o_1
XFILLER_0_21_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_39_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10304_ final_design.VGA_data_control.data_to_VGA\[31\] final_design.VGA_data_control.data_to_VGA\[30\]
+ final_design.VGA_data_control.data_to_VGA\[29\] final_design.VGA_data_control.data_to_VGA\[28\]
+ final_design.VGA_data_control.h_count\[1\] final_design.VGA_data_control.h_count\[2\]
+ vssd1 vssd1 vccd1 vccd1 _05158_ sky130_fd_sc_hd__mux4_1
X_14072_ clknet_leaf_14_clk _01269_ net1106 vssd1 vssd1 vccd1 vccd1 final_design.uart.working_data\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_11284_ _03613_ _05913_ vssd1 vssd1 vccd1 vccd1 _05982_ sky130_fd_sc_hd__nor2_1
XANTENNA__13094__CLK clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13023_ clknet_leaf_8_clk _00254_ net1154 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_10235_ _05109_ _05110_ vssd1 vssd1 vccd1 vccd1 _00009_ sky130_fd_sc_hd__nor2_1
Xfanout1000 net1001 vssd1 vssd1 vccd1 vccd1 net1000 sky130_fd_sc_hd__clkbuf_4
Xfanout1011 _05166_ vssd1 vssd1 vccd1 vccd1 net1011 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09127__X _04046_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1022 _06298_ vssd1 vssd1 vccd1 vccd1 net1022 sky130_fd_sc_hd__clkbuf_2
X_10166_ _05054_ _05058_ vssd1 vssd1 vccd1 vccd1 _05060_ sky130_fd_sc_hd__nand2_1
Xfanout1033 net1035 vssd1 vssd1 vccd1 vccd1 net1033 sky130_fd_sc_hd__buf_2
XANTENNA__13907__CLK clknet_leaf_36_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1044 final_design.VGA_adr\[10\] vssd1 vssd1 vccd1 vccd1 net1044 sky130_fd_sc_hd__clkbuf_2
Xfanout1055 net1056 vssd1 vssd1 vccd1 vccd1 net1055 sky130_fd_sc_hd__clkbuf_4
Xfanout1066 net1068 vssd1 vssd1 vccd1 vccd1 net1066 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_76_1721 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12288__B1 net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1077 net1080 vssd1 vssd1 vccd1 vccd1 net1077 sky130_fd_sc_hd__clkbuf_4
X_10097_ final_design.VGA_data_control.h_count\[1\] final_design.VGA_data_control.h_count\[2\]
+ vssd1 vssd1 vccd1 vccd1 _05013_ sky130_fd_sc_hd__and2_1
XANTENNA__11536__C _02095_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1088 net1090 vssd1 vssd1 vccd1 vccd1 net1088 sky130_fd_sc_hd__clkbuf_4
Xfanout1099 net1105 vssd1 vssd1 vccd1 vccd1 net1099 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_76_1765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13925_ clknet_leaf_50_clk _01156_ net1173 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[913\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_18_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkload4_A clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13856_ clknet_leaf_10_clk _01087_ net1101 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[844\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06486__X _01437_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12807_ net1359 vssd1 vssd1 vccd1 vccd1 _00248_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__09303__A net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13787_ clknet_leaf_65_clk _01018_ net1072 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[775\]
+ sky130_fd_sc_hd__dfrtp_1
X_10999_ _04042_ _05715_ _05724_ _04040_ vssd1 vssd1 vccd1 vccd1 _05725_ sky130_fd_sc_hd__a22o_1
XFILLER_0_70_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11263__A1 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12738_ net954 _06377_ _06378_ net796 final_design.VGA_adr\[2\] vssd1 vssd1 vccd1
+ vccd1 _01349_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_61_2283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_61_2294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12669_ final_design.VGA_data_control.ready_data\[22\] net1019 net974 final_design.data_from_mem\[22\]
+ vssd1 vssd1 vccd1 vccd1 _06322_ sky130_fd_sc_hd__a22o_1
XANTENNA__12212__B1 net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13437__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold505 final_design.cpu.reg_window\[148\] vssd1 vssd1 vccd1 vccd1 net1847 sky130_fd_sc_hd__dlygate4sd3_1
Xhold516 final_design.cpu.reg_window\[1004\] vssd1 vssd1 vccd1 vccd1 net1858 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07865__S1 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold527 final_design.cpu.reg_window\[832\] vssd1 vssd1 vccd1 vccd1 net1869 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_1889 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold538 final_design.cpu.reg_window\[777\] vssd1 vssd1 vccd1 vccd1 net1880 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold549 final_design.cpu.reg_window\[512\] vssd1 vssd1 vccd1 vccd1 net1891 sky130_fd_sc_hd__dlygate4sd3_1
X_08900_ final_design.CPU_instr_adr\[26\] net1015 _03842_ _03845_ vssd1 vssd1 vccd1
+ vccd1 _00237_ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_55_2076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_2087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09880_ net475 _04795_ vssd1 vssd1 vccd1 vccd1 _04799_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_55_2098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07617__S1 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08831_ net624 _03781_ vssd1 vssd1 vccd1 vccd1 _03782_ sky130_fd_sc_hd__nor2_1
XANTENNA__13587__CLK clknet_leaf_40_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11727__B net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10190__Y _05080_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1205 final_design.reqhand.data_from_UART\[5\] vssd1 vssd1 vccd1 vccd1 net2547
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07942__A1 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12900__Q net166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12279__B1 net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08762_ net1018 _02361_ vssd1 vssd1 vccd1 vccd1 _03713_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_40_1190 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09144__B1 _02325_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07713_ final_design.cpu.reg_window\[987\] final_design.cpu.reg_window\[1019\] net865
+ vssd1 vssd1 vccd1 vccd1 _02664_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_1805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08693_ _03359_ _03425_ _03636_ _03643_ vssd1 vssd1 vccd1 vccd1 _03644_ sky130_fd_sc_hd__and4_1
XFILLER_0_75_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_0_213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12294__A3 net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07644_ net712 _02594_ vssd1 vssd1 vccd1 vccd1 _02595_ sky130_fd_sc_hd__nor2_1
XFILLER_0_79_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11462__B net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07575_ _02522_ _02523_ _02524_ _02525_ net685 net703 vssd1 vssd1 vccd1 vccd1 _02526_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout343_A net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1085_A net1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09314_ net537 net535 net534 net533 net457 net466 vssd1 vssd1 vccd1 vccd1 _04233_
+ sky130_fd_sc_hd__mux4_2
XANTENNA__10057__A2 _04940_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06526_ _01465_ _01468_ _01475_ vssd1 vssd1 vccd1 vccd1 _01477_ sky130_fd_sc_hd__or3_4
XFILLER_0_75_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11889__S net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09245_ _04132_ _04162_ vssd1 vssd1 vccd1 vccd1 _04164_ sky130_fd_sc_hd__nor2_1
X_06457_ wb_manage.BUSY_O net1057 net34 vssd1 vssd1 vccd1 vccd1 _01410_ sky130_fd_sc_hd__and3b_2
XANTENNA_fanout510_A net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12574__A net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_1901 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1268 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12203__B1 net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09176_ _03631_ _03650_ vssd1 vssd1 vccd1 vccd1 _04095_ sky130_fd_sc_hd__or2_2
XANTENNA__08263__S net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11557__A2 net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08127_ final_design.cpu.reg_window\[77\] final_design.cpu.reg_window\[109\] net850
+ vssd1 vssd1 vccd1 vccd1 _03078_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09883__A _04341_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08058_ net721 _03008_ vssd1 vssd1 vccd1 vccd1 _03009_ sky130_fd_sc_hd__nor2_1
XFILLER_0_31_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout977_A _06299_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11309__A2 net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07009_ final_design.cpu.reg_window\[719\] final_design.cpu.reg_window\[751\] net887
+ vssd1 vssd1 vccd1 vccd1 _01960_ sky130_fd_sc_hd__mux2_1
XANTENNA__09907__C1 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10822__A net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09383__A0 _01657_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10020_ _04936_ _04937_ _04938_ vssd1 vssd1 vccd1 vccd1 _04939_ sky130_fd_sc_hd__a21oi_2
XANTENNA__11637__B net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout765_X net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12954__CLK clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08011__B net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11971_ _06173_ net286 net406 net1717 vssd1 vssd1 vccd1 vccd1 _00704_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout932_X net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12285__A3 net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13710_ clknet_leaf_43_clk _00941_ net1218 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[698\]
+ sky130_fd_sc_hd__dfrtp_1
X_10922_ net83 net1046 vssd1 vssd1 vccd1 vccd1 _05651_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_47_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07342__S net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06595__S1 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13641_ clknet_leaf_37_clk _00872_ net1228 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[629\]
+ sky130_fd_sc_hd__dfrtp_1
X_10853_ final_design.CPU_instr_adr\[20\] _03893_ net1060 vssd1 vssd1 vccd1 vccd1
+ _05585_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10048__A2 _04530_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13572_ clknet_leaf_54_clk _00803_ net1177 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[560\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09989__A2 _04773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10784_ net962 _05519_ vssd1 vssd1 vccd1 vccd1 _05520_ sky130_fd_sc_hd__nand2_1
X_12523_ _06185_ net353 net328 net1681 vssd1 vssd1 vccd1 vccd1 _01228_ sky130_fd_sc_hd__a22o_1
XFILLER_0_13_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08661__A2 _03610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12454_ net2003 net194 net335 vssd1 vssd1 vccd1 vccd1 _01161_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08949__B1 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11405_ net589 _06087_ _06088_ vssd1 vssd1 vccd1 vccd1 _06089_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_10_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12385_ net2197 _06017_ net270 vssd1 vssd1 vccd1 vccd1 _01096_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14124_ clknet_leaf_21_clk final_design.vga.v_next_count\[4\] net1160 vssd1 vssd1
+ vccd1 vccd1 final_design.VGA_data_control.v_count\[4\] sky130_fd_sc_hd__dfrtp_1
X_11336_ final_design.data_from_mem\[23\] net235 net233 vssd1 vssd1 vccd1 vccd1 _06028_
+ sky130_fd_sc_hd__a21o_2
XFILLER_0_61_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14055_ clknet_leaf_16_clk _00016_ net1091 vssd1 vssd1 vccd1 vccd1 final_design.uart.BAUD_counter\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_11267_ final_design.data_from_mem\[15\] _05914_ _05917_ vssd1 vssd1 vccd1 vccd1
+ _05967_ sky130_fd_sc_hd__a21o_1
X_13006_ net1337 _00237_ net1234 vssd1 vssd1 vccd1 vccd1 final_design.CPU_instr_adr\[26\]
+ sky130_fd_sc_hd__dfrtp_2
X_10218_ _05099_ vssd1 vssd1 vccd1 vccd1 _05100_ sky130_fd_sc_hd__inv_2
XFILLER_0_20_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08202__A net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11198_ final_design.data_from_mem\[7\] final_design.reqhand.data_from_UART\[7\]
+ net251 vssd1 vssd1 vccd1 vccd1 _05906_ sky130_fd_sc_hd__mux2_1
XANTENNA__11181__B1 net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11720__A2 net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10149_ final_design.VGA_data_control.h_count\[0\] _05013_ vssd1 vssd1 vccd1 vccd1
+ _05048_ sky130_fd_sc_hd__nand2_1
XFILLER_0_27_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12276__A3 net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1901 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13908_ clknet_leaf_8_clk _01139_ net1151 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[896\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_67_2481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07252__S net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11282__B net223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_2345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13839_ clknet_leaf_42_clk _01070_ net1223 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[827\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_63_2356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_2367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07360_ net759 _02310_ vssd1 vssd1 vccd1 vccd1 _02311_ sky130_fd_sc_hd__or2_1
XFILLER_0_35_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11787__A2 net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07291_ net532 _02240_ vssd1 vssd1 vccd1 vccd1 _02242_ sky130_fd_sc_hd__xor2_1
XANTENNA__11502__S net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09030_ _03688_ _03689_ vssd1 vssd1 vccd1 vccd1 _03961_ sky130_fd_sc_hd__nor2_1
XFILLER_0_2_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10626__B final_design.VGA_adr\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_57_2138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold302 final_design.cpu.reg_window\[171\] vssd1 vssd1 vccd1 vccd1 net1644 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08404__A2 _03352_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_2149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12200__A3 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold313 final_design.cpu.reg_window\[759\] vssd1 vssd1 vccd1 vccd1 net1655 sky130_fd_sc_hd__dlygate4sd3_1
Xhold324 final_design.cpu.reg_window\[225\] vssd1 vssd1 vccd1 vccd1 net1666 sky130_fd_sc_hd__dlygate4sd3_1
Xhold335 final_design.cpu.reg_window\[787\] vssd1 vssd1 vccd1 vccd1 net1677 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold346 final_design.cpu.reg_window\[470\] vssd1 vssd1 vccd1 vccd1 net1688 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkload30_A clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold357 final_design.cpu.reg_window\[48\] vssd1 vssd1 vccd1 vccd1 net1699 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11297__X _05994_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09932_ _04179_ _04850_ vssd1 vssd1 vccd1 vccd1 _04851_ sky130_fd_sc_hd__or2_1
Xhold368 final_design.cpu.reg_window\[665\] vssd1 vssd1 vccd1 vccd1 net1710 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12977__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold379 final_design.cpu.reg_window\[917\] vssd1 vssd1 vccd1 vccd1 net1721 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout804 _02295_ vssd1 vssd1 vccd1 vccd1 net804 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09365__B1 net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout815 net818 vssd1 vssd1 vccd1 vccd1 net815 sky130_fd_sc_hd__buf_2
Xfanout826 net828 vssd1 vssd1 vccd1 vccd1 net826 sky130_fd_sc_hd__clkbuf_4
Xfanout837 net841 vssd1 vssd1 vccd1 vccd1 net837 sky130_fd_sc_hd__clkbuf_4
X_09863_ _04690_ _04779_ net482 vssd1 vssd1 vccd1 vccd1 _04782_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout848 net852 vssd1 vssd1 vccd1 vccd1 net848 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout293_A _06228_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout859 net860 vssd1 vssd1 vccd1 vccd1 net859 sky130_fd_sc_hd__clkbuf_4
X_08814_ _03764_ vssd1 vssd1 vccd1 vccd1 _03765_ sky130_fd_sc_hd__inv_2
Xhold1002 final_design.cpu.reg_window\[112\] vssd1 vssd1 vccd1 vccd1 net2344 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1013 final_design.cpu.reg_window\[119\] vssd1 vssd1 vccd1 vccd1 net2355 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1000_A net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1024 final_design.cpu.reg_window\[510\] vssd1 vssd1 vccd1 vccd1 net2366 sky130_fd_sc_hd__dlygate4sd3_1
X_09794_ net484 _04712_ vssd1 vssd1 vccd1 vccd1 _04713_ sky130_fd_sc_hd__nand2_1
XANTENNA__09380__A3 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1035 final_design.reqhand.instruction\[2\] vssd1 vssd1 vccd1 vccd1 net2377 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1046 final_design.reqhand.instruction\[5\] vssd1 vssd1 vccd1 vccd1 net2388 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_1572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08745_ final_design.CPU_instr_adr\[8\] _02186_ vssd1 vssd1 vccd1 vccd1 _03696_ sky130_fd_sc_hd__and2_1
Xhold1057 final_design.cpu.reg_window\[292\] vssd1 vssd1 vccd1 vccd1 net2399 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout460_A net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1068 final_design.cpu.reg_window\[1013\] vssd1 vssd1 vccd1 vccd1 net2410 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1079 final_design.VGA_data_control.data_to_VGA\[5\] vssd1 vssd1 vccd1 vccd1 net2421
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12267__A3 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout558_A net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09668__B2 _04342_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13325__RESET_B net1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08676_ _03625_ _03626_ _03619_ _03621_ vssd1 vssd1 vccd1 vccd1 _03627_ sky130_fd_sc_hd__o211a_2
XFILLER_0_75_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_1411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_1668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07627_ final_design.cpu.reg_window\[348\] final_design.cpu.reg_window\[380\] net866
+ vssd1 vssd1 vccd1 vccd1 _02578_ sky130_fd_sc_hd__mux2_1
XANTENNA__11192__B net251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout725_A net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout346_X net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13602__CLK clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12424__B1 net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09515__S1 net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07558_ _01998_ _02028_ vssd1 vssd1 vccd1 vccd1 _02509_ sky130_fd_sc_hd__nor2_1
XFILLER_0_75_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11778__A2 net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06509_ net1041 net993 net990 _01376_ vssd1 vssd1 vccd1 vccd1 _01460_ sky130_fd_sc_hd__a31o_1
XANTENNA_clkbuf_3_2_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout513_X net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07489_ _02185_ _02186_ vssd1 vssd1 vccd1 vccd1 _02440_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_36_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11412__S net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09228_ _03638_ _04146_ vssd1 vssd1 vccd1 vccd1 _04147_ sky130_fd_sc_hd__nand2_1
XFILLER_0_49_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13752__CLK clknet_leaf_65_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09159_ net614 _03550_ _01597_ _02423_ vssd1 vssd1 vccd1 vccd1 _04078_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_20_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_1737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12170_ net1560 net237 net381 vssd1 vssd1 vccd1 vccd1 _00889_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout882_X net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11121_ _01373_ net1029 _04993_ vssd1 vssd1 vccd1 vccd1 _05837_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_13_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11950__A2 net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14108__CLK clknet_leaf_25_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10552__A net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold880 final_design.cpu.reg_window\[1003\] vssd1 vssd1 vccd1 vccd1 net2222 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09356__A0 _04058_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold891 final_design.cpu.reg_window\[950\] vssd1 vssd1 vccd1 vccd1 net2233 sky130_fd_sc_hd__dlygate4sd3_1
X_11052_ _05757_ _05775_ vssd1 vssd1 vccd1 vccd1 _05776_ sky130_fd_sc_hd__nor2_1
XANTENNA__09118__A net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08254__S1 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06709__A2 _01659_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10003_ _04919_ _04921_ vssd1 vssd1 vccd1 vccd1 _04922_ sky130_fd_sc_hd__nand2_1
XANTENNA__11702__A2 net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input21_A DAT_I[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13132__CLK clknet_leaf_46_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12258__A3 net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11954_ _06155_ net286 net410 net1944 vssd1 vssd1 vccd1 vccd1 _00689_ sky130_fd_sc_hd__a22o_1
XFILLER_0_38_1855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07072__S net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10905_ _05629_ _05633_ vssd1 vssd1 vccd1 vccd1 _05635_ sky130_fd_sc_hd__and2b_1
X_11885_ net230 net2028 net272 vssd1 vssd1 vccd1 vccd1 _00627_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13282__CLK clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13624_ clknet_leaf_65_clk _00855_ net1072 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[612\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11218__A1 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10836_ _05567_ _05568_ _05548_ vssd1 vssd1 vccd1 vccd1 _05569_ sky130_fd_sc_hd__o21ba_1
XANTENNA__12415__B1 net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13555_ clknet_leaf_38_clk _00786_ net1206 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[543\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10767_ _05479_ _05498_ _05478_ vssd1 vssd1 vccd1 vccd1 _05503_ sky130_fd_sc_hd__and3b_1
XANTENNA__10286__X _05142_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12430__A3 net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11322__S net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06645__A1 net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12506_ _06168_ net343 net326 net1656 vssd1 vssd1 vccd1 vccd1 _01211_ sky130_fd_sc_hd__a22o_1
XANTENNA__10441__A2 net1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13486_ clknet_leaf_43_clk _00717_ net1222 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[474\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10698_ _05436_ _05437_ vssd1 vssd1 vccd1 vccd1 _05438_ sky130_fd_sc_hd__nor2_1
XFILLER_0_81_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10446__B net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12437_ net2128 net225 net335 vssd1 vssd1 vccd1 vccd1 _01144_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_1796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_2750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09727__S net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09595__B1 net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_2761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12368_ net1562 net239 net268 vssd1 vssd1 vccd1 vccd1 _01079_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_2772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_2783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_2614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_2625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14107_ clknet_leaf_24_clk _01304_ net1163 vssd1 vssd1 vccd1 vccd1 final_design.reqhand.instruction\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_71_2636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11319_ net737 _03886_ _06012_ vssd1 vssd1 vccd1 vccd1 _06013_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11941__A2 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_71_2647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12153__S net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10462__A _02540_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12299_ net1762 net241 net365 vssd1 vssd1 vccd1 vccd1 _01013_ sky130_fd_sc_hd__mux2_1
X_14038_ clknet_leaf_15_clk _00028_ net1094 vssd1 vssd1 vccd1 vccd1 final_design.uart.BAUD_counter\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06860_ final_design.cpu.reg_window\[596\] final_design.cpu.reg_window\[628\] net947
+ vssd1 vssd1 vccd1 vccd1 _01811_ sky130_fd_sc_hd__mux2_1
XANTENNA__09315__X _04234_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_2554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06791_ _01738_ _01739_ _01740_ _01741_ net771 net790 vssd1 vssd1 vccd1 vccd1 _01742_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_69_2565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12249__A3 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_2576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_2418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08530_ _03468_ _03469_ _03480_ net876 vssd1 vssd1 vccd1 vccd1 _03481_ sky130_fd_sc_hd__a22oi_4
XTAP_TAPCELL_ROW_65_2429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13625__CLK clknet_leaf_54_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_1917 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08461_ final_design.cpu.reg_window\[516\] final_design.cpu.reg_window\[548\] net819
+ vssd1 vssd1 vccd1 vccd1 _03412_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07412_ net528 _02361_ vssd1 vssd1 vccd1 vccd1 _02363_ sky130_fd_sc_hd__and2_1
XFILLER_0_9_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12406__B1 net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08392_ final_design.cpu.reg_window\[966\] final_design.cpu.reg_window\[998\] net823
+ vssd1 vssd1 vccd1 vccd1 _03343_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13775__CLK clknet_leaf_43_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07343_ _02281_ _02282_ _02293_ net881 vssd1 vssd1 vccd1 vccd1 _02294_ sky130_fd_sc_hd__a22oi_4
XANTENNA__12328__S net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_14_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07274_ final_design.cpu.reg_window\[6\] final_design.cpu.reg_window\[38\] net901
+ vssd1 vssd1 vccd1 vccd1 _02225_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09013_ net623 _03944_ vssd1 vssd1 vccd1 vccd1 _03946_ sky130_fd_sc_hd__nor2_1
XFILLER_0_72_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08389__A1 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout306_A net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12185__A2 net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold110 net121 vssd1 vssd1 vccd1 vccd1 net1452 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold121 final_design.VGA_data_control.ready_data\[1\] vssd1 vssd1 vccd1 vccd1 net1463
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold132 net117 vssd1 vssd1 vccd1 vccd1 net1474 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_1_clk_A clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11393__B1 net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold143 final_design.cpu.reg_window\[719\] vssd1 vssd1 vccd1 vccd1 net1485 sky130_fd_sc_hd__dlygate4sd3_1
Xhold154 final_design.VGA_data_control.ready_data\[27\] vssd1 vssd1 vccd1 vccd1 net1496
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11932__A2 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold165 final_design.VGA_data_control.ready_data\[21\] vssd1 vssd1 vccd1 vccd1 net1507
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold176 net133 vssd1 vssd1 vccd1 vccd1 net1518 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10291__S1 net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09338__B1 _03523_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout601 _02514_ vssd1 vssd1 vccd1 vccd1 net601 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07157__S net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold187 final_design.VGA_data_control.ready_data\[19\] vssd1 vssd1 vccd1 vccd1 net1529
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold198 final_design.cpu.reg_window\[647\] vssd1 vssd1 vccd1 vccd1 net1540 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13155__CLK clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout612 _02513_ vssd1 vssd1 vccd1 vccd1 net612 sky130_fd_sc_hd__buf_4
X_09915_ net533 net532 net531 net529 net452 net460 vssd1 vssd1 vccd1 vccd1 _04834_
+ sky130_fd_sc_hd__mux4_1
Xfanout623 _02506_ vssd1 vssd1 vccd1 vccd1 net623 sky130_fd_sc_hd__clkbuf_2
Xfanout634 net635 vssd1 vssd1 vccd1 vccd1 net634 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout296_X net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout675_A net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout645 _05853_ vssd1 vssd1 vccd1 vccd1 net645 sky130_fd_sc_hd__buf_2
XFILLER_0_42_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout656 _05142_ vssd1 vssd1 vccd1 vccd1 net656 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11696__A1 net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout667 _01498_ vssd1 vssd1 vccd1 vccd1 net667 sky130_fd_sc_hd__buf_4
X_09846_ _04673_ _04764_ net449 vssd1 vssd1 vccd1 vccd1 _04765_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09353__A3 _04086_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout678 net690 vssd1 vssd1 vccd1 vccd1 net678 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout1003_X net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout689 net690 vssd1 vssd1 vccd1 vccd1 net689 sky130_fd_sc_hd__clkbuf_4
X_09777_ _04046_ _04350_ _04682_ _04695_ vssd1 vssd1 vccd1 vccd1 _04696_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout463_X net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout842_A _01818_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06989_ net544 _01939_ vssd1 vssd1 vccd1 vccd1 _01940_ sky130_fd_sc_hd__nor2_1
X_08728_ _01363_ _01968_ vssd1 vssd1 vccd1 vccd1 _03679_ sky130_fd_sc_hd__nor2_1
XFILLER_0_16_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09510__B1 net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11999__A2 net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout630_X net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08659_ net260 _03596_ _03609_ _03595_ vssd1 vssd1 vccd1 vccd1 _03610_ sky130_fd_sc_hd__o211a_2
XFILLER_0_51_1318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout728_X net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11670_ net805 _02358_ net803 vssd1 vssd1 vccd1 vccd1 _06193_ sky130_fd_sc_hd__nand3_1
X_10621_ _05347_ _05364_ vssd1 vssd1 vccd1 vccd1 _05365_ sky130_fd_sc_hd__nand2_1
XANTENNA__09401__A net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09813__A1 net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10959__B1 net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_12_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13340_ clknet_leaf_5_clk _00571_ net1081 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[328\]
+ sky130_fd_sc_hd__dfrtp_1
X_10552_ net964 _05298_ vssd1 vssd1 vccd1 vccd1 _05299_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06722__S1 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13271_ clknet_leaf_6_clk _00502_ net1134 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[259\]
+ sky130_fd_sc_hd__dfrtp_1
X_10483_ net36 _05220_ _05228_ _05229_ vssd1 vssd1 vccd1 vccd1 _05233_ sky130_fd_sc_hd__a31oi_2
X_12222_ net578 _06150_ net510 net378 net1841 vssd1 vssd1 vccd1 vccd1 _00940_ sky130_fd_sc_hd__a32o_1
XANTENNA_input69_A memory_size[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11923__A2 net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12153_ net192 net2359 net387 vssd1 vssd1 vccd1 vccd1 _00874_ sky130_fd_sc_hd__mux2_1
XFILLER_0_40_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11104_ net959 _05822_ _05824_ net957 vssd1 vssd1 vccd1 vccd1 _05825_ sky130_fd_sc_hd__o22a_1
XANTENNA__07067__S net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14080__CLK clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12084_ net2328 net393 net500 _06025_ vssd1 vssd1 vccd1 vccd1 _00809_ sky130_fd_sc_hd__a22o_1
XANTENNA__08227__S1 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11035_ _05720_ _05739_ _05738_ vssd1 vssd1 vccd1 vccd1 _05759_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_21_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13648__CLK clknet_leaf_36_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input24_X net24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10895__C1 net1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12986_ net1317 _00217_ net1165 vssd1 vssd1 vccd1 vccd1 final_design.CPU_instr_adr\[6\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__13798__CLK clknet_leaf_51_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11937_ _06138_ net290 net410 net1890 vssd1 vssd1 vccd1 vccd1 _00672_ sky130_fd_sc_hd__a22o_1
XFILLER_0_73_1598 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11868_ net428 net199 net553 net518 net1784 vssd1 vssd1 vccd1 vccd1 _00614_ sky130_fd_sc_hd__a32o_1
XFILLER_0_28_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10819_ _05551_ _05552_ vssd1 vssd1 vccd1 vccd1 _05553_ sky130_fd_sc_hd__nand2_1
X_13607_ clknet_leaf_62_clk _00838_ net1119 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[595\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11560__B net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12148__S net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13028__CLK clknet_leaf_54_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11799_ net648 _05869_ _06024_ vssd1 vssd1 vccd1 vccd1 _06236_ sky130_fd_sc_hd__and3_1
XANTENNA__09804__A1 net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13538_ clknet_leaf_3_clk _00769_ net1067 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[526\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_2823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_58_2200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_2834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07910__S0 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_77_2845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13469_ clknet_leaf_2_clk _00700_ net1077 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[457\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_2709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13178__CLK clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11288__A net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07961_ final_design.cpu.reg_window\[81\] final_design.cpu.reg_window\[113\] net848
+ vssd1 vssd1 vccd1 vccd1 _02912_ sky130_fd_sc_hd__mux2_1
XANTENNA__11127__B1 net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09700_ _04457_ _04618_ net474 vssd1 vssd1 vccd1 vccd1 _04619_ sky130_fd_sc_hd__mux2_1
X_06912_ final_design.cpu.reg_window\[82\] final_design.cpu.reg_window\[114\] net924
+ vssd1 vssd1 vccd1 vccd1 _01863_ sky130_fd_sc_hd__mux2_1
XANTENNA__11678__A1 net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07892_ final_design.cpu.reg_window\[407\] final_design.cpu.reg_window\[439\] net852
+ vssd1 vssd1 vccd1 vccd1 _02843_ sky130_fd_sc_hd__mux2_1
XANTENNA__08597__A net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09631_ net730 _04546_ _04549_ vssd1 vssd1 vccd1 vccd1 _04550_ sky130_fd_sc_hd__and3_1
X_06843_ final_design.cpu.reg_window\[404\] final_design.cpu.reg_window\[436\] net948
+ vssd1 vssd1 vccd1 vccd1 _01794_ sky130_fd_sc_hd__mux2_1
X_09562_ _04186_ _04480_ vssd1 vssd1 vccd1 vccd1 _04481_ sky130_fd_sc_hd__and2_1
XANTENNA__09205__B _04053_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06774_ _01718_ _01722_ vssd1 vssd1 vccd1 vccd1 _01725_ sky130_fd_sc_hd__nand2_1
X_08513_ final_design.cpu.reg_window\[2\] final_design.cpu.reg_window\[34\] net832
+ vssd1 vssd1 vccd1 vccd1 _03464_ sky130_fd_sc_hd__mux2_1
XANTENNA__09920__S net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09493_ _04208_ _04210_ net467 vssd1 vssd1 vccd1 vccd1 _04412_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout256_A net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08444_ final_design.cpu.reg_window\[388\] final_design.cpu.reg_window\[420\] net821
+ vssd1 vssd1 vccd1 vccd1 _03395_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_95 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06845__A net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08059__B1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12058__S net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08375_ _03297_ _03322_ _02211_ vssd1 vssd1 vccd1 vccd1 _03326_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout423_A net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1165_A net1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07326_ final_design.cpu.reg_window\[4\] final_design.cpu.reg_window\[36\] net902
+ vssd1 vssd1 vccd1 vccd1 _02277_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_22_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_22_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06704__S1 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11897__S net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07257_ final_design.cpu.reg_window\[519\] final_design.cpu.reg_window\[551\] net887
+ vssd1 vssd1 vccd1 vccd1 _02208_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout309_X net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_871 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07188_ final_design.cpu.reg_window\[9\] final_design.cpu.reg_window\[41\] net888
+ vssd1 vssd1 vccd1 vccd1 _02139_ sky130_fd_sc_hd__mux2_1
XANTENNA__11366__B1 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout792_A net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08457__S1 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1745 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_6_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10614__A2_N net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout420 net421 vssd1 vssd1 vccd1 vccd1 net420 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_6_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout431 _05847_ vssd1 vssd1 vccd1 vccd1 net431 sky130_fd_sc_hd__buf_4
XANTENNA_fanout678_X net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11926__A net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout442 net443 vssd1 vssd1 vccd1 vccd1 net442 sky130_fd_sc_hd__clkbuf_4
Xfanout453 net454 vssd1 vssd1 vccd1 vccd1 net453 sky130_fd_sc_hd__buf_4
Xfanout464 _03519_ vssd1 vssd1 vccd1 vccd1 net464 sky130_fd_sc_hd__buf_2
Xfanout475 net476 vssd1 vssd1 vccd1 vccd1 net475 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_35_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout486 net488 vssd1 vssd1 vccd1 vccd1 net486 sky130_fd_sc_hd__buf_2
XANTENNA__12330__A2 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09829_ net726 _04744_ _04747_ vssd1 vssd1 vccd1 vccd1 _04748_ sky130_fd_sc_hd__o21a_1
XANTENNA__11645__B net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout497 _03418_ vssd1 vssd1 vccd1 vccd1 net497 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_31_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13940__CLK clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10341__B2 final_design.data_from_mem\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12840_ clknet_leaf_19_clk _00078_ net1111 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.ready_data\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_1347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07196__S1 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11722_ net434 net577 _06219_ net296 net1731 vssd1 vssd1 vccd1 vccd1 _00492_ sky130_fd_sc_hd__a32o_1
XFILLER_0_51_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07350__S net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06943__S1 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11653_ net190 net632 vssd1 vssd1 vccd1 vccd1 _06184_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_29_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10604_ _04961_ _04787_ vssd1 vssd1 vccd1 vccd1 _05348_ sky130_fd_sc_hd__and2b_1
X_11584_ net192 net637 vssd1 vssd1 vccd1 vccd1 _06148_ sky130_fd_sc_hd__and2_1
XFILLER_0_0_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13320__CLK clknet_leaf_41_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13323_ clknet_leaf_53_clk _00554_ net1189 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[311\]
+ sky130_fd_sc_hd__dfrtp_1
X_10535_ net62 _05282_ vssd1 vssd1 vccd1 vccd1 _05283_ sky130_fd_sc_hd__nand2_1
XFILLER_0_36_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1889 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13254_ clknet_leaf_50_clk _00485_ net1172 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[242\]
+ sky130_fd_sc_hd__dfrtp_1
X_10466_ net68 net958 net955 final_design.CPU_instr_adr\[0\] vssd1 vssd1 vccd1 vccd1
+ _05218_ sky130_fd_sc_hd__o22a_1
XFILLER_0_51_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10724__B _04613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11357__B1 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12205_ net556 _06133_ net503 net376 net2300 vssd1 vssd1 vccd1 vccd1 _00923_ sky130_fd_sc_hd__a32o_1
XFILLER_0_0_927 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_61_clk_X clknet_leaf_61_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13185_ clknet_leaf_47_clk _00416_ net1198 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[173\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13470__CLK clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10397_ _03648_ _05180_ vssd1 vssd1 vccd1 vccd1 _05181_ sky130_fd_sc_hd__or2_4
X_12136_ net237 net2408 net385 vssd1 vssd1 vccd1 vccd1 _00857_ sky130_fd_sc_hd__mux2_1
XANTENNA__09970__B1 _04119_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11109__B1 net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07981__C1 net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12067_ net573 _05898_ net508 net395 net1590 vssd1 vssd1 vccd1 vccd1 _00792_ sky130_fd_sc_hd__a32o_1
XANTENNA__09722__A0 net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11018_ final_design.CPU_instr_adr\[27\] _05239_ _05742_ net1056 vssd1 vssd1 vccd1
+ vccd1 _05743_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__07959__S0 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10332__B2 final_design.data_from_mem\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06649__B _01599_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12609__B1 net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12969_ clknet_leaf_15_clk _00207_ net1092 vssd1 vssd1 vccd1 vccd1 final_design.uart.bits_received\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06490_ final_design.cpu.reg_window\[798\] final_design.cpu.reg_window\[830\] net935
+ vssd1 vssd1 vccd1 vccd1 _01441_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_16_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08209__X _03160_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_2907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_2918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_14_clk_X clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08160_ final_design.cpu.reg_window\[79\] final_design.cpu.reg_window\[111\] net807
+ vssd1 vssd1 vccd1 vccd1 _03111_ sky130_fd_sc_hd__mux2_1
X_07111_ final_design.reqhand.instruction\[12\] net973 _02060_ vssd1 vssd1 vccd1 vccd1
+ _02062_ sky130_fd_sc_hd__o21a_1
XFILLER_0_67_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09695__B _04613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06698__S0 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08091_ final_design.cpu.reg_window\[332\] final_design.cpu.reg_window\[364\] net828
+ vssd1 vssd1 vccd1 vccd1 _03042_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11510__S net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13813__CLK clknet_leaf_57_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload30 clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 clkload30/X sky130_fd_sc_hd__clkbuf_8
Xclkload41 clknet_leaf_32_clk vssd1 vssd1 vccd1 vccd1 clkload41/Y sky130_fd_sc_hd__clkinv_16
X_07042_ _01989_ _01990_ _01991_ _01992_ net765 net786 vssd1 vssd1 vccd1 vccd1 _01993_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_24_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08091__S net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_29_clk_X clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07016__A1 net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12560__A2 net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08993_ net258 _03927_ net1016 vssd1 vssd1 vccd1 vccd1 _03929_ sky130_fd_sc_hd__a21o_1
XANTENNA__13963__CLK clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08598__Y _03549_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07944_ _01755_ net602 vssd1 vssd1 vccd1 vccd1 _02895_ sky130_fd_sc_hd__and2_1
XANTENNA__07435__S net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07875_ final_design.cpu.reg_window\[596\] final_design.cpu.reg_window\[628\] net867
+ vssd1 vssd1 vccd1 vccd1 _02826_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10323__B2 final_design.data_from_mem\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout373_A _06272_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09614_ net492 _04491_ _04227_ vssd1 vssd1 vccd1 vccd1 _04533_ sky130_fd_sc_hd__o21a_1
X_06826_ net754 _01776_ vssd1 vssd1 vccd1 vccd1 _01777_ sky130_fd_sc_hd__or2_1
XFILLER_0_17_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09545_ _02936_ net445 net443 _02932_ _04463_ vssd1 vssd1 vccd1 vccd1 _04464_ sky130_fd_sc_hd__o221a_1
X_06757_ final_design.cpu.reg_window\[919\] final_design.cpu.reg_window\[951\] net932
+ vssd1 vssd1 vccd1 vccd1 _01708_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout540_A _02026_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout638_A net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout259_X net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09476_ _04393_ _04394_ net475 vssd1 vssd1 vccd1 vccd1 _04395_ sky130_fd_sc_hd__mux2_1
X_06688_ final_design.cpu.reg_window\[25\] final_design.cpu.reg_window\[57\] net936
+ vssd1 vssd1 vccd1 vccd1 _01639_ sky130_fd_sc_hd__mux2_1
XANTENNA__13343__CLK clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09492__A2 net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08427_ final_design.cpu.reg_window\[709\] final_design.cpu.reg_window\[741\] net840
+ vssd1 vssd1 vccd1 vccd1 _03378_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_1891 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout426_X net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout805_A _02095_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08358_ net707 _03302_ net722 vssd1 vssd1 vccd1 vccd1 _03309_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_24_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload2 clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 clkload2/Y sky130_fd_sc_hd__clkinvlp_4
XTAP_TAPCELL_ROW_43_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11587__B1 net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07309_ final_design.cpu.reg_window\[581\] final_design.cpu.reg_window\[613\] net921
+ vssd1 vssd1 vccd1 vccd1 _02260_ sky130_fd_sc_hd__mux2_1
XANTENNA__08452__B1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08289_ final_design.cpu.reg_window\[9\] final_design.cpu.reg_window\[41\] net807
+ vssd1 vssd1 vccd1 vccd1 _03240_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_1829 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13493__CLK clknet_leaf_56_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11420__S net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10320_ net1511 net1012 net988 final_design.data_from_mem\[5\] vssd1 vssd1 vccd1
+ vccd1 _00077_ sky130_fd_sc_hd__a22o_1
XFILLER_0_28_1640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout795_X net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10251_ _05119_ _05120_ vssd1 vssd1 vccd1 vccd1 _00015_ sky130_fd_sc_hd__nor2_1
XFILLER_0_63_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12551__A2 net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10182_ _05069_ _05071_ vssd1 vssd1 vccd1 vccd1 _05072_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout962_X net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10562__B2 net1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1204 net1227 vssd1 vssd1 vccd1 vccd1 net1204 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_37_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1215 net1217 vssd1 vssd1 vccd1 vccd1 net1215 sky130_fd_sc_hd__clkbuf_4
Xfanout1226 net1227 vssd1 vssd1 vccd1 vccd1 net1226 sky130_fd_sc_hd__clkbuf_2
Xfanout1237 net1244 vssd1 vssd1 vccd1 vccd1 net1237 sky130_fd_sc_hd__buf_2
Xfanout250 net251 vssd1 vssd1 vccd1 vccd1 net250 sky130_fd_sc_hd__buf_4
Xfanout261 _04071_ vssd1 vssd1 vccd1 vccd1 net261 sky130_fd_sc_hd__clkbuf_4
Xfanout272 net273 vssd1 vssd1 vccd1 vccd1 net272 sky130_fd_sc_hd__buf_4
XFILLER_0_76_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13941_ clknet_leaf_57_clk _01172_ net1144 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[929\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout283 net284 vssd1 vssd1 vccd1 vccd1 net283 sky130_fd_sc_hd__clkbuf_4
Xfanout294 net295 vssd1 vssd1 vccd1 vccd1 net294 sky130_fd_sc_hd__buf_4
XANTENNA__06613__S0 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13872_ clknet_leaf_34_clk _01103_ net1239 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[860\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07191__B1 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12067__A1 net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12823_ net1370 vssd1 vssd1 vccd1 vccd1 _00264_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__08684__B net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12754_ _06344_ _06351_ _06384_ vssd1 vssd1 vccd1 vccd1 _06391_ sky130_fd_sc_hd__or3_1
XFILLER_0_16_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06485__A net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09483__A2 net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06916__S1 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11705_ net204 net629 vssd1 vssd1 vccd1 vccd1 _06211_ sky130_fd_sc_hd__and2_1
XANTENNA__11290__A2 _05984_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12685_ final_design.VGA_data_control.ready_data\[30\] net1022 net977 final_design.data_from_mem\[30\]
+ vssd1 vssd1 vccd1 vccd1 _06330_ sky130_fd_sc_hd__a22o_1
XFILLER_0_38_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13836__CLK clknet_leaf_46_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11636_ net426 net556 _06175_ net298 net1497 vssd1 vssd1 vccd1 vccd1 _00450_ sky130_fd_sc_hd__a32o_1
XFILLER_0_38_996 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11567_ net559 net421 _06139_ net302 net1738 vssd1 vssd1 vccd1 vccd1 _00417_ sky130_fd_sc_hd__a32o_1
X_10518_ net1427 net1029 net1002 _05266_ vssd1 vssd1 vccd1 vccd1 _00176_ sky130_fd_sc_hd__a22o_1
XANTENNA__07341__S1 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13306_ clknet_leaf_6_clk _00537_ net1128 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[294\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold709 final_design.cpu.reg_window\[951\] vssd1 vssd1 vccd1 vccd1 net2051 sky130_fd_sc_hd__dlygate4sd3_1
Xwire695 _01753_ vssd1 vssd1 vccd1 vccd1 net695 sky130_fd_sc_hd__buf_4
X_11498_ net673 _06116_ vssd1 vssd1 vccd1 vccd1 _06117_ sky130_fd_sc_hd__nand2_1
XANTENNA__12860__CLK clknet_leaf_18_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10454__B net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13986__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13237_ clknet_leaf_6_clk _00468_ net1133 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[225\]
+ sky130_fd_sc_hd__dfrtp_1
X_10449_ net1426 net1035 _05208_ net248 vssd1 vssd1 vccd1 vccd1 _00165_ sky130_fd_sc_hd__a22o_1
XANTENNA__09538__A3 net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12542__A2 net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09943__B1 net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13168_ clknet_leaf_33_clk _00399_ net1231 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[156\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11750__A0 net207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12119_ net1995 net190 net391 vssd1 vssd1 vccd1 vccd1 _00843_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_41_clk_A clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11566__A net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13216__CLK clknet_leaf_11_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1913 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12161__S net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13099_ clknet_leaf_38_clk _00330_ net1188 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[87\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07255__S net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07108__X _02059_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07660_ _01507_ net604 vssd1 vssd1 vccd1 vccd1 _02611_ sky130_fd_sc_hd__nand2_1
XANTENNA__13366__CLK clknet_leaf_58_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_56_clk_A clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06611_ final_design.cpu.reg_window\[604\] final_design.cpu.reg_window\[636\] net947
+ vssd1 vssd1 vccd1 vccd1 _01562_ sky130_fd_sc_hd__mux2_1
XANTENNA__12058__A1 net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07591_ net602 _02540_ _02515_ _02503_ vssd1 vssd1 vccd1 vccd1 _02542_ sky130_fd_sc_hd__o211a_2
X_09330_ _01493_ _04248_ vssd1 vssd1 vccd1 vccd1 _04249_ sky130_fd_sc_hd__or2_2
XANTENNA__11505__S net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06542_ _01463_ _01474_ _01482_ vssd1 vssd1 vccd1 vccd1 _01493_ sky130_fd_sc_hd__or3_4
XFILLER_0_14_1717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10629__B final_design.VGA_adr\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09474__A2 net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09261_ net96 net97 _04179_ vssd1 vssd1 vccd1 vccd1 _04180_ sky130_fd_sc_hd__and3_1
XFILLER_0_8_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06473_ final_design.cpu.reg_window\[286\] final_design.cpu.reg_window\[318\] net932
+ vssd1 vssd1 vccd1 vccd1 _01424_ sky130_fd_sc_hd__mux2_1
X_08212_ net600 _03160_ _03135_ net541 vssd1 vssd1 vccd1 vccd1 _03163_ sky130_fd_sc_hd__o211a_1
XFILLER_0_12_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09192_ _03617_ _03649_ vssd1 vssd1 vccd1 vccd1 _04111_ sky130_fd_sc_hd__nor2_2
XFILLER_0_62_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11569__B1 net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08143_ _03090_ _03091_ _03092_ _03093_ net684 net703 vssd1 vssd1 vccd1 vccd1 _03094_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_44_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout219_A _05928_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08074_ net613 _03022_ _03023_ net547 vssd1 vssd1 vccd1 vccd1 _03025_ sky130_fd_sc_hd__a211oi_2
X_07025_ final_design.cpu.reg_window\[206\] final_design.cpu.reg_window\[238\] net893
+ vssd1 vssd1 vccd1 vccd1 _01976_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout1030_A net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12533__A2 net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09934__B1 net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1879 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11741__A0 net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout490_A _03453_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout588_A net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14141__CLK clknet_leaf_19_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold14 final_design.cpu.reg_window\[2\] vssd1 vssd1 vccd1 vccd1 net1356 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_32_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08976_ _01911_ _01912_ vssd1 vssd1 vccd1 vccd1 _03913_ sky130_fd_sc_hd__and2b_1
XANTENNA__12985__RESET_B net1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold25 final_design.cpu.reg_window\[17\] vssd1 vssd1 vccd1 vccd1 net1367 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_32_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold36 final_design.cpu.reg_window\[19\] vssd1 vssd1 vccd1 vccd1 net1378 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07165__S net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold47 net171 vssd1 vssd1 vccd1 vccd1 net1389 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_51_1955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13709__CLK clknet_leaf_48_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07927_ final_design.cpu.reg_window\[214\] final_design.cpu.reg_window\[246\] net837
+ vssd1 vssd1 vccd1 vccd1 _02878_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_51_1966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12297__A1 net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold58 final_design.reqhand.instruction\[21\] vssd1 vssd1 vccd1 vccd1 net1400 sky130_fd_sc_hd__dlygate4sd3_1
Xhold69 net103 vssd1 vssd1 vccd1 vccd1 net1411 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout755_A net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout376_X net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08596__S0 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07858_ final_design.cpu.reg_window\[404\] final_design.cpu.reg_window\[436\] net868
+ vssd1 vssd1 vccd1 vccd1 _02809_ sky130_fd_sc_hd__mux2_1
XANTENNA__12049__A1 net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06809_ final_design.cpu.reg_window\[213\] final_design.cpu.reg_window\[245\] net939
+ vssd1 vssd1 vccd1 vccd1 _01760_ sky130_fd_sc_hd__mux2_1
X_07789_ final_design.cpu.reg_window\[345\] final_design.cpu.reg_window\[377\] net856
+ vssd1 vssd1 vccd1 vccd1 _02740_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout922_A net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11415__S net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09528_ _04436_ _04446_ vssd1 vssd1 vccd1 vccd1 _04447_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_49_1873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_1884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09459_ _04107_ _04377_ _04376_ net481 vssd1 vssd1 vccd1 vccd1 _04378_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA_fanout710_X net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09870__C1 _04046_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12470_ _06130_ net348 net331 net2224 vssd1 vssd1 vccd1 vccd1 _01176_ sky130_fd_sc_hd__a22o_1
XFILLER_0_30_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12883__CLK clknet_leaf_18_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11421_ net1972 net215 net311 vssd1 vssd1 vccd1 vccd1 _00318_ sky130_fd_sc_hd__mux2_1
XANTENNA__12221__A1 net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1773 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14140_ clknet_leaf_17_clk net1246 net1115 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.h_count\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_50_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11352_ final_design.data_from_mem\[25\] net235 net233 vssd1 vssd1 vccd1 vccd1 _06042_
+ sky130_fd_sc_hd__a21o_2
X_10303_ final_design.VGA_data_control.h_count\[3\] _05156_ final_design.VGA_data_control.h_count\[5\]
+ vssd1 vssd1 vccd1 vccd1 _05157_ sky130_fd_sc_hd__o21ai_1
XANTENNA__10783__B2 net1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11980__B1 net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13239__CLK clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14071_ clknet_leaf_13_clk _01268_ net1106 vssd1 vssd1 vccd1 vccd1 final_design.uart.working_data\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_11283_ net432 net572 _05981_ net317 net1699 vssd1 vssd1 vccd1 vccd1 _00291_ sky130_fd_sc_hd__a32o_1
X_13022_ clknet_leaf_13_clk _00253_ net1088 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input51_A mem_adr_start[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10234_ final_design.uart.BAUD_counter\[12\] _05108_ net799 vssd1 vssd1 vccd1 vccd1
+ _05110_ sky130_fd_sc_hd__o21ai_1
XANTENNA__12524__A2 net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07087__S0 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06739__B1 _01504_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11732__B1 net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1001 _05239_ vssd1 vssd1 vccd1 vccd1 net1001 sky130_fd_sc_hd__buf_4
Xfanout1012 _05166_ vssd1 vssd1 vccd1 vccd1 net1012 sky130_fd_sc_hd__clkbuf_2
X_10165_ _05058_ vssd1 vssd1 vccd1 vccd1 _05059_ sky130_fd_sc_hd__inv_2
Xfanout1023 net1024 vssd1 vssd1 vccd1 vccd1 net1023 sky130_fd_sc_hd__clkbuf_4
Xfanout1034 net1035 vssd1 vssd1 vccd1 vccd1 net1034 sky130_fd_sc_hd__clkbuf_2
Xfanout1045 net1047 vssd1 vssd1 vccd1 vccd1 net1045 sky130_fd_sc_hd__clkbuf_2
XANTENNA__13389__CLK clknet_leaf_44_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1056 final_design.reqhand.current_client\[2\] vssd1 vssd1 vccd1 vccd1 net1056
+ sky130_fd_sc_hd__buf_4
XANTENNA__12288__A1 net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10096_ final_design.VGA_data_control.h_count\[0\] net1050 vssd1 vssd1 vccd1 vccd1
+ _05012_ sky130_fd_sc_hd__or2_1
Xfanout1067 net1068 vssd1 vssd1 vccd1 vccd1 net1067 sky130_fd_sc_hd__buf_2
Xfanout1078 net1080 vssd1 vssd1 vccd1 vccd1 net1078 sky130_fd_sc_hd__buf_2
XFILLER_0_76_1733 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1089 net1090 vssd1 vssd1 vccd1 vccd1 net1089 sky130_fd_sc_hd__buf_2
X_13924_ clknet_leaf_52_clk _01155_ net1171 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[912\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06767__X _01718_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1777 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13855_ clknet_leaf_7_clk _01086_ net1130 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[843\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_18_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12806_ net1383 vssd1 vssd1 vccd1 vccd1 _00247_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__11552__C net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10998_ _05722_ _05723_ vssd1 vssd1 vccd1 vccd1 _05724_ sky130_fd_sc_hd__or2_1
XFILLER_0_70_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13786_ clknet_leaf_58_clk _01017_ net1122 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[774\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_8_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12737_ _05058_ _06373_ _06376_ vssd1 vssd1 vccd1 vccd1 _06378_ sky130_fd_sc_hd__a21o_1
XANTENNA__11263__A2 _05960_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10471__B1 net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_2284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_2295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12668_ _06321_ net1464 net978 vssd1 vssd1 vccd1 vccd1 _01336_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14014__CLK clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11619_ net243 net630 vssd1 vssd1 vccd1 vccd1 _06167_ sky130_fd_sc_hd__and2_1
XANTENNA__12156__S net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12599_ net1403 net996 net982 final_design.data_from_mem\[17\] vssd1 vssd1 vccd1
+ vccd1 _01292_ sky130_fd_sc_hd__a22o_1
XFILLER_0_53_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08511__S0 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07110__Y _02061_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold506 final_design.cpu.reg_window\[465\] vssd1 vssd1 vccd1 vccd1 net1848 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11971__B1 net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold517 final_design.cpu.reg_window\[594\] vssd1 vssd1 vccd1 vccd1 net1859 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold528 final_design.cpu.reg_window\[660\] vssd1 vssd1 vccd1 vccd1 net1870 sky130_fd_sc_hd__dlygate4sd3_1
Xhold539 final_design.cpu.reg_window\[542\] vssd1 vssd1 vccd1 vccd1 net1881 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14164__CLK clknet_leaf_17_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12515__A2 net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_2077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_2088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_2099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08830_ _03779_ _03780_ vssd1 vssd1 vccd1 vccd1 _03781_ sky130_fd_sc_hd__xnor2_1
XANTENNA__06825__S0 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1206 final_design.cpu.reg_window\[818\] vssd1 vssd1 vccd1 vccd1 net2548 sky130_fd_sc_hd__dlygate4sd3_1
X_08761_ _01367_ _02361_ vssd1 vssd1 vccd1 vccd1 _03712_ sky130_fd_sc_hd__nor2_1
XFILLER_0_75_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07712_ final_design.cpu.reg_window\[795\] final_design.cpu.reg_window\[827\] net863
+ vssd1 vssd1 vccd1 vccd1 _02663_ sky130_fd_sc_hd__mux2_1
XANTENNA__08578__S0 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07780__Y _02731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08692_ _03456_ _03457_ _03554_ _03639_ vssd1 vssd1 vccd1 vccd1 _03643_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_0_203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07713__S net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07643_ _02590_ _02591_ _02592_ _02593_ net687 net704 vssd1 vssd1 vccd1 vccd1 _02594_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__06902__B1 _01821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_96 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07574_ final_design.cpu.reg_window\[159\] final_design.cpu.reg_window\[191\] net857
+ vssd1 vssd1 vccd1 vccd1 _02525_ sky130_fd_sc_hd__mux2_1
X_09313_ net541 net540 net539 _02091_ net459 net469 vssd1 vssd1 vccd1 vccd1 _04232_
+ sky130_fd_sc_hd__mux4_1
X_06525_ _01465_ _01468_ _01475_ vssd1 vssd1 vccd1 vccd1 _01476_ sky130_fd_sc_hd__nor3_2
XANTENNA__11254__A2 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout336_A net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_60_clk clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_60_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_8_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09244_ _04162_ vssd1 vssd1 vccd1 vccd1 _04163_ sky130_fd_sc_hd__inv_2
XFILLER_0_75_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06456_ _01405_ _01406_ _01407_ _01396_ vssd1 vssd1 vccd1 vccd1 _01409_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_8_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08544__S net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12203__A1 net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09175_ _03631_ _03650_ vssd1 vssd1 vccd1 vccd1 _04094_ sky130_fd_sc_hd__nor2_4
XFILLER_0_66_1913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout503_A net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1245_A net100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08126_ _03073_ _03074_ _03075_ _03076_ net684 net694 vssd1 vssd1 vccd1 vccd1 _03077_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_32_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11962__B1 net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_1_Right_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08057_ _03004_ _03005_ _03006_ _03007_ net682 net702 vssd1 vssd1 vccd1 vccd1 _03008_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout1033_X net1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07008_ _01955_ _01956_ _01957_ _01958_ net766 net785 vssd1 vssd1 vccd1 vccd1 _01959_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__12506__A2 net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11918__B _05845_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout493_X net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout872_A net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11714__B1 net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09383__A1 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11190__A1 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout660_X net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08959_ _02459_ _03897_ vssd1 vssd1 vccd1 vccd1 _03898_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout758_X net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13681__CLK clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11970_ _06172_ net279 net404 net1832 vssd1 vssd1 vccd1 vccd1 _00703_ sky130_fd_sc_hd__a22o_1
XFILLER_0_73_1917 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10921_ net83 net1046 vssd1 vssd1 vccd1 vccd1 _05650_ sky130_fd_sc_hd__and2_1
XANTENNA__07241__S0 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11653__B net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10852_ _04954_ net252 vssd1 vssd1 vccd1 vccd1 _05584_ sky130_fd_sc_hd__nor2_1
X_13640_ clknet_leaf_40_clk _00871_ net1219 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[628\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14037__CLK clknet_leaf_15_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10783_ final_design.CPU_instr_adr\[16\] net1000 _05516_ net1042 vssd1 vssd1 vccd1
+ vccd1 _05519_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_67_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13571_ clknet_leaf_0_clk _00802_ net1062 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[559\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12442__A1 net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12765__A final_design.VGA_adr\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_51_clk clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_51_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_52_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_1901 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12522_ _06184_ net355 net329 net1861 vssd1 vssd1 vccd1 vccd1 _01227_ sky130_fd_sc_hd__a22o_1
XFILLER_0_82_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08454__S net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input99_A memory_size[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13061__CLK clknet_leaf_49_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12453_ net1721 net196 net337 vssd1 vssd1 vccd1 vccd1 _01160_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11404_ _04127_ _04176_ net657 vssd1 vssd1 vccd1 vccd1 _06088_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_10_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12384_ net1706 net197 net270 vssd1 vssd1 vccd1 vccd1 _01095_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_10_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10300__S0 net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11953__B1 net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14123_ clknet_leaf_21_clk final_design.vga.v_next_count\[3\] net1159 vssd1 vssd1
+ vccd1 vccd1 final_design.VGA_data_control.v_count\[3\] sky130_fd_sc_hd__dfrtp_2
X_11335_ net737 _03869_ _06026_ vssd1 vssd1 vccd1 vccd1 _06027_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_1_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14054_ clknet_leaf_16_clk _00015_ net1091 vssd1 vssd1 vccd1 vccd1 final_design.uart.BAUD_counter\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_11266_ net2506 net314 _05966_ net425 vssd1 vssd1 vccd1 vccd1 _00289_ sky130_fd_sc_hd__a22o_1
XFILLER_0_43_1743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13005_ net1336 _00236_ net1233 vssd1 vssd1 vccd1 vccd1 final_design.CPU_instr_adr\[25\]
+ sky130_fd_sc_hd__dfrtp_2
X_10217_ final_design.uart.BAUD_counter\[6\] _05098_ vssd1 vssd1 vccd1 vccd1 _05099_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_43_1776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11197_ net427 net563 _05905_ net315 net1983 vssd1 vssd1 vccd1 vccd1 _00281_ sky130_fd_sc_hd__a32o_1
XANTENNA__11181__A1 net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10148_ _05012_ _05046_ _05047_ vssd1 vssd1 vccd1 vccd1 final_design.vga.h_next_count\[1\]
+ sky130_fd_sc_hd__and3_1
XFILLER_0_59_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10079_ net1 _04995_ _04993_ vssd1 vssd1 vccd1 vccd1 _00003_ sky130_fd_sc_hd__a21o_1
XANTENNA__07533__S net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13907_ clknet_leaf_36_clk _01138_ net1230 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[895\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_8_1913 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12681__B2 final_design.data_from_mem\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_2482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13838_ clknet_leaf_45_clk _01069_ net1216 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[826\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09429__A2 _04343_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_2346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_63_2357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_2368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13769_ clknet_leaf_36_clk _01000_ net1229 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[757\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_42_clk clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_42_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__13404__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07290_ _02239_ _02240_ vssd1 vssd1 vccd1 vccd1 _02241_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_45_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12197__A0 net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13554__CLK clknet_leaf_39_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09601__A2 _04088_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_2139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold303 final_design.cpu.reg_window\[902\] vssd1 vssd1 vccd1 vccd1 net1645 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11944__B1 net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold314 final_design.cpu.reg_window\[968\] vssd1 vssd1 vccd1 vccd1 net1656 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold325 final_design.cpu.reg_window\[37\] vssd1 vssd1 vccd1 vccd1 net1667 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_766 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12614__S _05080_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold336 final_design.cpu.reg_window\[66\] vssd1 vssd1 vccd1 vccd1 net1678 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold347 final_design.cpu.reg_window\[42\] vssd1 vssd1 vccd1 vccd1 net1689 sky130_fd_sc_hd__dlygate4sd3_1
Xhold358 final_design.cpu.reg_window\[535\] vssd1 vssd1 vccd1 vccd1 net1700 sky130_fd_sc_hd__dlygate4sd3_1
X_09931_ net95 _04178_ vssd1 vssd1 vccd1 vccd1 _04850_ sky130_fd_sc_hd__nor2_1
Xhold369 final_design.cpu.reg_window\[554\] vssd1 vssd1 vccd1 vccd1 net1711 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout805 _02095_ vssd1 vssd1 vccd1 vccd1 net805 sky130_fd_sc_hd__buf_2
Xfanout816 net817 vssd1 vssd1 vccd1 vccd1 net816 sky130_fd_sc_hd__clkbuf_4
X_09862_ net482 _04683_ _04780_ _04055_ vssd1 vssd1 vccd1 vccd1 _04781_ sky130_fd_sc_hd__a211o_1
Xfanout827 net828 vssd1 vssd1 vccd1 vccd1 net827 sky130_fd_sc_hd__buf_2
Xfanout838 net841 vssd1 vssd1 vccd1 vccd1 net838 sky130_fd_sc_hd__clkbuf_4
Xfanout849 net852 vssd1 vssd1 vccd1 vccd1 net849 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07915__A2 _02863_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08813_ final_design.CPU_instr_adr\[20\] _01823_ _03760_ vssd1 vssd1 vccd1 vccd1
+ _03764_ sky130_fd_sc_hd__a21bo_1
Xhold1003 final_design.cpu.reg_window\[285\] vssd1 vssd1 vccd1 vccd1 net2345 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09770__D1 net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1014 final_design.cpu.reg_window\[630\] vssd1 vssd1 vccd1 vccd1 net2356 sky130_fd_sc_hd__dlygate4sd3_1
X_09793_ _04710_ _04711_ net476 vssd1 vssd1 vccd1 vccd1 _04712_ sky130_fd_sc_hd__mux2_1
Xhold1025 final_design.cpu.reg_window\[625\] vssd1 vssd1 vccd1 vccd1 net2367 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1036 final_design.cpu.reg_window\[617\] vssd1 vssd1 vccd1 vccd1 net2378 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout286_A net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1047 final_design.cpu.reg_window\[628\] vssd1 vssd1 vccd1 vccd1 net2389 sky130_fd_sc_hd__dlygate4sd3_1
X_08744_ final_design.CPU_instr_adr\[9\] net667 _01537_ vssd1 vssd1 vccd1 vccd1 _03695_
+ sky130_fd_sc_hd__and3_1
Xhold1058 final_design.cpu.reg_window\[355\] vssd1 vssd1 vccd1 vccd1 net2400 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07128__B1 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1069 final_design.cpu.reg_window\[563\] vssd1 vssd1 vccd1 vccd1 net2411 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08675_ _02061_ _03616_ _01487_ vssd1 vssd1 vccd1 vccd1 _03626_ sky130_fd_sc_hd__a21o_1
XFILLER_0_75_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout453_A net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1195_A net1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10683__B1 net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07626_ _01570_ net607 vssd1 vssd1 vccd1 vccd1 _02577_ sky130_fd_sc_hd__nand2_1
XFILLER_0_18_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07557_ _02477_ _02505_ vssd1 vssd1 vccd1 vccd1 _02508_ sky130_fd_sc_hd__xnor2_1
XANTENNA__13084__CLK clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout620_A _02507_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout339_X net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout718_A _01720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_33_clk clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_33_clk sky130_fd_sc_hd__clkbuf_8
X_06508_ net1040 net995 net992 final_design.reqhand.instruction\[4\] vssd1 vssd1 vccd1
+ vccd1 _01459_ sky130_fd_sc_hd__o31a_1
XANTENNA__10435__B1 _05201_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06583__A net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07488_ _02214_ _02437_ _02213_ vssd1 vssd1 vccd1 vccd1 _02439_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_64_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06439_ wb_manage.BUSY_O net34 vssd1 vssd1 vccd1 vccd1 _01393_ sky130_fd_sc_hd__and2b_1
X_09227_ _03488_ _04145_ _03486_ vssd1 vssd1 vccd1 vccd1 _04146_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout1150_X net1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout506_X net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_1721 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09158_ _04075_ _04076_ net478 vssd1 vssd1 vccd1 vccd1 _04077_ sky130_fd_sc_hd__mux2_1
XANTENNA__09053__B1 net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06870__X _01821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10738__A1 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11935__B1 net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08109_ final_design.cpu.reg_window\[652\] final_design.cpu.reg_window\[684\] net813
+ vssd1 vssd1 vccd1 vccd1 _03060_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09089_ _02300_ _02433_ _04012_ vssd1 vssd1 vccd1 vccd1 _04013_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_82_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12921__CLK clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07618__S net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11120_ _05831_ _05835_ _05836_ _05830_ net2537 vssd1 vssd1 vccd1 vccd1 _00208_ sky130_fd_sc_hd__a32o_1
Xhold870 final_design.cpu.reg_window\[955\] vssd1 vssd1 vccd1 vccd1 net2212 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout875_X net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold881 final_design.cpu.reg_window\[271\] vssd1 vssd1 vccd1 vccd1 net2223 sky130_fd_sc_hd__dlygate4sd3_1
X_11051_ _05773_ _05774_ vssd1 vssd1 vccd1 vccd1 _05775_ sky130_fd_sc_hd__or2_1
Xhold892 final_design.cpu.reg_window\[632\] vssd1 vssd1 vccd1 vccd1 net2234 sky130_fd_sc_hd__dlygate4sd3_1
X_10002_ _04192_ _04920_ vssd1 vssd1 vccd1 vccd1 _04921_ sky130_fd_sc_hd__and2_1
XANTENNA__12360__B1 net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08449__S net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1861 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07353__S net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input14_A DAT_I[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11953_ _06154_ net292 net410 net2522 vssd1 vssd1 vccd1 vccd1 _00688_ sky130_fd_sc_hd__a22o_1
XFILLER_0_59_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12663__B2 final_design.data_from_mem\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13427__CLK clknet_leaf_39_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10904_ _05633_ _05629_ vssd1 vssd1 vccd1 vccd1 _05634_ sky130_fd_sc_hd__and2b_1
XFILLER_0_54_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11884_ _05848_ _06246_ vssd1 vssd1 vccd1 vccd1 _06247_ sky130_fd_sc_hd__or2_1
X_13623_ clknet_leaf_4_clk _00854_ net1084 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[611\]
+ sky130_fd_sc_hd__dfrtp_1
X_10835_ net78 net1044 vssd1 vssd1 vccd1 vccd1 _05568_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_81_2980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_24_clk clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_24_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_67_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09292__A0 _01626_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13554_ clknet_leaf_39_clk _00785_ net1205 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[542\]
+ sky130_fd_sc_hd__dfrtp_1
X_10766_ _05439_ _05501_ vssd1 vssd1 vccd1 vccd1 _05502_ sky130_fd_sc_hd__nor2_1
XFILLER_0_66_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13577__CLK clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12505_ _06167_ net342 net326 net2095 vssd1 vssd1 vccd1 vccd1 _01210_ sky130_fd_sc_hd__a22o_1
X_10697_ net39 _05435_ vssd1 vssd1 vccd1 vccd1 _05437_ sky130_fd_sc_hd__nor2_1
XFILLER_0_67_1529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13485_ clknet_leaf_44_clk _00716_ net1202 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[473\]
+ sky130_fd_sc_hd__dfrtp_1
X_12436_ net1608 net240 net334 vssd1 vssd1 vccd1 vccd1 _01143_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_2751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_2762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12434__S net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12367_ net1754 net227 net269 vssd1 vssd1 vccd1 vccd1 _01078_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_75_2773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_2615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14106_ clknet_leaf_23_clk _01303_ net1164 vssd1 vssd1 vccd1 vccd1 final_design.reqhand.instruction\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_71_2626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11318_ net663 _03882_ net737 vssd1 vssd1 vccd1 vccd1 _06012_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11558__B net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_2637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12298_ net2210 net229 net365 vssd1 vssd1 vccd1 vccd1 _01012_ sky130_fd_sc_hd__mux2_1
XANTENNA__10462__B net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14037_ clknet_leaf_15_clk _00017_ net1092 vssd1 vssd1 vccd1 vccd1 final_design.uart.BAUD_counter\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_11249_ net646 net212 vssd1 vssd1 vccd1 vccd1 _05952_ sky130_fd_sc_hd__and2_2
XANTENNA__12351__B1 net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06790_ final_design.cpu.reg_window\[662\] final_design.cpu.reg_window\[694\] net920
+ vssd1 vssd1 vccd1 vccd1 _01741_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_1901 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_2555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06668__A net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13876__RESET_B net1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_2566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_2577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_2419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10665__B1 _04990_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08460_ final_design.cpu.reg_window\[580\] final_design.cpu.reg_window\[612\] net819
+ vssd1 vssd1 vccd1 vccd1 _03411_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07411_ net528 _02361_ vssd1 vssd1 vccd1 vccd1 _02362_ sky130_fd_sc_hd__nor2_1
XFILLER_0_37_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08391_ final_design.cpu.reg_window\[774\] final_design.cpu.reg_window\[806\] net831
+ vssd1 vssd1 vccd1 vccd1 _03342_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_15_clk clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_15_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__11513__S net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07342_ _02287_ _02292_ net749 vssd1 vssd1 vccd1 vccd1 _02293_ sky130_fd_sc_hd__mux2_1
XANTENNA__08094__S net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07273_ final_design.cpu.reg_window\[70\] final_design.cpu.reg_window\[102\] net904
+ vssd1 vssd1 vccd1 vccd1 _02224_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_14_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12944__CLK clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09012_ _02032_ _02033_ vssd1 vssd1 vccd1 vccd1 _03945_ sky130_fd_sc_hd__and2b_1
XFILLER_0_2_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_40 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold100 final_design.reqhand.instruction\[28\] vssd1 vssd1 vccd1 vccd1 net1442 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_78_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout201_A _05996_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold111 net139 vssd1 vssd1 vccd1 vccd1 net1453 sky130_fd_sc_hd__dlygate4sd3_1
Xhold122 final_design.VGA_data_control.data_to_VGA\[21\] vssd1 vssd1 vccd1 vccd1 net1464
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold133 final_design.cpu.reg_window\[194\] vssd1 vssd1 vccd1 vccd1 net1475 sky130_fd_sc_hd__dlygate4sd3_1
Xhold144 final_design.cpu.reg_window\[214\] vssd1 vssd1 vccd1 vccd1 net1486 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12590__B1 net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11468__B net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold155 final_design.cpu.reg_window\[207\] vssd1 vssd1 vccd1 vccd1 net1497 sky130_fd_sc_hd__dlygate4sd3_1
Xhold166 final_design.VGA_data_control.ready_data\[30\] vssd1 vssd1 vccd1 vccd1 net1508
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_61_1640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold177 final_design.VGA_data_control.ready_data\[16\] vssd1 vssd1 vccd1 vccd1 net1519
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold188 final_design.VGA_data_control.data_to_VGA\[13\] vssd1 vssd1 vccd1 vccd1 net1530
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold199 final_design.cpu.reg_window\[712\] vssd1 vssd1 vccd1 vccd1 net1541 sky130_fd_sc_hd__dlygate4sd3_1
X_09914_ _03422_ net441 net438 _03421_ _04832_ vssd1 vssd1 vccd1 vccd1 _04833_ sky130_fd_sc_hd__o221a_1
Xfanout602 net603 vssd1 vssd1 vccd1 vccd1 net602 sky130_fd_sc_hd__buf_2
Xfanout613 net618 vssd1 vssd1 vccd1 vccd1 net613 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_0_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11145__A1 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout624 net625 vssd1 vssd1 vccd1 vccd1 net624 sky130_fd_sc_hd__buf_2
Xfanout635 _06123_ vssd1 vssd1 vccd1 vccd1 net635 sky130_fd_sc_hd__clkbuf_8
XANTENNA__12342__B1 net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout646 net648 vssd1 vssd1 vccd1 vccd1 net646 sky130_fd_sc_hd__clkbuf_4
XANTENNA_input6_A DAT_I[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08010__B2 net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09845_ _03229_ _04503_ vssd1 vssd1 vccd1 vccd1 _04764_ sky130_fd_sc_hd__or2_1
Xfanout657 net658 vssd1 vssd1 vccd1 vccd1 net657 sky130_fd_sc_hd__clkbuf_2
Xfanout668 net670 vssd1 vssd1 vccd1 vccd1 net668 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout570_A net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout679 net681 vssd1 vssd1 vccd1 vccd1 net679 sky130_fd_sc_hd__buf_4
XANTENNA_fanout668_A net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout289_X net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09776_ _04409_ _04694_ _04689_ vssd1 vssd1 vccd1 vccd1 _04695_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_20_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06988_ net743 net667 net664 net773 _01821_ vssd1 vssd1 vccd1 vccd1 _01939_ sky130_fd_sc_hd__o221a_2
XFILLER_0_9_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08727_ _01939_ final_design.CPU_instr_adr\[16\] vssd1 vssd1 vccd1 vccd1 _03678_
+ sky130_fd_sc_hd__and2b_1
XANTENNA__12645__B2 final_design.data_from_mem\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout835_A net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10656__B1 net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08658_ _02642_ _03607_ _03608_ _02545_ _03604_ vssd1 vssd1 vccd1 vccd1 _03609_ sky130_fd_sc_hd__a221oi_2
X_07609_ final_design.cpu.reg_window\[541\] final_design.cpu.reg_window\[573\] net866
+ vssd1 vssd1 vccd1 vccd1 _02560_ sky130_fd_sc_hd__mux2_1
XANTENNA__06584__Y _01535_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08589_ final_design.cpu.reg_window\[896\] final_design.cpu.reg_window\[928\] net827
+ vssd1 vssd1 vccd1 vccd1 _03540_ sky130_fd_sc_hd__mux2_1
XANTENNA__11423__S net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10620_ _05362_ _05363_ vssd1 vssd1 vccd1 vccd1 _05364_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_12_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09813__A2 net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_12_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10551_ _04042_ _05296_ _05297_ _05295_ net960 vssd1 vssd1 vccd1 vccd1 _05298_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_12_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11620__A2 net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10482_ _05231_ _05232_ net1470 net1030 vssd1 vssd1 vccd1 vccd1 _00174_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__09026__B1 net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13270_ clknet_leaf_57_clk _00501_ net1138 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[258\]
+ sky130_fd_sc_hd__dfrtp_1
X_12221_ net582 _06149_ net514 net378 net1947 vssd1 vssd1 vccd1 vccd1 _00939_ sky130_fd_sc_hd__a32o_1
XANTENNA__11384__A1 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07588__B1 net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12152_ net195 net2356 net387 vssd1 vssd1 vccd1 vccd1 _00873_ sky130_fd_sc_hd__mux2_1
XANTENNA__10773__A_N net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08033__A net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11103_ final_design.CPU_instr_adr\[31\] _03804_ net1059 vssd1 vssd1 vccd1 vccd1
+ _05824_ sky130_fd_sc_hd__mux2_1
XANTENNA__09329__A1 net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12083_ net579 _06018_ net511 net394 net2190 vssd1 vssd1 vccd1 vccd1 _00808_ sky130_fd_sc_hd__a32o_1
XANTENNA__12333__B1 net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11034_ _04421_ net252 vssd1 vssd1 vccd1 vccd1 _05758_ sky130_fd_sc_hd__nor2_1
XANTENNA__07872__A net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12985_ net1316 _00216_ net1165 vssd1 vssd1 vccd1 vccd1 final_design.CPU_instr_adr\[5\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_19_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11936_ _06137_ net278 net408 net2498 vssd1 vssd1 vccd1 vccd1 _00671_ sky130_fd_sc_hd__a22o_1
XFILLER_0_73_1566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_1905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07811__S net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11867_ _06108_ net287 net518 net2451 vssd1 vssd1 vccd1 vccd1 _00613_ sky130_fd_sc_hd__a22o_1
X_13606_ clknet_leaf_50_clk _00837_ net1172 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[594\]
+ sky130_fd_sc_hd__dfrtp_1
X_10818_ _05530_ _05533_ _05550_ vssd1 vssd1 vccd1 vccd1 _05552_ sky130_fd_sc_hd__or3b_1
X_11798_ net2521 net415 net289 _06018_ vssd1 vssd1 vccd1 vccd1 _00552_ sky130_fd_sc_hd__a22o_1
XFILLER_0_54_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13537_ clknet_leaf_47_clk _00768_ net1203 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[525\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10749_ net74 net1043 vssd1 vssd1 vccd1 vccd1 _05486_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_77_2824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_2201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_2835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07910__S1 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_2846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13468_ clknet_leaf_5_clk _00699_ net1077 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[456\]
+ sky130_fd_sc_hd__dfrtp_1
X_12419_ _06017_ net640 net354 _06280_ vssd1 vssd1 vccd1 vccd1 _01128_ sky130_fd_sc_hd__a31o_1
XANTENNA__12164__S net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11375__A1 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13399_ clknet_leaf_6_clk _00630_ net1130 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[387\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14004__RESET_B net1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07960_ net714 _02910_ vssd1 vssd1 vccd1 vccd1 _02911_ sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_4_clk clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_4_clk sky130_fd_sc_hd__clkbuf_8
X_06911_ net756 _01861_ vssd1 vssd1 vccd1 vccd1 _01862_ sky130_fd_sc_hd__nor2_1
X_07891_ final_design.cpu.reg_window\[471\] final_design.cpu.reg_window\[503\] net849
+ vssd1 vssd1 vccd1 vccd1 _02842_ sky130_fd_sc_hd__mux2_1
XANTENNA__11678__A2 net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11508__S net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09630_ _02868_ _04547_ _04548_ net449 vssd1 vssd1 vccd1 vccd1 _04549_ sky130_fd_sc_hd__a211o_1
X_06842_ final_design.cpu.reg_window\[468\] final_design.cpu.reg_window\[500\] net948
+ vssd1 vssd1 vccd1 vccd1 _01793_ sky130_fd_sc_hd__mux2_1
X_09561_ net73 _04185_ net74 vssd1 vssd1 vccd1 vccd1 _04480_ sky130_fd_sc_hd__o21ai_1
XANTENNA__13742__CLK clknet_leaf_43_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06773_ _01723_ vssd1 vssd1 vccd1 vccd1 _01724_ sky130_fd_sc_hd__inv_2
XANTENNA__12627__B2 final_design.data_from_mem\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08512_ final_design.cpu.reg_window\[66\] final_design.cpu.reg_window\[98\] net837
+ vssd1 vssd1 vccd1 vccd1 _03463_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09492_ net552 _01717_ net551 net550 net458 net468 vssd1 vssd1 vccd1 vccd1 _04411_
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_37_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08443_ final_design.cpu.reg_window\[452\] final_design.cpu.reg_window\[484\] net821
+ vssd1 vssd1 vccd1 vccd1 _03394_ sky130_fd_sc_hd__mux2_1
XANTENNA__11850__A2 net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout249_A _04986_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13892__CLK clknet_leaf_52_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08059__A1 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08374_ net610 _03321_ _03323_ _02211_ vssd1 vssd1 vccd1 vccd1 _03325_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_4_1459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07325_ final_design.cpu.reg_window\[68\] final_design.cpu.reg_window\[100\] net902
+ vssd1 vssd1 vccd1 vccd1 _02276_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_22_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11063__B1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_22_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1060_A final_design.reqhand.current_client\[3\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_2_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout416_A net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07256_ final_design.cpu.reg_window\[583\] final_design.cpu.reg_window\[615\] net887
+ vssd1 vssd1 vccd1 vccd1 _02207_ sky130_fd_sc_hd__mux2_1
XANTENNA__09008__B1 net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13122__CLK clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07187_ final_design.cpu.reg_window\[73\] final_design.cpu.reg_window\[105\] net888
+ vssd1 vssd1 vccd1 vccd1 _02138_ sky130_fd_sc_hd__mux2_1
XANTENNA__11366__A1 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07665__S0 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout785_A net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13272__CLK clknet_leaf_63_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout410 net411 vssd1 vssd1 vccd1 vccd1 net410 sky130_fd_sc_hd__clkbuf_8
Xfanout421 net422 vssd1 vssd1 vccd1 vccd1 net421 sky130_fd_sc_hd__buf_4
Xfanout432 _05847_ vssd1 vssd1 vccd1 vccd1 net432 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_6_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07692__A _01599_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11926__B net240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout443 net444 vssd1 vssd1 vccd1 vccd1 net443 sky130_fd_sc_hd__clkbuf_4
Xfanout454 net455 vssd1 vssd1 vccd1 vccd1 net454 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout573_X net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout952_A net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11418__S net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout465 net466 vssd1 vssd1 vccd1 vccd1 net465 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_35_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08534__A2 _03481_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout476 _03484_ vssd1 vssd1 vccd1 vccd1 net476 sky130_fd_sc_hd__clkbuf_4
X_09828_ _04182_ _04746_ vssd1 vssd1 vccd1 vccd1 _04747_ sky130_fd_sc_hd__nand2_1
Xfanout487 net488 vssd1 vssd1 vccd1 vccd1 net487 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout498 net501 vssd1 vssd1 vccd1 vccd1 net498 sky130_fd_sc_hd__buf_4
XFILLER_0_57_1517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09759_ _04659_ _04677_ vssd1 vssd1 vccd1 vccd1 _04678_ sky130_fd_sc_hd__or2_1
XANTENNA__12618__A1 final_design.reqhand.data_from_UART\[4\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_69_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_1241 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12770_ net1043 _06333_ vssd1 vssd1 vccd1 vccd1 _01357_ sky130_fd_sc_hd__and2_1
XFILLER_0_74_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09495__B1 net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11721_ net188 net628 vssd1 vssd1 vccd1 vccd1 _06219_ sky130_fd_sc_hd__and2_1
XANTENNA__11661__B net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11652_ net433 net574 _06183_ net301 net1501 vssd1 vssd1 vccd1 vccd1 _00458_ sky130_fd_sc_hd__a32o_1
XFILLER_0_65_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10603_ _05329_ _05345_ _05344_ vssd1 vssd1 vccd1 vccd1 _05347_ sky130_fd_sc_hd__o21bai_4
XFILLER_0_65_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11583_ net430 net569 _06147_ net303 net1686 vssd1 vssd1 vccd1 vccd1 _00425_ sky130_fd_sc_hd__a32o_1
XFILLER_0_25_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input81_A memory_size[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13322_ clknet_leaf_59_clk _00553_ net1143 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[310\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10534_ net668 _05269_ _05281_ vssd1 vssd1 vccd1 vccd1 _05282_ sky130_fd_sc_hd__o21a_1
XFILLER_0_10_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11389__A net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10465_ final_design.CPU_instr_adr\[0\] net68 net1054 vssd1 vssd1 vccd1 vccd1 _05217_
+ sky130_fd_sc_hd__mux2_1
X_13253_ clknet_leaf_49_clk _00484_ net1184 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[241\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11357__A1 net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13615__CLK clknet_leaf_44_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10724__C net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12554__B1 net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12204_ _06132_ net498 net376 net2225 vssd1 vssd1 vccd1 vccd1 _00922_ sky130_fd_sc_hd__a22o_1
XFILLER_0_62_1223 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13184_ clknet_leaf_12_clk _00415_ net1086 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[172\]
+ sky130_fd_sc_hd__dfrtp_1
X_10396_ _01481_ net725 net668 _05174_ vssd1 vssd1 vccd1 vccd1 _05180_ sky130_fd_sc_hd__or4_1
X_12135_ net225 net2384 net387 vssd1 vssd1 vccd1 vccd1 _00856_ sky130_fd_sc_hd__mux2_1
XANTENNA__09970__B2 _04066_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13765__CLK clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12066_ net563 _05891_ net504 net392 net1658 vssd1 vssd1 vccd1 vccd1 _00791_ sky130_fd_sc_hd__a32o_1
XANTENNA__09722__A1 net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09183__C1 _01567_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11017_ _05740_ _05741_ vssd1 vssd1 vccd1 vccd1 _05742_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07959__S1 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12609__B2 final_design.data_from_mem\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12968_ clknet_leaf_13_clk _00206_ net1088 vssd1 vssd1 vccd1 vccd1 final_design.uart.bits_received\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_0_clk_A clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11293__B1 net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11919_ net178 _06248_ _06251_ net274 net2386 vssd1 vssd1 vccd1 vccd1 _00657_ sky130_fd_sc_hd__a32o_1
XANTENNA__12159__S net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12899_ clknet_leaf_62_clk _00137_ net1123 vssd1 vssd1 vccd1 vccd1 net171 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_16_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_16_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13145__CLK clknet_leaf_57_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1779 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_2908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_2919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07110_ final_design.reqhand.instruction\[12\] net973 _02060_ vssd1 vssd1 vccd1 vccd1
+ _02061_ sky130_fd_sc_hd__o21ai_4
X_08090_ _02064_ net599 vssd1 vssd1 vccd1 vccd1 _03041_ sky130_fd_sc_hd__nand2_1
XFILLER_0_82_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06681__A _01627_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06698__S1 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload20 clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 clkload20/Y sky130_fd_sc_hd__bufinv_16
X_07041_ final_design.cpu.reg_window\[654\] final_design.cpu.reg_window\[686\] net897
+ vssd1 vssd1 vccd1 vccd1 _01992_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkload31 clknet_leaf_55_clk vssd1 vssd1 vccd1 vccd1 clkload31/Y sky130_fd_sc_hd__inv_16
XFILLER_0_63_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13295__CLK clknet_leaf_41_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload42 clknet_leaf_34_clk vssd1 vssd1 vccd1 vccd1 clkload42/Y sky130_fd_sc_hd__inv_6
XANTENNA__12545__B1 net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_1487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09961__A1 _04871_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08992_ _03927_ vssd1 vssd1 vccd1 vccd1 _03928_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_wire541_X net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07943_ net876 _02875_ _02881_ _02887_ _02893_ vssd1 vssd1 vccd1 vccd1 _02894_ sky130_fd_sc_hd__o32a_4
XFILLER_0_76_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07874_ final_design.cpu.reg_window\[660\] final_design.cpu.reg_window\[692\] net867
+ vssd1 vssd1 vccd1 vccd1 _02825_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_1837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09613_ _04510_ _04511_ _04531_ vssd1 vssd1 vccd1 vccd1 _04532_ sky130_fd_sc_hd__a21oi_1
X_06825_ _01772_ _01773_ _01774_ _01775_ net778 net792 vssd1 vssd1 vccd1 vccd1 _01776_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_74_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout366_A net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_3050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09544_ _02933_ _04094_ vssd1 vssd1 vccd1 vccd1 _04463_ sky130_fd_sc_hd__nand2_1
X_06756_ final_design.cpu.reg_window\[983\] final_design.cpu.reg_window\[1015\] net929
+ vssd1 vssd1 vccd1 vccd1 _01707_ sky130_fd_sc_hd__mux2_1
XANTENNA__12076__A2 net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06687_ final_design.cpu.reg_window\[89\] final_design.cpu.reg_window\[121\] net935
+ vssd1 vssd1 vccd1 vccd1 _01638_ sky130_fd_sc_hd__mux2_1
X_09475_ net534 net533 net532 net530 net457 net466 vssd1 vssd1 vccd1 vccd1 _04394_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_17_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout533_A _02211_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09492__A3 net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08426_ _03373_ _03374_ _03375_ _03376_ net680 net700 vssd1 vssd1 vccd1 vccd1 _03377_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_47_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14070__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08357_ net716 _03307_ vssd1 vssd1 vccd1 vccd1 _03308_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_24_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout700_A net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout321_X net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11587__A1 net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13638__CLK clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout419_X net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload3 clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 clkload3/Y sky130_fd_sc_hd__clkinv_8
XTAP_TAPCELL_ROW_43_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07308_ _02255_ _02256_ _02257_ _02258_ net770 net789 vssd1 vssd1 vccd1 vccd1 _02259_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_33_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08452__A1 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08288_ final_design.cpu.reg_window\[73\] final_design.cpu.reg_window\[105\] net807
+ vssd1 vssd1 vccd1 vccd1 _03239_ sky130_fd_sc_hd__mux2_1
XANTENNA__10384__Y _05173_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07239_ final_design.cpu.reg_window\[71\] final_design.cpu.reg_window\[103\] net887
+ vssd1 vssd1 vccd1 vccd1 _02190_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12536__B1 net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10250_ final_design.uart.BAUD_counter\[18\] _05118_ net798 vssd1 vssd1 vccd1 vccd1
+ _05120_ sky130_fd_sc_hd__o21ai_1
XANTENNA__12000__A2 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13788__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout690_X net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout788_X net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09952__A1 net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10181_ _05067_ _05068_ _05070_ vssd1 vssd1 vccd1 vccd1 _05071_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_37_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06766__A1 net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1205 net1207 vssd1 vssd1 vccd1 vccd1 net1205 sky130_fd_sc_hd__clkbuf_4
Xfanout1216 net1217 vssd1 vssd1 vccd1 vccd1 net1216 sky130_fd_sc_hd__buf_2
Xfanout1227 net1245 vssd1 vssd1 vccd1 vccd1 net1227 sky130_fd_sc_hd__buf_2
XANTENNA_fanout955_X net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout240 _05890_ vssd1 vssd1 vccd1 vccd1 net240 sky130_fd_sc_hd__buf_2
Xfanout1238 net1244 vssd1 vssd1 vccd1 vccd1 net1238 sky130_fd_sc_hd__clkbuf_4
Xfanout251 _04961_ vssd1 vssd1 vccd1 vccd1 net251 sky130_fd_sc_hd__buf_4
XANTENNA__13018__CLK clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09704__A1 _04116_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout262 net263 vssd1 vssd1 vccd1 vccd1 net262 sky130_fd_sc_hd__buf_1
Xfanout273 net275 vssd1 vssd1 vccd1 vccd1 net273 sky130_fd_sc_hd__buf_4
XANTENNA__09704__B2 net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13940_ clknet_leaf_8_clk _01171_ net1152 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[928\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout284 _06228_ vssd1 vssd1 vccd1 vccd1 net284 sky130_fd_sc_hd__clkbuf_4
Xfanout295 _06194_ vssd1 vssd1 vccd1 vccd1 net295 sky130_fd_sc_hd__clkbuf_8
XANTENNA__07810__S0 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13871_ clknet_leaf_42_clk _01102_ net1223 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[859\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06613__S1 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07191__A1 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12822_ net1372 vssd1 vssd1 vccd1 vccd1 _00263_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__13168__CLK clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11275__B1 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12753_ _06351_ _06384_ _06344_ vssd1 vssd1 vccd1 vccd1 _06390_ sky130_fd_sc_hd__o21ai_1
XANTENNA__09483__A3 net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11704_ net432 net572 _06210_ net297 net1801 vssd1 vssd1 vccd1 vccd1 _00483_ sky130_fd_sc_hd__a32o_1
X_12684_ _06329_ net1432 net980 vssd1 vssd1 vccd1 vccd1 _01344_ sky130_fd_sc_hd__mux2_1
XANTENNA__11027__B1 net1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11635_ net206 net630 vssd1 vssd1 vccd1 vccd1 _06175_ sky130_fd_sc_hd__and2_1
XFILLER_0_0_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07877__S0 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11566_ net208 net634 vssd1 vssd1 vccd1 vccd1 _06139_ sky130_fd_sc_hd__and2_1
XFILLER_0_0_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13305_ clknet_leaf_56_clk _00536_ net1146 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[293\]
+ sky130_fd_sc_hd__dfrtp_1
X_10517_ _05249_ _05265_ vssd1 vssd1 vccd1 vccd1 _05266_ sky130_fd_sc_hd__xnor2_1
X_11497_ _02359_ _05838_ vssd1 vssd1 vccd1 vccd1 _06116_ sky130_fd_sc_hd__nor2_4
XANTENNA__12527__B1 net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13236_ clknet_leaf_12_clk _00467_ net1088 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[224\]
+ sky130_fd_sc_hd__dfrtp_1
X_10448_ _02731_ net592 vssd1 vssd1 vccd1 vccd1 _05208_ sky130_fd_sc_hd__nor2_1
XFILLER_0_46_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13167_ clknet_leaf_42_clk _00398_ net1220 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[155\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12442__S net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10379_ net22 net1023 net1007 final_design.data_from_mem\[28\] vssd1 vssd1 vccd1
+ vccd1 _00132_ sky130_fd_sc_hd__o22a_1
XFILLER_0_21_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12118_ net2271 net192 net391 vssd1 vssd1 vccd1 vccd1 _00842_ sky130_fd_sc_hd__mux2_1
XANTENNA__09317__A net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11566__B net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13098_ clknet_leaf_61_clk _00329_ net1140 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[86\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12049_ net1826 net195 net397 vssd1 vssd1 vccd1 vccd1 _00777_ sky130_fd_sc_hd__mux2_1
XANTENNA__11502__A1 net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06610_ final_design.cpu.reg_window\[668\] final_design.cpu.reg_window\[700\] net946
+ vssd1 vssd1 vccd1 vccd1 _01561_ sky130_fd_sc_hd__mux2_1
X_07590_ _02504_ net617 vssd1 vssd1 vccd1 vccd1 _02541_ sky130_fd_sc_hd__nor2_1
XANTENNA__14093__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06541_ _01482_ _01464_ net880 vssd1 vssd1 vccd1 vccd1 _01492_ sky130_fd_sc_hd__and3b_1
XFILLER_0_75_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11805__A2 net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09474__A3 net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09260_ net95 _04178_ vssd1 vssd1 vccd1 vccd1 _04179_ sky130_fd_sc_hd__and2_1
X_06472_ final_design.cpu.reg_window\[350\] final_design.cpu.reg_window\[382\] net933
+ vssd1 vssd1 vccd1 vccd1 _01423_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09202__D _04120_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08211_ net612 _03160_ _03161_ net541 vssd1 vssd1 vccd1 vccd1 _03162_ sky130_fd_sc_hd__a211oi_4
XANTENNA__06693__B1 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09191_ net478 _04083_ vssd1 vssd1 vccd1 vccd1 _04110_ sky130_fd_sc_hd__and2_1
XANTENNA__12617__S _05080_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11521__S net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08142_ final_design.cpu.reg_window\[909\] final_design.cpu.reg_window\[941\] net854
+ vssd1 vssd1 vccd1 vccd1 _03093_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13930__CLK clknet_leaf_60_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08073_ net602 _03022_ _02998_ vssd1 vssd1 vccd1 vccd1 _03024_ sky130_fd_sc_hd__o21ai_1
XANTENNA__12518__B1 net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07024_ _01971_ _01972_ _01973_ _01974_ net768 net788 vssd1 vssd1 vccd1 vccd1 _01975_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_60_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09934__A1 net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07954__B net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1023_A net1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07446__S net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08975_ _03748_ _03911_ vssd1 vssd1 vccd1 vccd1 _03912_ sky130_fd_sc_hd__xnor2_1
Xhold15 net109 vssd1 vssd1 vccd1 vccd1 net1357 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_32_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout483_A net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold26 final_design.cpu.reg_window\[15\] vssd1 vssd1 vccd1 vccd1 net1368 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_32_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold37 net122 vssd1 vssd1 vccd1 vccd1 net1379 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_51_1945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07926_ final_design.cpu.reg_window\[22\] final_design.cpu.reg_window\[54\] net837
+ vssd1 vssd1 vccd1 vccd1 _02877_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_51_1956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold48 final_design.VGA_data_control.data_to_VGA\[31\] vssd1 vssd1 vccd1 vccd1 net1390
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold59 final_design.VGA_data_control.data_to_VGA\[2\] vssd1 vssd1 vccd1 vccd1 net1401
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_51_1967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09698__B1 net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1011 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09162__A2 _03550_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08596__S1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13310__CLK clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout650_A _05849_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07857_ final_design.cpu.reg_window\[468\] final_design.cpu.reg_window\[500\] net868
+ vssd1 vssd1 vccd1 vccd1 _02808_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout271_X net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout748_A _01438_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout369_X net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06808_ _01757_ _01758_ vssd1 vssd1 vccd1 vccd1 _01759_ sky130_fd_sc_hd__nand2_1
X_07788_ _01660_ net604 vssd1 vssd1 vccd1 vccd1 _02739_ sky130_fd_sc_hd__nand2_1
XANTENNA__12954__RESET_B net1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09527_ net472 _04336_ _04223_ vssd1 vssd1 vccd1 vccd1 _04446_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_78_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_1874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06739_ net742 net667 _01504_ _01689_ vssd1 vssd1 vccd1 vccd1 _01690_ sky130_fd_sc_hd__o211a_2
XANTENNA_fanout915_A net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_60_clk_X clknet_leaf_60_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13460__CLK clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09458_ _04308_ net470 _04054_ vssd1 vssd1 vccd1 vccd1 _04377_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_45_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08409_ _02267_ net610 vssd1 vssd1 vccd1 vccd1 _03360_ sky130_fd_sc_hd__or2_1
XFILLER_0_47_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout703_X net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09389_ net465 _03553_ _04061_ vssd1 vssd1 vccd1 vccd1 _04308_ sky130_fd_sc_hd__or3_1
XFILLER_0_30_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11431__S net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_720 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11420_ net1838 net216 net310 vssd1 vssd1 vccd1 vccd1 _00317_ sky130_fd_sc_hd__mux2_1
XANTENNA__07859__S0 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09622__B1 net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11351_ net737 _03853_ _06040_ vssd1 vssd1 vccd1 vccd1 _06041_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_21_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06987__A1 net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10783__A2 net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12509__B1 net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10302_ final_design.VGA_data_control.data_to_VGA\[15\] final_design.VGA_data_control.data_to_VGA\[14\]
+ final_design.VGA_data_control.data_to_VGA\[13\] final_design.VGA_data_control.data_to_VGA\[12\]
+ net1050 net1049 vssd1 vssd1 vccd1 vccd1 _05156_ sky130_fd_sc_hd__mux4_1
XFILLER_0_43_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14070_ clknet_leaf_14_clk _01267_ net1106 vssd1 vssd1 vccd1 vccd1 final_design.uart.working_data\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_11282_ net650 net223 vssd1 vssd1 vccd1 vccd1 _05981_ sky130_fd_sc_hd__and2_1
XANTENNA__12770__B _06333_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13021_ clknet_leaf_2_clk _00252_ net1064 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11667__A net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10233_ final_design.uart.BAUD_counter\[12\] _05108_ vssd1 vssd1 vccd1 vccd1 _05109_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_30_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07087__S1 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11732__A1 net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07356__S net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input44_A mem_adr_start[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10164_ final_design.VGA_data_control.VGA_request_address\[1\] final_design.VGA_data_control.VGA_request_address\[0\]
+ vssd1 vssd1 vccd1 vccd1 _05058_ sky130_fd_sc_hd__and2_2
XANTENNA__09137__A net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1002 net1003 vssd1 vssd1 vccd1 vccd1 net1002 sky130_fd_sc_hd__clkbuf_4
Xfanout1013 net1017 vssd1 vssd1 vccd1 vccd1 net1013 sky130_fd_sc_hd__buf_4
Xfanout1024 _05169_ vssd1 vssd1 vccd1 vccd1 net1024 sky130_fd_sc_hd__clkbuf_4
Xfanout1035 net1036 vssd1 vssd1 vccd1 vccd1 net1035 sky130_fd_sc_hd__clkbuf_4
Xfanout1046 final_design.VGA_adr\[10\] vssd1 vssd1 vccd1 vccd1 net1046 sky130_fd_sc_hd__clkbuf_2
X_10095_ final_design.VGA_data_control.h_count\[5\] _05010_ vssd1 vssd1 vccd1 vccd1
+ _05011_ sky130_fd_sc_hd__or2_1
XFILLER_0_76_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1057 final_design.reqhand.current_client\[3\] vssd1 vssd1 vccd1 vccd1 net1057
+ sky130_fd_sc_hd__clkbuf_4
Xfanout1068 net1069 vssd1 vssd1 vccd1 vccd1 net1068 sky130_fd_sc_hd__clkbuf_4
XANTENNA_clkbuf_leaf_13_clk_X clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1079 net1080 vssd1 vssd1 vccd1 vccd1 net1079 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11496__A0 net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07880__A _01504_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13923_ clknet_leaf_0_clk _01154_ net1071 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[911\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_1745 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_1789 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13803__CLK clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13854_ clknet_leaf_14_clk _01085_ net1103 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[842\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_18_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12805_ net1349 vssd1 vssd1 vccd1 vccd1 _00246_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_clkbuf_leaf_28_clk_X clknet_leaf_28_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13785_ clknet_leaf_55_clk _01016_ net1178 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[773\]
+ sky130_fd_sc_hd__dfrtp_1
X_10997_ _05717_ _05721_ vssd1 vssd1 vccd1 vccd1 _05723_ sky130_fd_sc_hd__and2b_1
XANTENNA__07879__X _02830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12736_ _05059_ _06372_ _06376_ vssd1 vssd1 vccd1 vccd1 _06377_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_61_2274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13953__CLK clknet_leaf_47_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12667_ final_design.VGA_data_control.ready_data\[21\] net1019 net974 final_design.data_from_mem\[21\]
+ vssd1 vssd1 vccd1 vccd1 _06321_ sky130_fd_sc_hd__a22o_1
XANTENNA__12437__S net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_2285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_2296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11618_ net564 net421 _06166_ net299 net1484 vssd1 vssd1 vccd1 vccd1 _00441_ sky130_fd_sc_hd__a32o_1
XFILLER_0_4_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12598_ net1385 net996 net982 final_design.data_from_mem\[16\] vssd1 vssd1 vccd1
+ vccd1 _01291_ sky130_fd_sc_hd__a22o_1
XFILLER_0_13_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08511__S1 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07624__C1 _01535_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11549_ net569 net422 _06130_ net303 net2066 vssd1 vssd1 vccd1 vccd1 _00408_ sky130_fd_sc_hd__a32o_1
Xhold507 final_design.cpu.reg_window\[834\] vssd1 vssd1 vccd1 vccd1 net1849 sky130_fd_sc_hd__dlygate4sd3_1
Xhold518 final_design.cpu.reg_window\[329\] vssd1 vssd1 vccd1 vccd1 net1860 sky130_fd_sc_hd__dlygate4sd3_1
Xhold529 final_design.cpu.reg_window\[1007\] vssd1 vssd1 vccd1 vccd1 net1871 sky130_fd_sc_hd__dlygate4sd3_1
X_12790__21 clknet_leaf_30_clk vssd1 vssd1 vccd1 vccd1 net1331 sky130_fd_sc_hd__inv_2
XFILLER_0_0_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13219_ clknet_leaf_0_clk _00450_ net1062 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[207\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12172__S net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_2078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14199_ net1257 vssd1 vssd1 vccd1 vccd1 gpio_oeb[11] sky130_fd_sc_hd__buf_2
XFILLER_0_21_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_2089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07266__S net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13333__CLK clknet_leaf_56_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06825__S1 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1207 final_design.uart.BAUD_counter\[31\] vssd1 vssd1 vccd1 vccd1 net2549 sky130_fd_sc_hd__dlygate4sd3_1
X_08760_ _03709_ _03710_ vssd1 vssd1 vccd1 vccd1 _03711_ sky130_fd_sc_hd__and2b_1
X_07711_ final_design.cpu.reg_window\[859\] final_design.cpu.reg_window\[891\] net863
+ vssd1 vssd1 vccd1 vccd1 _02662_ sky130_fd_sc_hd__mux2_1
XANTENNA__09144__A2 net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08578__S1 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08691_ _03554_ _03639_ vssd1 vssd1 vccd1 vccd1 _03642_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_69_Left_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11516__S net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13483__CLK clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07642_ final_design.cpu.reg_window\[924\] final_design.cpu.reg_window\[956\] net866
+ vssd1 vssd1 vccd1 vccd1 _02593_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06902__A1 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07573_ final_design.cpu.reg_window\[223\] final_design.cpu.reg_window\[255\] net857
+ vssd1 vssd1 vccd1 vccd1 _02524_ sky130_fd_sc_hd__mux2_1
X_09312_ _04092_ _04218_ vssd1 vssd1 vccd1 vccd1 _04231_ sky130_fd_sc_hd__or2_4
X_06524_ _01454_ _01455_ _01471_ net968 vssd1 vssd1 vccd1 vccd1 _01475_ sky130_fd_sc_hd__a211o_2
X_09243_ _04134_ _04159_ _04161_ _02995_ vssd1 vssd1 vccd1 vccd1 _04162_ sky130_fd_sc_hd__a211o_1
X_06455_ _01405_ _01406_ _01407_ _01396_ vssd1 vssd1 vccd1 vccd1 _01408_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout231_A net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout329_A _06284_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09174_ net527 _04092_ vssd1 vssd1 vccd1 vccd1 _04093_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_78_Left_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07030__A net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08125_ final_design.cpu.reg_window\[269\] final_design.cpu.reg_window\[301\] net850
+ vssd1 vssd1 vccd1 vccd1 _03076_ sky130_fd_sc_hd__mux2_1
XANTENNA__10094__C _05008_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1238_A net1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08056_ final_design.cpu.reg_window\[146\] final_design.cpu.reg_window\[178\] net839
+ vssd1 vssd1 vccd1 vccd1 _03007_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_1600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout698_A net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07007_ final_design.cpu.reg_window\[911\] final_design.cpu.reg_window\[943\] net892
+ vssd1 vssd1 vccd1 vccd1 _01958_ sky130_fd_sc_hd__mux2_1
XFILLER_0_29_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09907__A1 _04072_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08266__S0 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11714__A1 net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07029__X _01980_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout865_A net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13826__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08958_ _01855_ _01856_ vssd1 vssd1 vccd1 vccd1 _03897_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_58_1420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07909_ final_design.cpu.reg_window\[535\] final_design.cpu.reg_window\[567\] net849
+ vssd1 vssd1 vccd1 vccd1 _02860_ sky130_fd_sc_hd__mux2_1
X_08889_ net624 _03833_ _03834_ _03835_ net256 vssd1 vssd1 vccd1 vccd1 _03836_ sky130_fd_sc_hd__a311o_1
XANTENNA__07146__A1 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06587__Y _01538_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11426__S net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10920_ _04550_ net248 net670 vssd1 vssd1 vccd1 vccd1 _05649_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_54_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10150__B1 net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07241__S1 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_1339 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12850__CLK clknet_leaf_19_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10851_ net1004 _05582_ _05583_ net1036 net1361 vssd1 vssd1 vccd1 vccd1 _00192_ sky130_fd_sc_hd__a32o_1
XANTENNA__13976__CLK clknet_leaf_65_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13570_ clknet_leaf_3_clk _00801_ net1067 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[558\]
+ sky130_fd_sc_hd__dfrtp_1
X_10782_ net959 _05516_ _05517_ net956 vssd1 vssd1 vccd1 vccd1 _05518_ sky130_fd_sc_hd__o22a_1
XANTENNA__09843__B1 net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12765__B net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12521_ _06183_ net352 net329 net1834 vssd1 vssd1 vccd1 vccd1 _01226_ sky130_fd_sc_hd__a22o_1
XFILLER_0_26_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11650__B1 net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10453__B2 net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13206__CLK clknet_leaf_60_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_40_clk_A clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1913 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12452_ net2261 net198 net336 vssd1 vssd1 vccd1 vccd1 _01159_ sky130_fd_sc_hd__mux2_1
X_11403_ net657 _06084_ _06086_ vssd1 vssd1 vccd1 vccd1 _06087_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_10_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12383_ net1557 _06003_ net269 vssd1 vssd1 vccd1 vccd1 _01094_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_10_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_1793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10300__S1 net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14122_ clknet_leaf_21_clk final_design.vga.v_next_count\[2\] net1159 vssd1 vssd1
+ vccd1 vccd1 final_design.VGA_data_control.v_count\[2\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_65_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11334_ net663 _03864_ net737 vssd1 vssd1 vccd1 vccd1 _06026_ sky130_fd_sc_hd__a21oi_1
XANTENNA__13356__CLK clknet_leaf_45_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_55_clk_A clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07621__A2 _02570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11397__A net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1891 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14053_ clknet_leaf_16_clk _00014_ net1093 vssd1 vssd1 vccd1 vccd1 final_design.uart.BAUD_counter\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_11265_ net646 net561 net208 vssd1 vssd1 vccd1 vccd1 _05966_ sky130_fd_sc_hd__and3_1
XFILLER_0_82_1793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10508__A2 net1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07086__S net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13004_ net1335 _00235_ net1233 vssd1 vssd1 vccd1 vccd1 final_design.CPU_instr_adr\[24\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_73_2690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10216_ _05098_ net799 _05097_ vssd1 vssd1 vccd1 vccd1 _00033_ sky130_fd_sc_hd__and3b_1
X_11196_ net646 net237 vssd1 vssd1 vccd1 vccd1 _05905_ sky130_fd_sc_hd__and2_1
XANTENNA__11181__A2 net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10147_ final_design.VGA_data_control.h_count\[0\] net1050 vssd1 vssd1 vccd1 vccd1
+ _05047_ sky130_fd_sc_hd__nand2_1
XANTENNA__11469__A0 net209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10078_ wb_manage.curr_state\[2\] wb_manage.curr_state\[1\] vssd1 vssd1 vccd1 vccd1
+ _04995_ sky130_fd_sc_hd__or2_1
X_13906_ clknet_leaf_44_clk _01137_ net1212 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[894\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07688__A2 _02635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_67_2483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07115__A _02058_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10692__A1 net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_2494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13837_ clknet_leaf_53_clk _01068_ net1190 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[825\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10692__B2 _04042_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_2347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_2358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_2369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13768_ clknet_leaf_40_clk _00999_ net1220 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[756\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08637__A1 net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09834__B1 net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09330__A _01493_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06648__B1 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12719_ _06355_ _06358_ _06356_ vssd1 vssd1 vccd1 vccd1 _06360_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12167__S net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_0_clk clk vssd1 vssd1 vccd1 vccd1 clknet_0_clk sky130_fd_sc_hd__clkbuf_16
XANTENNA__10476__A net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13699_ clknet_leaf_0_clk _00930_ net1061 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[687\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14131__CLK clknet_leaf_18_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_731 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13664__RESET_B net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09062__A1 net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold304 final_design.cpu.reg_window\[49\] vssd1 vssd1 vccd1 vccd1 net1646 sky130_fd_sc_hd__dlygate4sd3_1
Xhold315 final_design.cpu.reg_window\[691\] vssd1 vssd1 vccd1 vccd1 net1657 sky130_fd_sc_hd__dlygate4sd3_1
Xhold326 final_design.cpu.reg_window\[532\] vssd1 vssd1 vccd1 vccd1 net1668 sky130_fd_sc_hd__dlygate4sd3_1
Xhold337 final_design.cpu.reg_window\[527\] vssd1 vssd1 vccd1 vccd1 net1679 sky130_fd_sc_hd__dlygate4sd3_1
Xhold348 final_design.cpu.reg_window\[763\] vssd1 vssd1 vccd1 vccd1 net1690 sky130_fd_sc_hd__dlygate4sd3_1
X_09930_ _04178_ _04829_ _04847_ vssd1 vssd1 vccd1 vccd1 _04849_ sky130_fd_sc_hd__o21bai_1
XANTENNA__06820__B1 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold359 final_design.cpu.reg_window\[91\] vssd1 vssd1 vccd1 vccd1 net1701 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_15_Right_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13849__CLK clknet_leaf_55_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout806 net809 vssd1 vssd1 vccd1 vccd1 net806 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_21_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout817 net818 vssd1 vssd1 vccd1 vccd1 net817 sky130_fd_sc_hd__clkbuf_4
X_09861_ net476 _04397_ net489 vssd1 vssd1 vccd1 vccd1 _04780_ sky130_fd_sc_hd__o21a_1
Xfanout828 net829 vssd1 vssd1 vccd1 vccd1 net828 sky130_fd_sc_hd__buf_2
XANTENNA_clkload16_A clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout839 net841 vssd1 vssd1 vccd1 vccd1 net839 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11594__X _06153_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08812_ _03759_ _03762_ vssd1 vssd1 vccd1 vccd1 _03763_ sky130_fd_sc_hd__nand2_1
Xhold1004 final_design.cpu.reg_window\[815\] vssd1 vssd1 vccd1 vccd1 net2346 sky130_fd_sc_hd__dlygate4sd3_1
X_09792_ net540 net539 _02091_ net537 net455 net461 vssd1 vssd1 vccd1 vccd1 _04711_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__10380__B1 net1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1015 final_design.cpu.reg_window\[1021\] vssd1 vssd1 vccd1 vccd1 net2357 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1026 final_design.cpu.reg_window\[627\] vssd1 vssd1 vccd1 vccd1 net2368 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12873__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09505__A _04421_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08743_ _03693_ vssd1 vssd1 vccd1 vccd1 _03694_ sky130_fd_sc_hd__inv_2
Xhold1037 final_design.cpu.reg_window\[275\] vssd1 vssd1 vccd1 vccd1 net2379 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13999__CLK clknet_leaf_43_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1048 final_design.cpu.reg_window\[937\] vssd1 vssd1 vccd1 vccd1 net2390 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1059 final_design.cpu.reg_window\[304\] vssd1 vssd1 vccd1 vccd1 net2401 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07128__A1 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout181_A _06074_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12121__A1 net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout279_A net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09999__X _04918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08674_ _03622_ _03623_ _03624_ _03618_ vssd1 vssd1 vccd1 vccd1 _03625_ sky130_fd_sc_hd__o211a_1
XFILLER_0_75_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07625_ _02573_ _02575_ vssd1 vssd1 vccd1 vccd1 _02576_ sky130_fd_sc_hd__nor2_1
XANTENNA__11880__B1 net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13229__CLK clknet_leaf_48_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_24_Right_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1090_A net1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout446_A _04088_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_631 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1188_A net1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07556_ _01469_ _02094_ vssd1 vssd1 vccd1 vccd1 _02507_ sky130_fd_sc_hd__nand2_4
XANTENNA__12424__A2 net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06507_ _01377_ net1040 net994 net991 vssd1 vssd1 vccd1 vccd1 _01458_ sky130_fd_sc_hd__or4_2
XFILLER_0_9_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11632__B1 net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10435__B2 net246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07487_ _02215_ _02437_ vssd1 vssd1 vccd1 vccd1 _02438_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout613_A net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09226_ _03521_ _03640_ _03520_ vssd1 vssd1 vccd1 vccd1 _04145_ sky130_fd_sc_hd__o21bai_2
XANTENNA__13379__CLK clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09053__A1 net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09157_ net548 net546 net545 net544 net459 net469 vssd1 vssd1 vccd1 vccd1 _04076_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout401_X net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09425__A_N _04342_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1733 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11935__A1 _06136_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09386__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08108_ final_design.cpu.reg_window\[716\] final_design.cpu.reg_window\[748\] net813
+ vssd1 vssd1 vccd1 vccd1 _03059_ sky130_fd_sc_hd__mux2_1
XANTENNA__09239__X _04158_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1777 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09088_ _02300_ _02433_ net619 vssd1 vssd1 vccd1 vccd1 _04012_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout982_A net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_33_Right_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12751__D _05058_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08039_ net717 _02989_ net875 vssd1 vssd1 vccd1 vccd1 _02990_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_31_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08239__S0 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold860 final_design.cpu.reg_window\[867\] vssd1 vssd1 vccd1 vccd1 net2202 sky130_fd_sc_hd__dlygate4sd3_1
Xhold871 final_design.cpu.reg_window\[876\] vssd1 vssd1 vccd1 vccd1 net2213 sky130_fd_sc_hd__dlygate4sd3_1
Xhold882 final_design.cpu.reg_window\[933\] vssd1 vssd1 vccd1 vccd1 net2224 sky130_fd_sc_hd__dlygate4sd3_1
X_11050_ _01387_ _05772_ vssd1 vssd1 vccd1 vccd1 _05774_ sky130_fd_sc_hd__and2_1
Xhold893 final_design.cpu.reg_window\[996\] vssd1 vssd1 vccd1 vccd1 net2235 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout770_X net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_1496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10001_ net83 _04191_ net84 vssd1 vssd1 vccd1 vccd1 _04920_ sky130_fd_sc_hd__o21ai_1
XANTENNA__10371__B1 net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14004__CLK clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1873 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09134__B net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11952_ _06153_ net288 net411 net2074 vssd1 vssd1 vccd1 vccd1 _00687_ sky130_fd_sc_hd__a22o_1
XFILLER_0_73_1737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_42_Right_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10903_ net82 _05610_ _05632_ vssd1 vssd1 vccd1 vccd1 _05633_ sky130_fd_sc_hd__a21o_1
XANTENNA__11871__B1 net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11883_ net672 _06116_ vssd1 vssd1 vccd1 vccd1 _06246_ sky130_fd_sc_hd__nand2_1
XANTENNA__14154__CLK clknet_leaf_18_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13622_ clknet_leaf_62_clk _00853_ net1124 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[610\]
+ sky130_fd_sc_hd__dfrtp_1
X_10834_ net78 net1044 vssd1 vssd1 vccd1 vccd1 _05567_ sky130_fd_sc_hd__and2_1
XFILLER_0_71_1461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12415__A2 net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06774__A _01718_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_2970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_81_2981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10426__B2 net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13553_ clknet_leaf_34_clk _00784_ net1236 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[541\]
+ sky130_fd_sc_hd__dfrtp_1
X_10765_ _05438_ _05457_ _05478_ _05498_ vssd1 vssd1 vccd1 vccd1 _05501_ sky130_fd_sc_hd__nand4_1
XANTENNA__09292__A1 _01657_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12504_ _06166_ net346 net327 net1552 vssd1 vssd1 vccd1 vccd1 _01209_ sky130_fd_sc_hd__a22o_1
X_13484_ clknet_leaf_46_clk _00715_ net1215 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[472\]
+ sky130_fd_sc_hd__dfrtp_1
X_10696_ net39 _05435_ vssd1 vssd1 vccd1 vccd1 _05436_ sky130_fd_sc_hd__and2_1
X_12435_ net1665 net227 net335 vssd1 vssd1 vccd1 vccd1 _01142_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_51_Right_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07809__S net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12366_ net1849 net242 net268 vssd1 vssd1 vccd1 vccd1 _01077_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06713__S net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_75_2752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_75_2763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_2774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14105_ clknet_leaf_24_clk _01302_ net1163 vssd1 vssd1 vccd1 vccd1 final_design.reqhand.instruction\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_71_2616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11317_ net2545 net316 _06011_ net435 vssd1 vssd1 vccd1 vccd1 _00295_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_71_2627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_2638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12297_ net1906 net231 net365 vssd1 vssd1 vccd1 vccd1 _01011_ sky130_fd_sc_hd__mux2_1
X_14036_ clknet_leaf_16_clk _00006_ net1092 vssd1 vssd1 vccd1 vccd1 final_design.uart.BAUD_counter\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12896__CLK clknet_leaf_25_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11248_ net591 _05949_ _05950_ vssd1 vssd1 vccd1 vccd1 _05951_ sky130_fd_sc_hd__and3_2
XANTENNA__12450__S net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10362__B1 net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11179_ _04846_ net651 net588 _05889_ vssd1 vssd1 vccd1 vccd1 _05890_ sky130_fd_sc_hd__o211a_1
XANTENNA__09325__A net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11574__B net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12103__A1 net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_60_Right_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_69_2556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1913 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_2567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_69_2578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11862__B1 net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11590__A net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07410_ net744 net666 net692 _01496_ _02360_ vssd1 vssd1 vccd1 vccd1 _02361_ sky130_fd_sc_hd__o221a_2
XFILLER_0_15_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08390_ final_design.cpu.reg_window\[838\] final_design.cpu.reg_window\[870\] net831
+ vssd1 vssd1 vccd1 vccd1 _03341_ sky130_fd_sc_hd__mux2_1
XANTENNA__12406__A2 net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13845__RESET_B net1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13521__CLK clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07341_ _02288_ _02289_ _02290_ _02291_ net767 net781 vssd1 vssd1 vccd1 vccd1 _02292_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__11614__B1 net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06716__S0 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10968__A2 net1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07272_ final_design.cpu.reg_window\[134\] final_design.cpu.reg_window\[166\] net904
+ vssd1 vssd1 vccd1 vccd1 _02223_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_14_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09011_ _03735_ _03741_ vssd1 vssd1 vccd1 vccd1 _03944_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_14_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13671__CLK clknet_leaf_63_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11378__C1 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold101 final_design.reqhand.instruction\[15\] vssd1 vssd1 vccd1 vccd1 net1443 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_63_1917 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold112 net159 vssd1 vssd1 vccd1 vccd1 net1454 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold123 final_design.VGA_data_control.ready_data\[11\] vssd1 vssd1 vccd1 vccd1 net1465
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11393__A2 net235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold134 final_design.cpu.reg_window\[718\] vssd1 vssd1 vccd1 vccd1 net1476 sky130_fd_sc_hd__dlygate4sd3_1
Xhold145 final_design.VGA_data_control.ready_data\[2\] vssd1 vssd1 vccd1 vccd1 net1487
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12590__B2 final_design.data_from_mem\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold156 final_design.cpu.reg_window\[714\] vssd1 vssd1 vccd1 vccd1 net1498 sky130_fd_sc_hd__dlygate4sd3_1
Xhold167 final_design.VGA_data_control.ready_data\[15\] vssd1 vssd1 vccd1 vccd1 net1509
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold178 final_design.cpu.reg_window\[217\] vssd1 vssd1 vccd1 vccd1 net1520 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09338__A2 net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09913_ _03423_ _04087_ vssd1 vssd1 vccd1 vccd1 _04832_ sky130_fd_sc_hd__nand2_1
XANTENNA__14027__CLK clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold189 final_design.reqhand.instruction\[7\] vssd1 vssd1 vccd1 vccd1 net1531 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout603 net607 vssd1 vssd1 vccd1 vccd1 net603 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout614 net615 vssd1 vssd1 vccd1 vccd1 net614 sky130_fd_sc_hd__buf_2
XFILLER_0_22_1636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout396_A net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout625 _02506_ vssd1 vssd1 vccd1 vccd1 net625 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_0_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout636 net637 vssd1 vssd1 vccd1 vccd1 net636 sky130_fd_sc_hd__buf_4
Xfanout647 net648 vssd1 vssd1 vccd1 vccd1 net647 sky130_fd_sc_hd__buf_2
X_09844_ _04761_ _04762_ _04760_ vssd1 vssd1 vccd1 vccd1 _04763_ sky130_fd_sc_hd__a21oi_1
Xfanout658 _05142_ vssd1 vssd1 vccd1 vccd1 net658 sky130_fd_sc_hd__buf_4
XANTENNA_fanout1103_A net1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10353__B1 _05170_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout669 net670 vssd1 vssd1 vccd1 vccd1 net669 sky130_fd_sc_hd__clkbuf_4
X_09775_ net494 _04693_ vssd1 vssd1 vccd1 vccd1 _04694_ sky130_fd_sc_hd__nand2_1
XFILLER_0_20_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout563_A net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06987_ net886 _01930_ _01936_ _01923_ _01924_ vssd1 vssd1 vccd1 vccd1 _01938_ sky130_fd_sc_hd__a32o_2
XANTENNA__13051__CLK clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14177__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08726_ final_design.CPU_instr_adr\[17\] _01909_ vssd1 vssd1 vccd1 vccd1 _03677_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_55_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11853__B1 net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08657_ net604 _02635_ _02611_ _01453_ vssd1 vssd1 vccd1 vccd1 _03608_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout351_X net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout828_A net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06955__S0 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout449_X net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07608_ final_design.cpu.reg_window\[605\] final_design.cpu.reg_window\[637\] net866
+ vssd1 vssd1 vccd1 vccd1 _02559_ sky130_fd_sc_hd__mux2_1
X_08588_ final_design.cpu.reg_window\[960\] final_design.cpu.reg_window\[992\] net827
+ vssd1 vssd1 vccd1 vccd1 _03539_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11605__A0 net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07539_ final_design.cpu.reg_window\[863\] final_design.cpu.reg_window\[895\] net939
+ vssd1 vssd1 vccd1 vccd1 _02490_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09813__A3 net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10550_ final_design.CPU_instr_adr\[5\] _05277_ vssd1 vssd1 vccd1 vccd1 _05297_ sky130_fd_sc_hd__nand2_1
X_09209_ _02868_ _02900_ vssd1 vssd1 vccd1 vccd1 _04128_ sky130_fd_sc_hd__nor2_1
XANTENNA__09026__A1 net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10481_ _05221_ _05228_ _05230_ net1005 vssd1 vssd1 vccd1 vccd1 _05232_ sky130_fd_sc_hd__a31o_1
XANTENNA__10844__A net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12220_ net575 _06148_ net509 net379 net1823 vssd1 vssd1 vccd1 vccd1 _00938_ sky130_fd_sc_hd__a32o_1
XFILLER_0_27_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11659__B net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07588__A1 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09982__C1 net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12151_ _06017_ net2447 net386 vssd1 vssd1 vccd1 vccd1 _00872_ sky130_fd_sc_hd__mux2_1
X_11102_ final_design.CPU_instr_adr\[31\] _05822_ net1056 vssd1 vssd1 vccd1 vccd1
+ _05823_ sky130_fd_sc_hd__mux2_1
X_12082_ net2419 net394 _06264_ _06011_ vssd1 vssd1 vccd1 vccd1 _00807_ sky130_fd_sc_hd__a22o_1
Xhold690 final_design.cpu.reg_window\[93\] vssd1 vssd1 vccd1 vccd1 net2032 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11675__A net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11033_ _05673_ _05753_ _05754_ _05756_ vssd1 vssd1 vccd1 vccd1 _05757_ sky130_fd_sc_hd__a31oi_4
XANTENNA__09734__C1 net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12984_ net1315 _00215_ net1166 vssd1 vssd1 vccd1 vccd1 final_design.CPU_instr_adr\[4\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__13544__CLK clknet_leaf_41_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11935_ _06136_ net282 net409 net2083 vssd1 vssd1 vccd1 vccd1 _00670_ sky130_fd_sc_hd__a22o_1
XFILLER_0_34_1529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06708__S _01415_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11866_ net2499 net519 _06243_ net433 vssd1 vssd1 vccd1 vccd1 _00612_ sky130_fd_sc_hd__a22o_1
XFILLER_0_71_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13605_ clknet_leaf_49_clk _00836_ net1181 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[593\]
+ sky130_fd_sc_hd__dfrtp_1
X_10817_ _05530_ _05533_ _05550_ vssd1 vssd1 vccd1 vccd1 _05551_ sky130_fd_sc_hd__o21bai_1
X_11797_ net2536 net414 _06235_ net435 vssd1 vssd1 vccd1 vccd1 _00551_ sky130_fd_sc_hd__a22o_1
XANTENNA__13694__CLK clknet_leaf_11_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07276__B1 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13536_ clknet_leaf_11_clk _00767_ net1086 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[524\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10748_ net74 net1043 vssd1 vssd1 vccd1 vccd1 _05485_ sky130_fd_sc_hd__and2_1
XANTENNA__07815__A2 _02763_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_2825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_2202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_2836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13467_ clknet_leaf_65_clk _00698_ net1070 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[455\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12445__S net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10679_ _05419_ vssd1 vssd1 vccd1 vccd1 _05420_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_77_2847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11202__X _05910_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12021__B1 net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12418_ final_design.cpu.reg_window\[885\] net340 vssd1 vssd1 vccd1 vccd1 _06280_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_51_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13398_ clknet_leaf_59_clk _00629_ net1142 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[386\]
+ sky130_fd_sc_hd__dfrtp_1
X_12349_ net2548 net361 net348 _05997_ vssd1 vssd1 vccd1 vccd1 _01061_ sky130_fd_sc_hd__a22o_1
XFILLER_0_23_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10583__B1 net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_1901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13074__CLK clknet_leaf_39_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14019_ clknet_leaf_1_clk _01250_ net1071 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[1007\]
+ sky130_fd_sc_hd__dfrtp_1
X_06910_ _01857_ _01858_ _01859_ _01860_ net773 net791 vssd1 vssd1 vccd1 vccd1 _01861_
+ sky130_fd_sc_hd__mux4_1
X_07890_ final_design.cpu.reg_window\[279\] final_design.cpu.reg_window\[311\] net851
+ vssd1 vssd1 vccd1 vccd1 _02841_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_1445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06841_ final_design.cpu.reg_window\[276\] final_design.cpu.reg_window\[308\] net948
+ vssd1 vssd1 vccd1 vccd1 _01792_ sky130_fd_sc_hd__mux2_1
XANTENNA__10886__B2 net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09560_ _04356_ _04358_ _04390_ _04424_ _04478_ vssd1 vssd1 vccd1 vccd1 _04479_ sky130_fd_sc_hd__o2111a_1
XANTENNA__12088__B1 net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06772_ _01718_ _01722_ vssd1 vssd1 vccd1 vccd1 _01723_ sky130_fd_sc_hd__or2_1
XFILLER_0_78_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08511_ _03458_ _03459_ _03460_ _03461_ net679 net700 vssd1 vssd1 vccd1 vccd1 _03462_
+ sky130_fd_sc_hd__mux4_1
X_09491_ _04408_ _04409_ vssd1 vssd1 vccd1 vccd1 _04410_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_77_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08442_ final_design.cpu.reg_window\[260\] final_design.cpu.reg_window\[292\] net822
+ vssd1 vssd1 vccd1 vccd1 _03393_ sky130_fd_sc_hd__mux2_1
XANTENNA__12911__CLK clknet_leaf_61_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10648__B final_design.VGA_adr\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08373_ net597 _03321_ _03297_ _02211_ vssd1 vssd1 vccd1 vccd1 _03324_ sky130_fd_sc_hd__o211a_1
XFILLER_0_74_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07324_ _02271_ _02272_ _02273_ _02274_ net767 net787 vssd1 vssd1 vccd1 vccd1 _02275_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_45_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_1375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12260__B1 net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1173 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09008__A1 net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07255_ final_design.cpu.reg_window\[647\] final_design.cpu.reg_window\[679\] net890
+ vssd1 vssd1 vccd1 vccd1 _02206_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout311_A _06092_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1053_A net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout409_A net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1861 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12012__B1 net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07186_ final_design.cpu.reg_window\[137\] final_design.cpu.reg_window\[169\] net888
+ vssd1 vssd1 vccd1 vccd1 _02137_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12563__A1 net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13417__CLK clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07665__S1 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_1889 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout680_A net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout400 net401 vssd1 vssd1 vccd1 vccd1 net400 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_6_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout411 _06252_ vssd1 vssd1 vccd1 vccd1 net411 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_6_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout399_X net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout422 _05877_ vssd1 vssd1 vccd1 vccd1 net422 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout778_A net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout433 _05847_ vssd1 vssd1 vccd1 vccd1 net433 sky130_fd_sc_hd__buf_2
XANTENNA__06589__A _01535_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11926__C net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout444 _04090_ vssd1 vssd1 vccd1 vccd1 net444 sky130_fd_sc_hd__buf_2
Xfanout455 _03552_ vssd1 vssd1 vccd1 vccd1 net455 sky130_fd_sc_hd__clkbuf_4
Xfanout466 _03518_ vssd1 vssd1 vccd1 vccd1 net466 sky130_fd_sc_hd__buf_2
X_09827_ net99 _04181_ vssd1 vssd1 vccd1 vccd1 _04746_ sky130_fd_sc_hd__nand2_1
Xfanout477 net480 vssd1 vssd1 vccd1 vccd1 net477 sky130_fd_sc_hd__clkbuf_4
XANTENNA__13567__CLK clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout488 _03454_ vssd1 vssd1 vccd1 vccd1 net488 sky130_fd_sc_hd__buf_2
XANTENNA_fanout945_A net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout566_X net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout499 net501 vssd1 vssd1 vccd1 vccd1 net499 sky130_fd_sc_hd__buf_2
XANTENNA__12079__B1 net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09758_ net450 _04675_ _04672_ net726 vssd1 vssd1 vccd1 vccd1 _04677_ sky130_fd_sc_hd__a211o_1
XFILLER_0_74_1821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08709_ _01359_ _01599_ vssd1 vssd1 vccd1 vccd1 _03660_ sky130_fd_sc_hd__nor2_1
XANTENNA__11826__A0 net206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout733_X net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09689_ net484 _04607_ vssd1 vssd1 vccd1 vccd1 _04608_ sky130_fd_sc_hd__nand2_1
XFILLER_0_70_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11434__S net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11720_ net436 net582 _06218_ net296 net1748 vssd1 vssd1 vccd1 vccd1 _00491_ sky130_fd_sc_hd__a32o_1
XFILLER_0_7_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11651_ net192 net633 vssd1 vssd1 vccd1 vccd1 _06183_ sky130_fd_sc_hd__and2_1
XFILLER_0_65_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10602_ net1416 net1030 net1002 _05346_ vssd1 vssd1 vccd1 vccd1 _00180_ sky130_fd_sc_hd__a22o_1
X_11582_ net194 _06123_ vssd1 vssd1 vccd1 vccd1 _06147_ sky130_fd_sc_hd__and2_1
XANTENNA__12251__B1 net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13321_ clknet_leaf_37_clk _00552_ net1229 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[309\]
+ sky130_fd_sc_hd__dfrtp_1
X_10533_ net801 _05276_ _05280_ net961 vssd1 vssd1 vccd1 vccd1 _05281_ sky130_fd_sc_hd__o22a_1
XFILLER_0_49_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_1871 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1901 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13252_ clknet_leaf_54_clk _00483_ net1179 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[240\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12003__B1 net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input74_A memory_size[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10464_ _04940_ net250 vssd1 vssd1 vccd1 vccd1 _05216_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_23_Left_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07105__S0 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12203_ net564 _06131_ net505 net377 net1618 vssd1 vssd1 vccd1 vccd1 _00921_ sky130_fd_sc_hd__a32o_1
XFILLER_0_0_907 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11357__A2 net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13097__CLK clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13183_ clknet_leaf_7_clk _00414_ net1145 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[171\]
+ sky130_fd_sc_hd__dfrtp_1
X_10395_ net801 net1002 _05179_ net1029 net169 vssd1 vssd1 vccd1 vccd1 _00140_ sky130_fd_sc_hd__a32o_1
XFILLER_0_62_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12134_ net240 net2448 net384 vssd1 vssd1 vccd1 vccd1 _00855_ sky130_fd_sc_hd__mux2_1
XANTENNA__09970__A2 net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12306__A1 net219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07981__A1 net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09707__C1 net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12065_ net2276 net392 net499 _05884_ vssd1 vssd1 vccd1 vccd1 _00790_ sky130_fd_sc_hd__a22o_1
XFILLER_0_19_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09183__B1 _03523_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11016_ _05720_ _05722_ vssd1 vssd1 vccd1 vccd1 _05741_ sky130_fd_sc_hd__nor2_1
XANTENNA__09722__A2 net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12934__CLK clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12609__A2 net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_32_Left_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09486__A1 _01566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12967_ clknet_leaf_12_clk _00205_ net1088 vssd1 vssd1 vccd1 vccd1 final_design.uart.bits_received\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11293__A1 net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11918_ final_design.cpu.reg_window\[414\] _05845_ vssd1 vssd1 vccd1 vccd1 _06251_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_34_1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12490__B1 net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12898_ clknet_leaf_29_clk _00136_ net1195 vssd1 vssd1 vccd1 vccd1 net133 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_75_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_16_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11849_ _06099_ net280 net517 net2275 vssd1 vssd1 vccd1 vccd1 _00599_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_16_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13090__RESET_B net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_2909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12242__B1 net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09789__A2 _04343_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_1471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13519_ clknet_leaf_42_clk _00750_ net1222 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[507\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12175__S net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_41_Left_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06681__B _01630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload10 clknet_leaf_57_clk vssd1 vssd1 vccd1 vccd1 clkload10/Y sky130_fd_sc_hd__inv_8
Xclkload21 clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 clkload21/Y sky130_fd_sc_hd__inv_8
X_07040_ final_design.cpu.reg_window\[718\] final_design.cpu.reg_window\[750\] net897
+ vssd1 vssd1 vccd1 vccd1 _01991_ sky130_fd_sc_hd__mux2_1
Xclkload32 clknet_leaf_41_clk vssd1 vssd1 vccd1 vccd1 clkload32/Y sky130_fd_sc_hd__inv_6
XFILLER_0_67_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload43 clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 clkload43/Y sky130_fd_sc_hd__inv_6
XFILLER_0_2_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09484__S net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08991_ _03792_ _03926_ vssd1 vssd1 vccd1 vccd1 _03927_ sky130_fd_sc_hd__or2_1
XFILLER_0_45_1499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_1791 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07942_ net718 _02892_ net876 vssd1 vssd1 vccd1 vccd1 _02893_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_76_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10843__A2_N net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07873_ final_design.cpu.reg_window\[724\] final_design.cpu.reg_window\[756\] net867
+ vssd1 vssd1 vccd1 vccd1 _02824_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_50_Left_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09612_ _04529_ _04530_ vssd1 vssd1 vccd1 vccd1 _04531_ sky130_fd_sc_hd__xnor2_1
X_06824_ final_design.cpu.reg_window\[917\] final_design.cpu.reg_window\[949\] net937
+ vssd1 vssd1 vccd1 vccd1 _01775_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_1849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_30_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08660__A_N _02542_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_3040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09543_ net495 _04461_ _04231_ vssd1 vssd1 vccd1 vccd1 _04462_ sky130_fd_sc_hd__a21oi_1
X_06755_ final_design.cpu.reg_window\[791\] final_design.cpu.reg_window\[823\] net929
+ vssd1 vssd1 vccd1 vccd1 _01706_ sky130_fd_sc_hd__mux2_1
XANTENNA__11808__B1 net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_3051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09477__A1 _02325_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout261_A _04071_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout359_A _06277_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09474_ net539 net538 net537 net535 net457 net466 vssd1 vssd1 vccd1 vccd1 _04393_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_8_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06686_ _01633_ _01634_ _01635_ _01636_ net774 net792 vssd1 vssd1 vccd1 vccd1 _01637_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__12481__B1 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08425_ final_design.cpu.reg_window\[901\] final_design.cpu.reg_window\[933\] net840
+ vssd1 vssd1 vccd1 vccd1 _03376_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout1170_A net1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08356_ _03303_ _03304_ _03305_ _03306_ net674 net696 vssd1 vssd1 vccd1 vccd1 _03307_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_24_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12233__B1 net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06872__A _01504_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload4 clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 clkload4/Y sky130_fd_sc_hd__inv_8
XANTENNA__11587__A2 net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07307_ final_design.cpu.reg_window\[901\] final_design.cpu.reg_window\[933\] net921
+ vssd1 vssd1 vccd1 vccd1 _02258_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_43_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08287_ net707 _03237_ vssd1 vssd1 vccd1 vccd1 _03238_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout314_X net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1056_X net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07238_ final_design.cpu.reg_window\[135\] final_design.cpu.reg_window\[167\] net887
+ vssd1 vssd1 vccd1 vccd1 _02189_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07169_ final_design.cpu.reg_window\[714\] final_design.cpu.reg_window\[746\] net899
+ vssd1 vssd1 vccd1 vccd1 _02120_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10180_ final_design.uart.BAUD_counter\[29\] final_design.uart.BAUD_counter\[28\]
+ final_design.uart.BAUD_counter\[31\] final_design.uart.BAUD_counter\[30\] vssd1
+ vssd1 vccd1 vccd1 _05070_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout683_X net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11429__S net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1206 net1207 vssd1 vssd1 vccd1 vccd1 net1206 sky130_fd_sc_hd__clkbuf_4
X_12773__4 clknet_leaf_26_clk vssd1 vssd1 vccd1 vccd1 net1314 sky130_fd_sc_hd__inv_2
XANTENNA__12957__CLK clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1217 net1227 vssd1 vssd1 vccd1 vccd1 net1217 sky130_fd_sc_hd__clkbuf_2
Xfanout1228 net1235 vssd1 vssd1 vccd1 vccd1 net1228 sky130_fd_sc_hd__clkbuf_4
Xfanout230 net231 vssd1 vssd1 vccd1 vccd1 net230 sky130_fd_sc_hd__clkbuf_2
Xfanout241 net242 vssd1 vssd1 vccd1 vccd1 net241 sky130_fd_sc_hd__buf_2
Xfanout1239 net1244 vssd1 vssd1 vccd1 vccd1 net1239 sky130_fd_sc_hd__clkbuf_2
Xfanout252 net253 vssd1 vssd1 vccd1 vccd1 net252 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07208__A net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout263 _04071_ vssd1 vssd1 vccd1 vccd1 net263 sky130_fd_sc_hd__clkbuf_4
Xfanout274 net275 vssd1 vssd1 vccd1 vccd1 net274 sky130_fd_sc_hd__clkbuf_8
Xfanout285 net286 vssd1 vssd1 vccd1 vccd1 net285 sky130_fd_sc_hd__clkbuf_4
Xfanout296 net297 vssd1 vssd1 vccd1 vccd1 net296 sky130_fd_sc_hd__buf_4
XANTENNA__08912__B1 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13870_ clknet_leaf_45_clk _01101_ net1216 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[858\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07810__S1 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12821_ net1378 vssd1 vssd1 vccd1 vccd1 _00262_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__09423__A _03627_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12067__A3 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12752_ final_design.VGA_adr\[5\] net796 _06383_ _06388_ _06389_ vssd1 vssd1 vccd1
+ vccd1 _01352_ sky130_fd_sc_hd__a221o_1
XANTENNA__11275__A1 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12472__B1 net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10288__B net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11703_ net222 net629 vssd1 vssd1 vccd1 vccd1 _06210_ sky130_fd_sc_hd__and2_1
XFILLER_0_56_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12683_ final_design.VGA_data_control.ready_data\[29\] net1021 net977 final_design.data_from_mem\[29\]
+ vssd1 vssd1 vccd1 vccd1 _06329_ sky130_fd_sc_hd__a22o_1
XANTENNA__11027__A1 net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12224__B1 net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11634_ net425 net559 _06174_ net298 net2187 vssd1 vssd1 vccd1 vccd1 _00449_ sky130_fd_sc_hd__a32o_1
XFILLER_0_21_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11565_ net434 net577 _06138_ net304 net2488 vssd1 vssd1 vccd1 vccd1 _00416_ sky130_fd_sc_hd__a32o_1
XANTENNA__07877__S1 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06454__A1 net1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13304_ clknet_leaf_63_clk _00535_ net1119 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[292\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10516_ _05263_ _05264_ vssd1 vssd1 vccd1 vccd1 _05265_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_0_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11496_ net176 net2370 net308 vssd1 vssd1 vccd1 vccd1 _00370_ sky130_fd_sc_hd__mux2_1
XANTENNA__13732__CLK clknet_leaf_54_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13235_ clknet_leaf_39_clk _00466_ net1207 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[223\]
+ sky130_fd_sc_hd__dfrtp_1
X_10447_ net149 net1036 _05207_ net249 vssd1 vssd1 vccd1 vccd1 _00164_ sky130_fd_sc_hd__a22o_1
XANTENNA__06721__S net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13166_ clknet_leaf_45_clk _00397_ net1213 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[154\]
+ sky130_fd_sc_hd__dfrtp_1
X_10378_ net21 net1024 net1006 final_design.data_from_mem\[27\] vssd1 vssd1 vccd1
+ vccd1 _00131_ sky130_fd_sc_hd__o22a_1
XFILLER_0_20_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12117_ net1773 net195 net391 vssd1 vssd1 vccd1 vccd1 _00841_ sky130_fd_sc_hd__mux2_1
X_13097_ clknet_leaf_35_clk _00328_ net1236 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[85\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13882__CLK clknet_leaf_58_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12048_ net2469 net196 net398 vssd1 vssd1 vccd1 vccd1 _00776_ sky130_fd_sc_hd__mux2_1
XANTENNA__13112__CLK clknet_leaf_62_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11582__B _06123_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13999_ clknet_leaf_43_clk _01230_ net1222 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[987\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_1713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06540_ _01464_ _01475_ _01483_ vssd1 vssd1 vccd1 vccd1 _01491_ sky130_fd_sc_hd__or3_4
XFILLER_0_1_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11266__B2 net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_1877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06471_ final_design.data_from_mem\[16\] net971 _01421_ vssd1 vssd1 vccd1 vccd1 _01422_
+ sky130_fd_sc_hd__a21oi_4
XANTENNA__13262__CLK clknet_leaf_45_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08210_ _02000_ net611 vssd1 vssd1 vccd1 vccd1 _03161_ sky130_fd_sc_hd__nor2_1
XANTENNA__06693__A1 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07788__A _01660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11018__B2 net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12215__B1 net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08383__S net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09190_ net495 _04107_ vssd1 vssd1 vccd1 vccd1 _04109_ sky130_fd_sc_hd__nand2_4
XANTENNA__06692__A net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11569__A2 net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08141_ final_design.cpu.reg_window\[973\] final_design.cpu.reg_window\[1005\] net854
+ vssd1 vssd1 vccd1 vccd1 _03092_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08072_ _01881_ net618 vssd1 vssd1 vccd1 vccd1 _03023_ sky130_fd_sc_hd__nor2_1
XFILLER_0_15_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07023_ final_design.cpu.reg_window\[398\] final_design.cpu.reg_window\[430\] net898
+ vssd1 vssd1 vccd1 vccd1 _01974_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07727__S net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09395__B1 net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08974_ _03676_ _03677_ vssd1 vssd1 vccd1 vccd1 _03911_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout1016_A net1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold16 net113 vssd1 vssd1 vccd1 vccd1 net1358 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_32_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07925_ final_design.cpu.reg_window\[86\] final_design.cpu.reg_window\[118\] net837
+ vssd1 vssd1 vccd1 vccd1 _02876_ sky130_fd_sc_hd__mux2_1
Xhold27 final_design.cpu.reg_window\[16\] vssd1 vssd1 vccd1 vccd1 net1369 sky130_fd_sc_hd__dlygate4sd3_1
Xhold38 final_design.cpu.reg_window\[6\] vssd1 vssd1 vccd1 vccd1 net1380 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_51_1946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold49 final_design.VGA_data_control.data_to_VGA\[28\] vssd1 vssd1 vccd1 vccd1 net1391
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_51_1957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout476_A _03484_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07856_ final_design.cpu.reg_window\[276\] final_design.cpu.reg_window\[308\] net868
+ vssd1 vssd1 vccd1 vccd1 _02807_ sky130_fd_sc_hd__mux2_1
XANTENNA__08370__B2 net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11492__B _06093_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06807_ net551 _01755_ vssd1 vssd1 vccd1 vccd1 _01758_ sky130_fd_sc_hd__nand2_1
X_07787_ _02737_ vssd1 vssd1 vccd1 vccd1 _02738_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout264_X net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout643_A net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13605__CLK clknet_leaf_49_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09526_ _04342_ _04439_ _04441_ _04444_ vssd1 vssd1 vccd1 vccd1 _04445_ sky130_fd_sc_hd__o22a_1
XFILLER_0_52_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06738_ net742 net879 vssd1 vssd1 vccd1 vccd1 _01689_ sky130_fd_sc_hd__nand2_1
XFILLER_0_17_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_49_1875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_1897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09457_ _04304_ _04307_ net475 vssd1 vssd1 vccd1 vccd1 _04376_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_45_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1190 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06669_ final_design.cpu.reg_window\[602\] final_design.cpu.reg_window\[634\] net936
+ vssd1 vssd1 vccd1 vccd1 _01620_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout431_X net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout908_A net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07698__A net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08408_ _03324_ _03325_ _03355_ _03357_ vssd1 vssd1 vccd1 vccd1 _03359_ sky130_fd_sc_hd__o22a_1
XANTENNA__11009__B2 net1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12206__B1 net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09388_ net530 net529 _02325_ net528 net456 net465 vssd1 vssd1 vccd1 vccd1 _04307_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__07308__S0 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13755__CLK clknet_leaf_65_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08339_ net610 _03287_ _03288_ net534 vssd1 vssd1 vccd1 vccd1 _03290_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_62_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07859__S1 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12221__A3 net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11350_ net661 _03847_ net733 vssd1 vssd1 vccd1 vccd1 _06040_ sky130_fd_sc_hd__o21a_1
XFILLER_0_61_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10301_ _01384_ _05154_ vssd1 vssd1 vccd1 vccd1 _05155_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout898_X net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11980__A2 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11281_ net590 _05978_ _05979_ vssd1 vssd1 vccd1 vccd1 _05980_ sky130_fd_sc_hd__and3_1
XANTENNA__10852__A _04954_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13020_ clknet_leaf_3_clk _00251_ net1066 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_10232_ _05108_ net799 _05107_ vssd1 vssd1 vccd1 vccd1 _00008_ sky130_fd_sc_hd__and3b_1
XANTENNA__11667__B net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06739__A2 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11732__A2 net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10163_ final_design.VGA_data_control.VGA_request_address\[0\] _05054_ final_design.VGA_data_control.VGA_request_address\[1\]
+ vssd1 vssd1 vccd1 vccd1 _05057_ sky130_fd_sc_hd__a21o_1
Xfanout1003 _05173_ vssd1 vssd1 vccd1 vccd1 net1003 sky130_fd_sc_hd__clkbuf_8
XANTENNA__09138__A0 net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08041__B net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1014 net1017 vssd1 vssd1 vccd1 vccd1 net1014 sky130_fd_sc_hd__clkbuf_4
Xfanout1025 _05168_ vssd1 vssd1 vccd1 vccd1 net1025 sky130_fd_sc_hd__clkbuf_4
Xfanout1036 _04994_ vssd1 vssd1 vccd1 vccd1 net1036 sky130_fd_sc_hd__clkbuf_8
XANTENNA__13135__CLK clknet_leaf_42_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1047 final_design.VGA_adr\[10\] vssd1 vssd1 vccd1 vccd1 net1047 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_input37_A mem_adr_start[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10094_ final_design.VGA_data_control.h_count\[8\] final_design.VGA_data_control.h_count\[9\]
+ _05008_ vssd1 vssd1 vccd1 vccd1 _05010_ sky130_fd_sc_hd__or3_1
Xfanout1058 final_design.reqhand.current_client\[3\] vssd1 vssd1 vccd1 vccd1 net1058
+ sky130_fd_sc_hd__buf_2
XANTENNA__12288__A3 net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1069 net1118 vssd1 vssd1 vccd1 vccd1 net1069 sky130_fd_sc_hd__buf_2
X_13922_ clknet_leaf_4_clk _01153_ net1083 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[910\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09424__Y _04343_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1123 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_18_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13853_ clknet_leaf_1_clk _01084_ net1081 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[841\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13285__CLK clknet_leaf_48_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12804_ net1356 vssd1 vssd1 vccd1 vccd1 _00245_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_2_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10996_ _05721_ _05717_ vssd1 vssd1 vccd1 vccd1 _05722_ sky130_fd_sc_hd__and2b_1
X_13784_ clknet_leaf_65_clk _01015_ net1073 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[772\]
+ sky130_fd_sc_hd__dfrtp_1
X_12735_ _06374_ _06375_ _06370_ vssd1 vssd1 vccd1 vccd1 _06376_ sky130_fd_sc_hd__a21o_1
XFILLER_0_70_1356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09861__A1 net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08664__A2 _02061_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06675__A1 net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10471__A2 net1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12666_ _06320_ net1602 net978 vssd1 vssd1 vccd1 vccd1 _01335_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_61_2275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_2286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_2297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11617_ net237 net630 vssd1 vssd1 vccd1 vccd1 _06166_ sky130_fd_sc_hd__and2_1
XFILLER_0_68_1230 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12597_ net1443 net996 net982 final_design.data_from_mem\[15\] vssd1 vssd1 vccd1
+ vccd1 _01290_ sky130_fd_sc_hd__a22o_1
XANTENNA__12212__A3 net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11548_ net224 net635 vssd1 vssd1 vccd1 vccd1 _06130_ sky130_fd_sc_hd__and2_1
XFILLER_0_53_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_1116 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11971__A2 net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold508 final_design.cpu.reg_window\[602\] vssd1 vssd1 vccd1 vccd1 net1850 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_34_990 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11858__A net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold519 final_design.cpu.reg_window\[984\] vssd1 vssd1 vccd1 vccd1 net1861 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12453__S net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11479_ net198 net2503 net308 vssd1 vssd1 vccd1 vccd1 _00359_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07547__S net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13218_ clknet_leaf_3_clk _00449_ net1066 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[206\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09328__A net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14198_ net1256 vssd1 vssd1 vccd1 vccd1 gpio_oeb[10] sky130_fd_sc_hd__buf_2
XFILLER_0_0_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_2079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13149_ clknet_leaf_2_clk _00380_ net1064 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[137\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_1870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14060__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1208 final_design.CPU_instr_adr\[5\] vssd1 vssd1 vccd1 vccd1 net2550 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12279__A3 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07710_ net719 _02660_ vssd1 vssd1 vccd1 vccd1 _02661_ sky130_fd_sc_hd__nor2_1
XANTENNA__13628__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08690_ _02419_ net452 vssd1 vssd1 vccd1 vccd1 _03641_ sky130_fd_sc_hd__nand2_1
XANTENNA__08378__S net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07282__S net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07641_ final_design.cpu.reg_window\[988\] final_design.cpu.reg_window\[1020\] net872
+ vssd1 vssd1 vccd1 vccd1 _02592_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_0_216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06902__A2 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1630 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07572_ final_design.cpu.reg_window\[31\] final_design.cpu.reg_window\[63\] net857
+ vssd1 vssd1 vccd1 vccd1 _02523_ sky130_fd_sc_hd__mux2_1
XANTENNA__11239__B2 net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09311_ _04222_ _04229_ _04218_ vssd1 vssd1 vccd1 vccd1 _04230_ sky130_fd_sc_hd__a21o_1
X_06523_ _01466_ _01467_ _01471_ net968 vssd1 vssd1 vccd1 vccd1 _01474_ sky130_fd_sc_hd__or4_4
XANTENNA__13778__CLK clknet_leaf_39_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11532__S net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09242_ _02994_ _03026_ vssd1 vssd1 vccd1 vccd1 _04161_ sky130_fd_sc_hd__nor2_1
X_06454_ net1057 net1039 final_design.reqhand.current_client\[1\] vssd1 vssd1 vccd1
+ vccd1 _01407_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_7_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09173_ _03635_ net659 vssd1 vssd1 vccd1 vccd1 _04092_ sky130_fd_sc_hd__or2_2
XANTENNA__12203__A3 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout224_A _05897_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_1926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08124_ final_design.cpu.reg_window\[333\] final_design.cpu.reg_window\[365\] net854
+ vssd1 vssd1 vccd1 vccd1 _03075_ sky130_fd_sc_hd__mux2_1
XANTENNA__11411__A1 net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07030__B _01980_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11962__A2 net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08055_ final_design.cpu.reg_window\[210\] final_design.cpu.reg_window\[242\] net844
+ vssd1 vssd1 vccd1 vccd1 _03006_ sky130_fd_sc_hd__mux2_1
XFILLER_0_29_1770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07006_ final_design.cpu.reg_window\[975\] final_design.cpu.reg_window\[1007\] net892
+ vssd1 vssd1 vccd1 vccd1 _01957_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_38_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07457__S net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13158__CLK clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08266__S1 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout593_A _05199_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11714__A2 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09383__A3 net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08957_ _03751_ _03895_ vssd1 vssd1 vccd1 vccd1 _03896_ sky130_fd_sc_hd__xor2_1
XANTENNA_fanout381_X net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout760_A _01426_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout858_A net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07908_ final_design.cpu.reg_window\[599\] final_design.cpu.reg_window\[631\] net846
+ vssd1 vssd1 vccd1 vccd1 _02859_ sky130_fd_sc_hd__mux2_1
X_08888_ net624 _03832_ vssd1 vssd1 vccd1 vccd1 _03835_ sky130_fd_sc_hd__nor2_1
XANTENNA__13122__RESET_B net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07045__X _01996_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07839_ _02786_ _02787_ _02788_ _02789_ net685 net706 vssd1 vssd1 vccd1 vccd1 _02790_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout646_X net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10850_ _05559_ _05564_ _05581_ vssd1 vssd1 vccd1 vccd1 _05583_ sky130_fd_sc_hd__o21ai_1
XANTENNA__12427__B1 net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07920__S net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09509_ _02936_ _04426_ _04160_ _03029_ vssd1 vssd1 vccd1 vccd1 _04428_ sky130_fd_sc_hd__o211ai_1
X_10781_ final_design.CPU_instr_adr\[16\] _03928_ net1060 vssd1 vssd1 vccd1 vccd1
+ _05517_ sky130_fd_sc_hd__mux2_1
X_12520_ _06182_ net349 net327 net1718 vssd1 vssd1 vccd1 vccd1 _01225_ sky130_fd_sc_hd__a22o_1
XANTENNA__11650__A1 net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10453__A2 net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10566__B final_design.VGA_adr\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12451_ net1876 net199 net334 vssd1 vssd1 vccd1 vccd1 _01158_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_1761 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11402_ _01501_ _05946_ _06085_ net645 vssd1 vssd1 vccd1 vccd1 _06086_ sky130_fd_sc_hd__a22o_2
X_12382_ net1942 net202 net270 vssd1 vssd1 vccd1 vccd1 _01093_ sky130_fd_sc_hd__mux2_1
XANTENNA__11402__B2 net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09071__A2 net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14121_ clknet_leaf_21_clk final_design.vga.v_next_count\[1\] net1159 vssd1 vssd1
+ vccd1 vccd1 final_design.VGA_data_control.v_count\[1\] sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_10_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11333_ net2334 net315 _06025_ net430 vssd1 vssd1 vccd1 vccd1 _00297_ sky130_fd_sc_hd__a22o_1
XANTENNA__11953__A2 net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14052_ clknet_leaf_16_clk _00013_ net1093 vssd1 vssd1 vccd1 vccd1 final_design.uart.BAUD_counter\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14083__CLK clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11264_ _04613_ net652 net588 _05964_ vssd1 vssd1 vccd1 vccd1 _05965_ sky130_fd_sc_hd__o211a_2
X_13003_ net1334 _00234_ net1233 vssd1 vssd1 vccd1 vccd1 final_design.CPU_instr_adr\[23\]
+ sky130_fd_sc_hd__dfrtp_2
X_10215_ final_design.uart.BAUD_counter\[5\] final_design.uart.BAUD_counter\[4\] _05094_
+ vssd1 vssd1 vccd1 vccd1 _05098_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_73_2691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11195_ _04723_ net651 net588 _05903_ vssd1 vssd1 vccd1 vccd1 _05904_ sky130_fd_sc_hd__o211a_1
XFILLER_0_78_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10146_ final_design.VGA_data_control.h_count\[0\] _05046_ vssd1 vssd1 vccd1 vccd1
+ final_design.vga.h_next_count\[0\] sky130_fd_sc_hd__and2b_1
XFILLER_0_59_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09154__Y _04073_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10077_ wb_manage.curr_state\[2\] wb_manage.curr_state\[1\] vssd1 vssd1 vccd1 vccd1
+ _04994_ sky130_fd_sc_hd__nor2_1
XANTENNA__08198__S net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_1554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13905_ clknet_leaf_35_clk _01136_ net1243 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[893\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13920__CLK clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkload2_A clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_2484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13836_ clknet_leaf_46_clk _01067_ net1217 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[824\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_67_2495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_2348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_2359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10979_ net959 _05703_ _05705_ net956 vssd1 vssd1 vccd1 vccd1 _05706_ sky130_fd_sc_hd__o22a_1
X_13767_ clknet_leaf_62_clk _00998_ net1123 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[755\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12448__S net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08637__A2 _02961_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06648__A1 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12718_ _06355_ _06356_ _06358_ vssd1 vssd1 vccd1 vccd1 _06359_ sky130_fd_sc_hd__a21o_2
X_13698_ clknet_leaf_11_clk _00929_ net1097 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[686\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_13_1571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12649_ final_design.VGA_data_control.ready_data\[12\] net1020 net975 final_design.data_from_mem\[12\]
+ vssd1 vssd1 vccd1 vccd1 _06312_ sky130_fd_sc_hd__a22o_1
XFILLER_0_26_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13300__CLK clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11944__A2 net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold305 final_design.cpu.reg_window\[243\] vssd1 vssd1 vccd1 vccd1 net1647 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12183__S net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10492__A net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold316 final_design.cpu.reg_window\[548\] vssd1 vssd1 vccd1 vccd1 net1658 sky130_fd_sc_hd__dlygate4sd3_1
Xhold327 final_design.cpu.reg_window\[593\] vssd1 vssd1 vccd1 vccd1 net1669 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_61_1801 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07277__S net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold338 final_design.cpu.reg_window\[590\] vssd1 vssd1 vccd1 vccd1 net1680 sky130_fd_sc_hd__dlygate4sd3_1
Xhold349 final_design.cpu.reg_window\[168\] vssd1 vssd1 vccd1 vccd1 net1691 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06820__A1 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout807 net809 vssd1 vssd1 vccd1 vccd1 net807 sky130_fd_sc_hd__clkbuf_4
X_09860_ _04641_ _04778_ net471 vssd1 vssd1 vccd1 vccd1 _04779_ sky130_fd_sc_hd__mux2_1
XANTENNA__13450__CLK clknet_leaf_60_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout818 net829 vssd1 vssd1 vccd1 vccd1 net818 sky130_fd_sc_hd__clkbuf_2
Xfanout829 _01818_ vssd1 vssd1 vccd1 vccd1 net829 sky130_fd_sc_hd__clkbuf_4
X_08811_ _03760_ _03761_ vssd1 vssd1 vccd1 vccd1 _03762_ sky130_fd_sc_hd__and2_1
X_09791_ net535 net534 net533 net532 net452 net461 vssd1 vssd1 vccd1 vccd1 _04710_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_77_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10380__B2 final_design.data_from_mem\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1005 final_design.cpu.reg_window\[266\] vssd1 vssd1 vccd1 vccd1 net2347 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1016 final_design.cpu.reg_window\[673\] vssd1 vssd1 vccd1 vccd1 net2358 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11527__S net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08742_ net667 _01537_ final_design.CPU_instr_adr\[9\] vssd1 vssd1 vccd1 vccd1 _03693_
+ sky130_fd_sc_hd__a21oi_1
Xhold1027 final_design.cpu.reg_window\[192\] vssd1 vssd1 vccd1 vccd1 net2369 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09505__B _04423_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1038 final_design.cpu.reg_window\[801\] vssd1 vssd1 vccd1 vccd1 net2380 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1049 final_design.cpu.reg_window\[314\] vssd1 vssd1 vccd1 vccd1 net2391 sky130_fd_sc_hd__dlygate4sd3_1
X_08673_ _01999_ _02062_ vssd1 vssd1 vccd1 vccd1 _03624_ sky130_fd_sc_hd__nand2_1
XFILLER_0_16_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07624_ net607 _02570_ _02546_ _01535_ vssd1 vssd1 vccd1 vccd1 _02575_ sky130_fd_sc_hd__o211a_1
XFILLER_0_36_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12409__B1 net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11770__B net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07555_ _01469_ _02094_ vssd1 vssd1 vccd1 vccd1 _02506_ sky130_fd_sc_hd__and2_2
XFILLER_0_76_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1083_A net1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09825__B2 net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout439_A _04095_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06506_ final_design.data_from_mem\[4\] net1041 net993 net990 vssd1 vssd1 vccd1 vccd1
+ _01457_ sky130_fd_sc_hd__and4_1
XANTENNA__11632__A1 net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07486_ _02242_ _02436_ _02241_ vssd1 vssd1 vccd1 vccd1 _02437_ sky130_fd_sc_hd__o21ai_1
XANTENNA__10386__B net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09225_ _03262_ _03293_ vssd1 vssd1 vccd1 vccd1 _04144_ sky130_fd_sc_hd__and2_1
X_06437_ net35 vssd1 vssd1 vccd1 vccd1 _01392_ sky130_fd_sc_hd__inv_2
XFILLER_0_17_732 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout606_A net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout227_X net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09156_ _01717_ net551 net550 _01815_ net458 net468 vssd1 vssd1 vccd1 vccd1 _04075_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_17_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06880__A net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1745 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11935__A2 net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08107_ _03054_ _03055_ _03056_ _03057_ net676 net697 vssd1 vssd1 vccd1 vccd1 _03058_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_20_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09087_ net2550 _04011_ net1037 vssd1 vssd1 vccd1 vccd1 _00216_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_20_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_1144 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08261__B1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1789 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08038_ _02985_ _02986_ _02987_ _02988_ net677 net692 vssd1 vssd1 vccd1 vccd1 _02989_
+ sky130_fd_sc_hd__mux4_1
Xhold850 final_design.cpu.reg_window\[280\] vssd1 vssd1 vccd1 vccd1 net2192 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout975_A _06299_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold861 final_design.cpu.reg_window\[869\] vssd1 vssd1 vccd1 vccd1 net2203 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08239__S1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_27_clk_X clknet_leaf_27_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold872 final_design.cpu.reg_window\[924\] vssd1 vssd1 vccd1 vccd1 net2214 sky130_fd_sc_hd__dlygate4sd3_1
Xhold883 final_design.cpu.reg_window\[679\] vssd1 vssd1 vccd1 vccd1 net2225 sky130_fd_sc_hd__dlygate4sd3_1
Xhold894 final_design.cpu.reg_window\[322\] vssd1 vssd1 vccd1 vccd1 net2236 sky130_fd_sc_hd__dlygate4sd3_1
X_10000_ _04918_ vssd1 vssd1 vccd1 vccd1 _04919_ sky130_fd_sc_hd__inv_2
XANTENNA__12360__A2 net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10371__A1 net14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13943__CLK clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout763_X net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09989_ _04370_ _04773_ _04409_ vssd1 vssd1 vccd1 vccd1 _04908_ sky130_fd_sc_hd__a21bo_1
XANTENNA__10371__B2 final_design.data_from_mem\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11437__S net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_4_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1705 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_1885 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11951_ _06152_ net292 net410 net2195 vssd1 vssd1 vccd1 vccd1 _00686_ sky130_fd_sc_hd__a22o_1
XANTENNA__11320__B1 net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10902_ _05630_ _05631_ _05610_ vssd1 vssd1 vccd1 vccd1 _05632_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_73_1749 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11871__A1 net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11882_ net177 net640 net288 net519 net1946 vssd1 vssd1 vccd1 vccd1 _00626_ sky130_fd_sc_hd__a32o_1
XFILLER_0_58_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10833_ _04571_ net252 _04990_ vssd1 vssd1 vccd1 vccd1 _05566_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_67_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13621_ clknet_leaf_58_clk _00852_ net1132 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[609\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_81_2960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06774__B _01722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_2971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1484 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_2982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10426__A2 net1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09150__B _04053_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10764_ net1004 _05499_ _05500_ net1032 net1355 vssd1 vssd1 vccd1 vccd1 _00188_ sky130_fd_sc_hd__a32o_1
X_13552_ clknet_leaf_36_clk _00783_ net1236 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[540\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10296__B net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13323__CLK clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09292__A2 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_1700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_123 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12503_ _06165_ net348 net327 net1582 vssd1 vssd1 vccd1 vccd1 _01208_ sky130_fd_sc_hd__a22o_1
XFILLER_0_82_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13483_ clknet_leaf_53_clk _00714_ net1188 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[471\]
+ sky130_fd_sc_hd__dfrtp_1
X_10695_ net670 _05424_ _05434_ net965 _05433_ vssd1 vssd1 vccd1 vccd1 _05435_ sky130_fd_sc_hd__o221a_1
XFILLER_0_67_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11900__S net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12434_ net2110 net241 net335 vssd1 vssd1 vccd1 vccd1 _01141_ sky130_fd_sc_hd__mux2_1
XANTENNA__08481__S net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11387__B1 _05843_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12365_ net1882 net229 net269 vssd1 vssd1 vccd1 vccd1 _01076_ sky130_fd_sc_hd__mux2_1
XANTENNA__13473__CLK clknet_leaf_49_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_2753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_2130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_2764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14104_ clknet_leaf_24_clk _01301_ net1163 vssd1 vssd1 vccd1 vccd1 final_design.reqhand.instruction\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_11316_ net649 net585 net198 vssd1 vssd1 vccd1 vccd1 _06011_ sky130_fd_sc_hd__and3_1
XANTENNA__06802__A1 final_design.data_from_mem\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_2775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_2617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12296_ _05867_ _06260_ vssd1 vssd1 vccd1 vccd1 _06275_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_71_2628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_2639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14035_ clknet_leaf_40_clk _01266_ net1210 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[1023\]
+ sky130_fd_sc_hd__dfrtp_1
X_11247_ _04639_ _04653_ net652 vssd1 vssd1 vccd1 vccd1 _05950_ sky130_fd_sc_hd__a21o_1
XANTENNA__12351__A2 _06264_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07825__S net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11178_ net653 _05886_ _05888_ vssd1 vssd1 vccd1 vccd1 _05889_ sky130_fd_sc_hd__or3_1
XANTENNA__10362__B2 final_design.data_from_mem\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10129_ final_design.vga.v_current_state\[0\] _05034_ _04999_ vssd1 vssd1 vccd1 vccd1
+ _05035_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_69_2546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_2557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_2568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_69_2579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10665__A2 net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11590__B net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13819_ clknet_leaf_65_clk _01050_ net1072 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[807\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_4_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12178__S net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09807__A1 net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07340_ final_design.cpu.reg_window\[516\] final_design.cpu.reg_window\[548\] net900
+ vssd1 vssd1 vccd1 vccd1 _02291_ sky130_fd_sc_hd__mux2_1
XANTENNA__11614__A1 net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06716__S1 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07271_ final_design.cpu.reg_window\[198\] final_design.cpu.reg_window\[230\] net901
+ vssd1 vssd1 vccd1 vccd1 _02222_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_14_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09010_ _01364_ net1038 _03943_ vssd1 vssd1 vccd1 vccd1 _00225_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_14_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13816__CLK clknet_leaf_65_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11378__B1 _06064_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold102 final_design.reqhand.instruction\[8\] vssd1 vssd1 vccd1 vccd1 net1444 sky130_fd_sc_hd__dlygate4sd3_1
Xhold113 final_design.VGA_data_control.data_to_VGA\[17\] vssd1 vssd1 vccd1 vccd1 net1455
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold124 final_design.VGA_data_control.data_to_VGA\[18\] vssd1 vssd1 vccd1 vccd1 net1466
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09991__B1 net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12590__A2 net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold135 final_design.reqhand.instruction\[24\] vssd1 vssd1 vccd1 vccd1 net1477 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12840__CLK clknet_leaf_19_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold146 final_design.cpu.reg_window\[196\] vssd1 vssd1 vccd1 vccd1 net1488 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09418__S0 net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold157 final_design.cpu.reg_window\[723\] vssd1 vssd1 vccd1 vccd1 net1499 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13966__CLK clknet_leaf_45_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold168 final_design.reqhand.instruction\[0\] vssd1 vssd1 vccd1 vccd1 net1510 sky130_fd_sc_hd__dlygate4sd3_1
X_09912_ _04149_ _04830_ net447 vssd1 vssd1 vccd1 vccd1 _04831_ sky130_fd_sc_hd__a21oi_1
Xhold179 final_design.VGA_data_control.ready_data\[7\] vssd1 vssd1 vccd1 vccd1 net1521
+ sky130_fd_sc_hd__dlygate4sd3_1
Xfanout604 net605 vssd1 vssd1 vccd1 vccd1 net604 sky130_fd_sc_hd__buf_2
Xfanout615 net616 vssd1 vssd1 vccd1 vccd1 net615 sky130_fd_sc_hd__buf_2
Xfanout626 net627 vssd1 vssd1 vccd1 vccd1 net626 sky130_fd_sc_hd__buf_4
XFILLER_0_10_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12342__A2 net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout637 _06123_ vssd1 vssd1 vccd1 vccd1 net637 sky130_fd_sc_hd__clkbuf_4
X_09843_ _03230_ _04495_ net321 vssd1 vssd1 vccd1 vccd1 _04762_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08420__A net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout648 _05849_ vssd1 vssd1 vccd1 vccd1 net648 sky130_fd_sc_hd__buf_4
XANTENNA__10353__A1 net24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout291_A net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout659 _03649_ vssd1 vssd1 vccd1 vccd1 net659 sky130_fd_sc_hd__buf_4
XANTENNA_fanout389_A _06265_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06986_ net886 _01930_ _01936_ _01923_ _01924_ vssd1 vssd1 vccd1 vccd1 _01937_ sky130_fd_sc_hd__a32oi_4
X_09774_ net493 _04690_ _04692_ vssd1 vssd1 vccd1 vccd1 _04693_ sky130_fd_sc_hd__o21a_1
X_08725_ final_design.CPU_instr_adr\[17\] _01909_ vssd1 vssd1 vccd1 vccd1 _03676_
+ sky130_fd_sc_hd__nor2_1
XANTENNA__11302__B1 net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout556_A net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08656_ _01535_ _02572_ _03606_ vssd1 vssd1 vccd1 vccd1 _03607_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_7_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_54_clk_A clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13346__CLK clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06955__S1 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07607_ net711 _02551_ net724 vssd1 vssd1 vccd1 vccd1 _02558_ sky130_fd_sc_hd__o21ai_1
X_08587_ final_design.cpu.reg_window\[768\] final_design.cpu.reg_window\[800\] net827
+ vssd1 vssd1 vccd1 vccd1 _03538_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout723_A net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout344_X net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07538_ net755 _02482_ net747 vssd1 vssd1 vccd1 vccd1 _02489_ sky130_fd_sc_hd__o21a_1
XFILLER_0_14_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_12_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout511_X net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07469_ _01489_ _01495_ _01820_ _01817_ _01816_ vssd1 vssd1 vccd1 vccd1 _02420_ sky130_fd_sc_hd__a32oi_4
XANTENNA__13496__CLK clknet_leaf_65_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09208_ _04126_ _04123_ net262 vssd1 vssd1 vccd1 vccd1 _04127_ sky130_fd_sc_hd__and3b_1
X_10480_ _05228_ _05230_ _05221_ vssd1 vssd1 vccd1 vccd1 _05231_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12772__3_A clknet_leaf_25_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11369__B1 _06056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09139_ net538 net537 net535 net534 net456 net465 vssd1 vssd1 vccd1 vccd1 _04058_
+ sky130_fd_sc_hd__mux4_2
X_12150_ net198 net2389 net386 vssd1 vssd1 vccd1 vccd1 _00871_ sky130_fd_sc_hd__mux2_1
X_11101_ _05820_ _05821_ vssd1 vssd1 vccd1 vccd1 _05822_ sky130_fd_sc_hd__xnor2_1
XANTENNA__11956__A net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12081_ net2411 net393 net499 _06004_ vssd1 vssd1 vccd1 vccd1 _00806_ sky130_fd_sc_hd__a22o_1
XANTENNA__06891__S0 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold680 final_design.uart.working_data\[8\] vssd1 vssd1 vccd1 vccd1 net2022 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold691 final_design.cpu.reg_window\[264\] vssd1 vssd1 vccd1 vccd1 net2033 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11032_ _05748_ _05755_ vssd1 vssd1 vccd1 vccd1 _05756_ sky130_fd_sc_hd__nand2_1
XANTENNA__12333__A2 net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10344__B2 final_design.data_from_mem\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11541__B1 net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14121__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06643__S0 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09713__X _04632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12983_ net1314 _00214_ net1166 vssd1 vssd1 vccd1 vccd1 final_design.CPU_instr_adr\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_77_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11934_ _06135_ net278 net408 net2509 vssd1 vssd1 vccd1 vccd1 _00669_ sky130_fd_sc_hd__a22o_1
XFILLER_0_24_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11865_ net203 net554 vssd1 vssd1 vccd1 vccd1 _06243_ sky130_fd_sc_hd__and2_1
XANTENNA__13839__CLK clknet_leaf_42_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13604_ clknet_leaf_54_clk _00835_ net1177 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[592\]
+ sky130_fd_sc_hd__dfrtp_1
X_10816_ net77 _05529_ _05549_ vssd1 vssd1 vccd1 vccd1 _05550_ sky130_fd_sc_hd__a21bo_1
X_11796_ net649 _05869_ net198 vssd1 vssd1 vccd1 vccd1 _06235_ sky130_fd_sc_hd__and3_1
XFILLER_0_82_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09896__S0 net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07276__A1 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_1888 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13535_ clknet_leaf_8_clk _00766_ net1153 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[523\]
+ sky130_fd_sc_hd__dfrtp_1
X_10747_ _05467_ _05470_ vssd1 vssd1 vccd1 vccd1 _05484_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_77_2826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_2203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10678_ _05406_ _05414_ _05417_ net38 vssd1 vssd1 vccd1 vccd1 _05419_ sky130_fd_sc_hd__a31oi_2
XANTENNA__06724__S net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13466_ clknet_leaf_58_clk _00697_ net1122 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[454\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12863__CLK clknet_leaf_18_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_2837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_2848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13989__CLK clknet_leaf_49_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09100__S net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12417_ _06109_ net358 net340 net2136 vssd1 vssd1 vccd1 vccd1 _01127_ sky130_fd_sc_hd__a22o_1
XFILLER_0_2_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13397_ clknet_leaf_56_clk _00628_ net1149 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[385\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09973__B1 _04341_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12348_ net2287 net362 net351 _05990_ vssd1 vssd1 vccd1 vccd1 _01060_ sky130_fd_sc_hd__a22o_1
XFILLER_0_50_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13219__CLK clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12279_ net558 _06209_ net504 net368 net1780 vssd1 vssd1 vccd1 vccd1 _00994_ sky130_fd_sc_hd__a32o_1
XANTENNA__12461__S net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14018_ clknet_leaf_4_clk _01249_ net1080 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[1006\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10335__B2 final_design.data_from_mem\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06840_ final_design.cpu.reg_window\[340\] final_design.cpu.reg_window\[372\] net948
+ vssd1 vssd1 vccd1 vccd1 _01791_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13369__CLK clknet_leaf_55_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12088__A1 net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06771_ net742 net721 net665 vssd1 vssd1 vccd1 vccd1 _01722_ sky130_fd_sc_hd__a21o_2
X_08510_ final_design.cpu.reg_window\[386\] final_design.cpu.reg_window\[418\] net837
+ vssd1 vssd1 vccd1 vccd1 _03461_ sky130_fd_sc_hd__mux2_1
XANTENNA__08387__S0 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09490_ _04093_ _04340_ vssd1 vssd1 vccd1 vccd1 _04409_ sky130_fd_sc_hd__or2_1
XANTENNA__11296__C1 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08386__S net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_43 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08441_ final_design.cpu.reg_window\[324\] final_design.cpu.reg_window\[356\] net822
+ vssd1 vssd1 vccd1 vccd1 _03392_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08372_ _02212_ net598 vssd1 vssd1 vccd1 vccd1 _03323_ sky130_fd_sc_hd__and2_1
XFILLER_0_58_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11599__B1 net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07323_ final_design.cpu.reg_window\[388\] final_design.cpu.reg_window\[420\] net902
+ vssd1 vssd1 vccd1 vccd1 _02274_ sky130_fd_sc_hd__mux2_1
XANTENNA__11063__A2 _01371_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12260__A1 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07254_ final_design.cpu.reg_window\[711\] final_design.cpu.reg_window\[743\] net887
+ vssd1 vssd1 vccd1 vccd1 _02205_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_1185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12933__Q net157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07185_ final_design.cpu.reg_window\[201\] final_design.cpu.reg_window\[233\] net889
+ vssd1 vssd1 vccd1 vccd1 _02136_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_41_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_1873 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout304_A net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1046_A final_design.VGA_adr\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08767__A1 final_design.CPU_instr_adr\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11771__B1 net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12371__S net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14144__CLK clknet_leaf_19_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout401 _06257_ vssd1 vssd1 vccd1 vccd1 net401 sky130_fd_sc_hd__buf_4
XANTENNA__07465__S net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout412 net413 vssd1 vssd1 vccd1 vccd1 net412 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_6_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout423 net424 vssd1 vssd1 vccd1 vccd1 net423 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_6_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout434 net437 vssd1 vssd1 vccd1 vccd1 net434 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10326__B2 final_design.data_from_mem\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout294_X net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout445 net446 vssd1 vssd1 vccd1 vccd1 net445 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06589__B _01538_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout456 net457 vssd1 vssd1 vccd1 vccd1 net456 sky130_fd_sc_hd__clkbuf_4
X_09826_ net726 _04744_ vssd1 vssd1 vccd1 vccd1 _04745_ sky130_fd_sc_hd__nor2_1
XANTENNA__06625__S0 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout467 net468 vssd1 vssd1 vccd1 vccd1 net467 sky130_fd_sc_hd__buf_2
XANTENNA_fanout1001_X net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout478 net479 vssd1 vssd1 vccd1 vccd1 net478 sky130_fd_sc_hd__buf_2
Xfanout489 net490 vssd1 vssd1 vccd1 vccd1 net489 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12079__A1 net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout840_A net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout461_X net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09757_ net450 _04675_ _04672_ vssd1 vssd1 vccd1 vccd1 _04676_ sky130_fd_sc_hd__a21o_1
X_06969_ final_design.cpu.reg_window\[208\] final_design.cpu.reg_window\[240\] net926
+ vssd1 vssd1 vccd1 vccd1 _01920_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout938_A net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1833 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08708_ final_design.CPU_instr_adr\[28\] _01570_ vssd1 vssd1 vccd1 vccd1 _03659_
+ sky130_fd_sc_hd__xor2_1
X_09688_ _04434_ _04606_ net474 vssd1 vssd1 vccd1 vccd1 _04607_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_1877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09495__A2 net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08639_ _03586_ _03588_ vssd1 vssd1 vccd1 vccd1 _03590_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout726_X net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11650_ net430 net569 _06182_ net299 net1486 vssd1 vssd1 vccd1 vccd1 _00457_ sky130_fd_sc_hd__a32o_1
XANTENNA__12886__CLK clknet_leaf_17_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10601_ _05329_ _05345_ vssd1 vssd1 vccd1 vccd1 _05346_ sky130_fd_sc_hd__xor2_1
XANTENNA__12251__A1 net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11581_ net437 net579 _06146_ net304 net2027 vssd1 vssd1 vccd1 vccd1 _00424_ sky130_fd_sc_hd__a32o_1
XANTENNA__09652__C1 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10532_ net958 _05275_ _05279_ net955 vssd1 vssd1 vccd1 vccd1 _05280_ sky130_fd_sc_hd__o22a_1
X_13320_ clknet_leaf_41_clk _00551_ net1224 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[308\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1883 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10463_ net1473 net1032 _05215_ net249 vssd1 vssd1 vccd1 vccd1 _00172_ sky130_fd_sc_hd__a22o_1
X_13251_ clknet_leaf_0_clk _00482_ net1062 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[239\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_46_1913 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10014__B1 _04341_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07105__S1 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11357__A3 _06046_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12202_ net569 _06130_ net507 net377 net1556 vssd1 vssd1 vccd1 vccd1 _00920_ sky130_fd_sc_hd__a32o_1
XANTENNA__12554__A2 net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13182_ clknet_leaf_13_clk _00413_ net1089 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[170\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input67_A mem_adr_start[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10394_ _03613_ _04991_ _04987_ vssd1 vssd1 vccd1 vccd1 _05179_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_27_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12133_ net226 net2341 net384 vssd1 vssd1 vccd1 vccd1 _00854_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07981__A2 _02929_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12064_ net2443 net393 net500 _05876_ vssd1 vssd1 vccd1 vccd1 _00789_ sky130_fd_sc_hd__a22o_1
XANTENNA__13511__CLK clknet_leaf_63_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11015_ _05738_ _05739_ vssd1 vssd1 vccd1 vccd1 _05740_ sky130_fd_sc_hd__nand2_1
XANTENNA__09722__A3 net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout990 _01414_ vssd1 vssd1 vccd1 vccd1 net990 sky130_fd_sc_hd__buf_2
XANTENNA__13661__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12966_ clknet_leaf_32_clk _00204_ net1234 vssd1 vssd1 vccd1 vccd1 net125 sky130_fd_sc_hd__dfrtp_1
XANTENNA__06719__S net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09486__A2 net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1917 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1851 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11917_ net181 net2321 net275 vssd1 vssd1 vccd1 vccd1 _00656_ sky130_fd_sc_hd__mux2_1
X_12897_ clknet_leaf_20_clk _00135_ net1158 vssd1 vssd1 vccd1 vccd1 final_design.data_from_mem\[31\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_16_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_1737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11848_ _06098_ net281 net518 net2400 vssd1 vssd1 vccd1 vccd1 _00598_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_16_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14017__CLK clknet_leaf_47_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12797__28 clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 net1338 sky130_fd_sc_hd__inv_2
XFILLER_0_51_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12456__S net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11779_ net2397 net412 net276 _05911_ vssd1 vssd1 vccd1 vccd1 _00538_ sky130_fd_sc_hd__a22o_1
XFILLER_0_3_1461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11213__X _05920_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13518_ clknet_leaf_43_clk _00749_ net1218 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[506\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload11 clknet_leaf_63_clk vssd1 vssd1 vccd1 vccd1 clkload11/Y sky130_fd_sc_hd__bufinv_16
Xclkload22 clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 clkload22/Y sky130_fd_sc_hd__clkinv_8
X_13449_ clknet_leaf_36_clk _00680_ net1230 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[437\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13041__CLK clknet_leaf_34_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14167__CLK clknet_leaf_18_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload33 clknet_leaf_42_clk vssd1 vssd1 vccd1 vccd1 clkload33/Y sky130_fd_sc_hd__clkinv_2
XFILLER_0_45_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkload44 clknet_leaf_36_clk vssd1 vssd1 vccd1 vccd1 clkload44/Y sky130_fd_sc_hd__inv_6
XANTENNA__12545__A2 net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09765__S net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12191__S net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08990_ final_design.CPU_instr_adr\[15\] _03791_ final_design.CPU_instr_adr\[16\]
+ vssd1 vssd1 vccd1 vccd1 _03926_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08241__Y _03192_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07285__S net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13191__CLK clknet_leaf_62_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09066__A net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire739_A _01490_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07941_ _02888_ _02889_ _02890_ _02891_ net680 net692 vssd1 vssd1 vccd1 vccd1 _02892_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_76_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07872_ net711 _02822_ vssd1 vssd1 vccd1 vccd1 _02823_ sky130_fd_sc_hd__nor2_1
XANTENNA__06607__S0 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09611_ net86 _04193_ vssd1 vssd1 vccd1 vccd1 _04530_ sky130_fd_sc_hd__xnor2_4
X_06823_ final_design.cpu.reg_window\[981\] final_design.cpu.reg_window\[1013\] net938
+ vssd1 vssd1 vccd1 vccd1 _01774_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_30_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11535__S net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_3030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06754_ final_design.cpu.reg_window\[855\] final_design.cpu.reg_window\[887\] net931
+ vssd1 vssd1 vccd1 vccd1 _01705_ sky130_fd_sc_hd__mux2_1
X_09542_ net484 _04366_ _04460_ vssd1 vssd1 vccd1 vccd1 _04461_ sky130_fd_sc_hd__o21bai_2
XANTENNA__09513__B _04094_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_3041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_3052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06685_ final_design.cpu.reg_window\[409\] final_design.cpu.reg_window\[441\] net934
+ vssd1 vssd1 vccd1 vccd1 _01636_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09473_ _04171_ _04391_ vssd1 vssd1 vccd1 vccd1 _04392_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout254_A net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08424_ final_design.cpu.reg_window\[965\] final_design.cpu.reg_window\[997\] net840
+ vssd1 vssd1 vccd1 vccd1 _03375_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_955 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08355_ final_design.cpu.reg_window\[135\] final_design.cpu.reg_window\[167\] net806
+ vssd1 vssd1 vccd1 vccd1 _03306_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_28_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12366__S net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_24_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout421_A net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1163_A net1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout519_A net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07306_ final_design.cpu.reg_window\[965\] final_design.cpu.reg_window\[997\] net921
+ vssd1 vssd1 vccd1 vccd1 _02257_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_43_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload5 clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 clkload5/Y sky130_fd_sc_hd__clkinv_4
XTAP_TAPCELL_ROW_43_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08286_ _03233_ _03234_ _03235_ _03236_ net674 net696 vssd1 vssd1 vccd1 vccd1 _03237_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_43_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11992__B1 net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07237_ final_design.cpu.reg_window\[199\] final_design.cpu.reg_window\[231\] net887
+ vssd1 vssd1 vccd1 vccd1 _02188_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout307_X net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1049_X net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12536__A2 net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09937__B1 _04109_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07099__S0 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07168_ net750 _02118_ vssd1 vssd1 vccd1 vccd1 _02119_ sky130_fd_sc_hd__or2_1
XANTENNA__11744__A0 net221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout790_A _01418_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout888_A net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07948__C1 _01750_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07099_ _02046_ _02047_ _02048_ _02049_ net766 net786 vssd1 vssd1 vccd1 vccd1 _02050_
+ sky130_fd_sc_hd__mux4_1
Xfanout1207 net1212 vssd1 vssd1 vccd1 vccd1 net1207 sky130_fd_sc_hd__buf_2
Xfanout1218 net1221 vssd1 vssd1 vccd1 vccd1 net1218 sky130_fd_sc_hd__clkbuf_4
Xfanout220 net221 vssd1 vssd1 vccd1 vccd1 net220 sky130_fd_sc_hd__clkbuf_2
Xfanout1229 net1232 vssd1 vssd1 vccd1 vccd1 net1229 sky130_fd_sc_hd__clkbuf_4
Xfanout231 net232 vssd1 vssd1 vccd1 vccd1 net231 sky130_fd_sc_hd__buf_2
XANTENNA_fanout676_X net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout242 _05875_ vssd1 vssd1 vccd1 vccd1 net242 sky130_fd_sc_hd__buf_2
Xfanout253 _04961_ vssd1 vssd1 vccd1 vccd1 net253 sky130_fd_sc_hd__clkbuf_8
XANTENNA__13684__CLK clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout264 net265 vssd1 vssd1 vccd1 vccd1 net264 sky130_fd_sc_hd__buf_4
Xfanout275 _06247_ vssd1 vssd1 vccd1 vccd1 net275 sky130_fd_sc_hd__clkbuf_8
XANTENNA__08373__C1 _02211_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout286 net287 vssd1 vssd1 vccd1 vccd1 net286 sky130_fd_sc_hd__clkbuf_2
Xfanout297 _06194_ vssd1 vssd1 vccd1 vccd1 net297 sky130_fd_sc_hd__buf_4
X_09809_ _04727_ vssd1 vssd1 vccd1 vccd1 _04728_ sky130_fd_sc_hd__inv_2
XANTENNA__11445__S net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1630 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12820_ net1382 vssd1 vssd1 vccd1 vccd1 _00261_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_69_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09423__B _04341_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12751_ _06351_ _06372_ net954 _05058_ vssd1 vssd1 vccd1 vccd1 _06389_ sky130_fd_sc_hd__and4b_1
XFILLER_0_69_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_1084 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11702_ net557 net420 _06209_ net294 net1634 vssd1 vssd1 vccd1 vccd1 _00482_ sky130_fd_sc_hd__a32o_1
X_12682_ _06328_ net1391 net981 vssd1 vssd1 vccd1 vccd1 _01343_ sky130_fd_sc_hd__mux2_1
XANTENNA__12224__A1 net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11633_ net207 net630 vssd1 vssd1 vccd1 vccd1 _06174_ sky130_fd_sc_hd__and2_1
XANTENNA__13064__CLK clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08979__A1 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08523__S0 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11564_ net209 net636 vssd1 vssd1 vccd1 vccd1 _06138_ sky130_fd_sc_hd__and2_1
XFILLER_0_37_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11983__B1 net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13303_ clknet_leaf_6_clk _00534_ net1132 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[291\]
+ sky130_fd_sc_hd__dfrtp_1
X_10515_ _05250_ _05260_ _05262_ net61 vssd1 vssd1 vccd1 vccd1 _05264_ sky130_fd_sc_hd__a31o_1
XANTENNA__07651__A1 net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11495_ net179 net2365 net308 vssd1 vssd1 vccd1 vccd1 _00369_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_1612 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09928__B1 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12527__A2 net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10446_ _02863_ net592 vssd1 vssd1 vccd1 vccd1 _05207_ sky130_fd_sc_hd__nor2_1
X_13234_ clknet_leaf_39_clk _00465_ net1205 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[222\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10377_ net20 net1025 net1008 final_design.data_from_mem\[26\] vssd1 vssd1 vccd1
+ vccd1 _00130_ sky130_fd_sc_hd__a22o_1
X_13165_ clknet_leaf_48_clk _00396_ net1202 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[153\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08600__B1 _02423_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12901__CLK clknet_leaf_25_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12116_ net1790 net196 net390 vssd1 vssd1 vccd1 vccd1 _00840_ sky130_fd_sc_hd__mux2_1
X_13096_ clknet_leaf_35_clk _00327_ net1240 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[84\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09156__A1 net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12047_ net1668 net198 net398 vssd1 vssd1 vccd1 vccd1 _00775_ sky130_fd_sc_hd__mux2_1
XANTENNA__11863__B net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07405__Y _02356_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1861 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13998_ clknet_leaf_43_clk _01229_ net1222 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[986\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08116__C1 net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12949_ clknet_leaf_29_clk _00187_ net1194 vssd1 vssd1 vccd1 vccd1 net106 sky130_fd_sc_hd__dfrtp_1
XANTENNA__11266__A2 net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13407__CLK clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1889 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06470_ final_design.reqhand.instruction\[16\] net969 vssd1 vssd1 vccd1 vccd1 _01421_
+ sky130_fd_sc_hd__and2_1
XANTENNA__12215__A1 net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12186__S net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08140_ final_design.cpu.reg_window\[781\] final_design.cpu.reg_window\[813\] net855
+ vssd1 vssd1 vccd1 vccd1 _03091_ sky130_fd_sc_hd__mux2_1
XANTENNA__07140__Y _02091_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13557__CLK clknet_leaf_57_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11974__B1 net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08071_ net879 _03021_ _03010_ _03009_ vssd1 vssd1 vccd1 vccd1 _03022_ sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_43_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12518__A2 net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07022_ final_design.cpu.reg_window\[462\] final_design.cpu.reg_window\[494\] net897
+ vssd1 vssd1 vccd1 vccd1 _01973_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11726__B1 net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkload39_A clknet_leaf_30_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07945__A2 _02894_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08973_ final_design.CPU_instr_adr\[18\] net1016 _03908_ _03910_ vssd1 vssd1 vccd1
+ vccd1 _00229_ sky130_fd_sc_hd__a22o_1
Xhold17 final_design.cpu.reg_window\[5\] vssd1 vssd1 vccd1 vccd1 net1359 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_32_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07924_ net710 _02874_ vssd1 vssd1 vccd1 vccd1 _02875_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_32_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold28 final_design.cpu.reg_window\[21\] vssd1 vssd1 vccd1 vccd1 net1370 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_51_1936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold39 net118 vssd1 vssd1 vccd1 vccd1 net1381 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12151__A0 _06017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1009_A _05166_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07253__S0 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07855_ final_design.cpu.reg_window\[340\] final_design.cpu.reg_window\[372\] net868
+ vssd1 vssd1 vccd1 vccd1 _02806_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout371_A _06274_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout469_A _03518_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06806_ net551 _01755_ vssd1 vssd1 vccd1 vccd1 _01757_ sky130_fd_sc_hd__or2_1
X_07786_ _02734_ _02736_ vssd1 vssd1 vccd1 vccd1 _02737_ sky130_fd_sc_hd__nor2_1
XFILLER_0_79_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09525_ _04116_ _04443_ _04442_ net320 vssd1 vssd1 vccd1 vccd1 _04444_ sky130_fd_sc_hd__a2bb2o_1
X_06737_ net877 vssd1 vssd1 vccd1 vccd1 _01688_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13087__CLK clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10465__A0 final_design.CPU_instr_adr\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout257_X net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_63_clk clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_63_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout636_A net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07979__A net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06668_ net753 _01618_ vssd1 vssd1 vccd1 vccd1 _01619_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_26_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09456_ net479 _04302_ _04374_ net319 vssd1 vssd1 vccd1 vccd1 _04375_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_49_1898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08407_ _03355_ _03357_ vssd1 vssd1 vccd1 vccd1 _03358_ sky130_fd_sc_hd__or2_2
XFILLER_0_4_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12096__S net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout424_X net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09387_ net491 _04305_ vssd1 vssd1 vccd1 vccd1 _04306_ sky130_fd_sc_hd__or2_1
X_06599_ final_design.cpu.reg_window\[476\] final_design.cpu.reg_window\[508\] net946
+ vssd1 vssd1 vccd1 vccd1 _01550_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout1166_X net1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07308__S1 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08338_ net598 _03287_ _03263_ vssd1 vssd1 vccd1 vccd1 _03289_ sky130_fd_sc_hd__o21a_1
XANTENNA__09622__A2 net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11965__B1 net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08269_ final_design.cpu.reg_window\[586\] final_design.cpu.reg_window\[618\] net815
+ vssd1 vssd1 vccd1 vccd1 _03220_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12924__CLK clknet_leaf_49_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10300_ final_design.VGA_data_control.data_to_VGA\[11\] final_design.VGA_data_control.data_to_VGA\[10\]
+ final_design.VGA_data_control.data_to_VGA\[9\] final_design.VGA_data_control.data_to_VGA\[8\]
+ net1050 net1049 vssd1 vssd1 vccd1 vccd1 _05154_ sky130_fd_sc_hd__mux4_1
XANTENNA__12963__RESET_B net1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12509__A2 net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11280_ _04681_ _04696_ net652 vssd1 vssd1 vccd1 vccd1 _05979_ sky130_fd_sc_hd__a21o_1
XANTENNA__10852__B net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout793_X net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10231_ final_design.uart.BAUD_counter\[11\] final_design.uart.BAUD_counter\[10\]
+ _05104_ vssd1 vssd1 vccd1 vccd1 _05108_ sky130_fd_sc_hd__and3_1
XANTENNA__06819__S0 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11193__A1 final_design.data_from_mem\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10162_ final_design.VGA_data_control.VGA_request_address\[0\] _05054_ _05056_ vssd1
+ vssd1 vccd1 vccd1 final_design.vga.h_next_count\[6\] sky130_fd_sc_hd__o21a_1
XANTENNA__11018__A2_N _05239_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07219__A net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout960_X net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1004 _05173_ vssd1 vssd1 vccd1 vccd1 net1004 sky130_fd_sc_hd__clkbuf_2
Xfanout1015 net1017 vssd1 vssd1 vccd1 vccd1 net1015 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09138__A1 net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1026 _05168_ vssd1 vssd1 vccd1 vccd1 net1026 sky130_fd_sc_hd__clkbuf_2
X_10093_ final_design.VGA_data_control.h_count\[8\] final_design.VGA_data_control.h_count\[9\]
+ vssd1 vssd1 vccd1 vccd1 _05009_ sky130_fd_sc_hd__nor2_1
Xfanout1037 _01410_ vssd1 vssd1 vccd1 vccd1 net1037 sky130_fd_sc_hd__buf_4
Xfanout1048 final_design.VGA_data_control.h_count\[4\] vssd1 vssd1 vccd1 vccd1 net1048
+ sky130_fd_sc_hd__clkbuf_2
XANTENNA__12142__A0 net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1059 net1060 vssd1 vssd1 vccd1 vccd1 net1059 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11683__B net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13921_ clknet_leaf_47_clk _01152_ net1203 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[909\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13852_ clknet_leaf_5_clk _01083_ net1083 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[840\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09153__B net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_1179 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12803_ net1386 vssd1 vssd1 vccd1 vccd1 _00244_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_74_1471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13783_ clknet_leaf_6_clk _01014_ net1129 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[771\]
+ sky130_fd_sc_hd__dfrtp_1
X_10995_ net86 _05698_ _05720_ vssd1 vssd1 vccd1 vccd1 _05721_ sky130_fd_sc_hd__a21o_1
Xclkbuf_leaf_54_clk clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_54_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__11903__S net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12734_ _06364_ _06367_ _06368_ final_design.VGA_data_control.v_count\[0\] vssd1
+ vssd1 vccd1 vccd1 _06375_ sky130_fd_sc_hd__o22a_1
XANTENNA__08484__S net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12665_ final_design.VGA_data_control.ready_data\[20\] net1019 net974 final_design.data_from_mem\[20\]
+ vssd1 vssd1 vccd1 vccd1 _06320_ sky130_fd_sc_hd__a22o_1
XFILLER_0_38_763 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_2276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_1753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_2287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12748__A2 _05058_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_2298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11616_ net569 net422 _06165_ net299 net1467 vssd1 vssd1 vccd1 vccd1 _00440_ sky130_fd_sc_hd__a32o_1
X_12596_ net1662 net998 net984 final_design.data_from_mem\[14\] vssd1 vssd1 vccd1
+ vccd1 _01289_ sky130_fd_sc_hd__a22o_1
XFILLER_0_13_1797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1242 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07624__A1 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11547_ net2531 net302 _06129_ net421 vssd1 vssd1 vccd1 vccd1 _00407_ sky130_fd_sc_hd__a22o_1
XFILLER_0_41_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_1475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold509 final_design.cpu.reg_window\[522\] vssd1 vssd1 vccd1 vccd1 net1851 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06732__S net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11858__B net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11478_ net197 net640 vssd1 vssd1 vccd1 vccd1 _06109_ sky130_fd_sc_hd__and2_1
XANTENNA__11708__B1 net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09377__A1 net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13217_ clknet_leaf_49_clk _00448_ net1184 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[205\]
+ sky130_fd_sc_hd__dfrtp_1
X_10429_ net526 _05190_ vssd1 vssd1 vccd1 vccd1 _05198_ sky130_fd_sc_hd__nor2_1
X_14197_ net1255 vssd1 vssd1 vccd1 vccd1 gpio_oeb[9] sky130_fd_sc_hd__buf_2
XFILLER_0_42_1415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13148_ clknet_leaf_3_clk _00379_ net1068 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[136\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10931__A1 net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10931__B2 net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13079_ clknet_leaf_5_clk _00310_ net1082 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[67\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1209 net166 vssd1 vssd1 vccd1 vccd1 net2551 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_75_1213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07640_ final_design.cpu.reg_window\[796\] final_design.cpu.reg_window\[828\] net866
+ vssd1 vssd1 vccd1 vccd1 _02591_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_0_217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_0_228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12436__A1 net240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07571_ final_design.cpu.reg_window\[95\] final_design.cpu.reg_window\[127\] net857
+ vssd1 vssd1 vccd1 vccd1 _02522_ sky130_fd_sc_hd__mux2_1
XANTENNA__11239__A2 net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_45_clk clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_45_clk sky130_fd_sc_hd__clkbuf_8
X_06522_ _01466_ _01467_ _01471_ _01472_ vssd1 vssd1 vccd1 vccd1 _01473_ sky130_fd_sc_hd__nor4_1
XANTENNA__11813__S net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09310_ _04226_ _04228_ vssd1 vssd1 vccd1 vccd1 _04229_ sky130_fd_sc_hd__nand2_1
XANTENNA__07799__A net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06453_ _01405_ _01406_ _01396_ vssd1 vssd1 vccd1 vccd1 _00001_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_5_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09241_ _04159_ vssd1 vssd1 vccd1 vccd1 _04160_ sky130_fd_sc_hd__inv_2
XANTENNA__12947__CLK clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09172_ _03635_ net659 vssd1 vssd1 vccd1 vccd1 _04091_ sky130_fd_sc_hd__nor2_1
XFILLER_0_7_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08123_ final_design.cpu.reg_window\[397\] final_design.cpu.reg_window\[429\] net854
+ vssd1 vssd1 vccd1 vccd1 _03074_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11947__B1 net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout217_A _05934_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08054_ final_design.cpu.reg_window\[18\] final_design.cpu.reg_window\[50\] net844
+ vssd1 vssd1 vccd1 vccd1 _03005_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_38_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12781__12 clknet_leaf_28_clk vssd1 vssd1 vccd1 vccd1 net1322 sky130_fd_sc_hd__inv_2
XFILLER_0_64_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07005_ final_design.cpu.reg_window\[783\] final_design.cpu.reg_window\[815\] net892
+ vssd1 vssd1 vccd1 vccd1 _01956_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_38_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xmax_cap740 _01484_ vssd1 vssd1 vccd1 vccd1 net740 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_38_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_1635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_983 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07379__B1 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1126_A net1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08040__A1 net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout586_A net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11784__A net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08956_ _03671_ _03672_ vssd1 vssd1 vccd1 vccd1 _03895_ sky130_fd_sc_hd__nand2_1
X_07907_ final_design.cpu.reg_window\[663\] final_design.cpu.reg_window\[695\] net848
+ vssd1 vssd1 vccd1 vccd1 _02858_ sky130_fd_sc_hd__mux2_1
XANTENNA__12675__B2 final_design.data_from_mem\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08887_ _01600_ _01601_ _02472_ vssd1 vssd1 vccd1 vccd1 _03834_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout374_X net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout753_A net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07838_ final_design.cpu.reg_window\[917\] final_design.cpu.reg_window\[949\] net860
+ vssd1 vssd1 vccd1 vccd1 _02789_ sky130_fd_sc_hd__mux2_1
XANTENNA__10150__A2 net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout920_A net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07769_ final_design.cpu.reg_window\[856\] final_design.cpu.reg_window\[888\] net864
+ vssd1 vssd1 vccd1 vccd1 _02720_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_36_clk clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_36_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout639_X net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09508_ _02934_ _03587_ _04426_ _03029_ _02932_ vssd1 vssd1 vccd1 vccd1 _04427_ sky130_fd_sc_hd__a311o_1
XANTENNA__09701__B _04619_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10780_ _05514_ _05515_ vssd1 vssd1 vccd1 vccd1 _05516_ sky130_fd_sc_hd__and2_1
XFILLER_0_78_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07303__B1 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09439_ _04191_ _04357_ vssd1 vssd1 vccd1 vccd1 _04358_ sky130_fd_sc_hd__nand2_1
XANTENNA__07854__A1 _01504_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11650__A2 net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13872__CLK clknet_leaf_34_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12450_ net1632 net202 net336 vssd1 vssd1 vccd1 vccd1 _01157_ sky130_fd_sc_hd__mux2_1
XANTENNA__11938__B1 net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11401_ final_design.data_from_mem\[31\] net236 net234 vssd1 vssd1 vccd1 vccd1 _06085_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_1_1773 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12381_ net2073 net203 net270 vssd1 vssd1 vccd1 vccd1 _01092_ sky130_fd_sc_hd__mux2_1
XANTENNA__11402__A2 _05946_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1584 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14120_ clknet_leaf_21_clk final_design.vga.v_next_count\[0\] net1159 vssd1 vssd1
+ vccd1 vccd1 final_design.VGA_data_control.v_count\[0\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__07648__S net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11332_ net648 net570 net194 vssd1 vssd1 vccd1 vccd1 _06025_ sky130_fd_sc_hd__and3_1
XANTENNA__13102__CLK clknet_leaf_45_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14051_ clknet_leaf_16_clk _00012_ net1093 vssd1 vssd1 vccd1 vccd1 final_design.uart.BAUD_counter\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_11263_ net644 _05960_ _05963_ vssd1 vssd1 vccd1 vccd1 _05964_ sky130_fd_sc_hd__a21o_1
XANTENNA__11166__A1 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09863__S net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13002_ net1333 _00233_ net1196 vssd1 vssd1 vccd1 vccd1 final_design.CPU_instr_adr\[22\]
+ sky130_fd_sc_hd__dfrtp_4
X_10214_ final_design.uart.BAUD_counter\[3\] final_design.uart.BAUD_counter\[4\] _05093_
+ final_design.uart.BAUD_counter\[5\] vssd1 vssd1 vccd1 vccd1 _05097_ sky130_fd_sc_hd__a31o_1
X_11194_ net653 _05900_ _05902_ vssd1 vssd1 vccd1 vccd1 _05903_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_73_2692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10145_ _05016_ _05045_ vssd1 vssd1 vccd1 vccd1 _05046_ sky130_fd_sc_hd__or2_1
XANTENNA__13252__CLK clknet_leaf_54_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08479__S net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07383__S net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10076_ net801 _04988_ _04992_ _01373_ vssd1 vssd1 vccd1 vccd1 _04993_ sky130_fd_sc_hd__a211oi_2
XANTENNA__09531__A1 net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13904_ clknet_leaf_33_clk _01135_ net1239 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[892\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_72_1408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13835_ clknet_leaf_52_clk _01066_ net1185 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[823\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_67_2485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_27_clk clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_27_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_67_2496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_63_2349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06727__S net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13766_ clknet_leaf_50_clk _00997_ net1173 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[754\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10978_ final_design.CPU_instr_adr\[25\] _03854_ net1059 vssd1 vssd1 vccd1 vccd1
+ _05705_ sky130_fd_sc_hd__mux2_1
XANTENNA__09834__A2 _04087_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12717_ _06347_ _06357_ _06349_ vssd1 vssd1 vccd1 vccd1 _06358_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_2_1504 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06648__A2 _01598_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13697_ clknet_leaf_47_clk _00928_ net1199 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[685\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09256__B1_N _02545_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12648_ _06311_ net1406 net978 vssd1 vssd1 vccd1 vccd1 _01326_ sky130_fd_sc_hd__mux2_1
XANTENNA__11929__B1 net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12579_ net2022 _06294_ _06286_ vssd1 vssd1 vccd1 vccd1 _01274_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_1657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11588__B net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold306 final_design.cpu.reg_window\[523\] vssd1 vssd1 vccd1 vccd1 net1648 sky130_fd_sc_hd__dlygate4sd3_1
Xhold317 final_design.cpu.reg_window\[576\] vssd1 vssd1 vccd1 vccd1 net1659 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold328 final_design.cpu.reg_window\[683\] vssd1 vssd1 vccd1 vccd1 net1670 sky130_fd_sc_hd__dlygate4sd3_1
Xhold339 final_design.cpu.reg_window\[985\] vssd1 vssd1 vccd1 vccd1 net1681 sky130_fd_sc_hd__dlygate4sd3_1
X_14249_ net1303 vssd1 vssd1 vccd1 vccd1 gpio_out[27] sky130_fd_sc_hd__buf_2
XFILLER_0_61_1813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11157__A1 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12354__B1 net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout808 net809 vssd1 vssd1 vccd1 vccd1 net808 sky130_fd_sc_hd__clkbuf_2
Xfanout819 net824 vssd1 vssd1 vccd1 vccd1 net819 sky130_fd_sc_hd__clkbuf_4
X_08810_ final_design.CPU_instr_adr\[21\] _01788_ vssd1 vssd1 vccd1 vccd1 _03761_
+ sky130_fd_sc_hd__or2_1
X_09790_ net491 _04607_ vssd1 vssd1 vccd1 vccd1 _04709_ sky130_fd_sc_hd__nand2_1
XANTENNA__06584__A1 net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10380__A2 net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1006 final_design.cpu.reg_window\[543\] vssd1 vssd1 vccd1 vccd1 net2348 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1017 final_design.cpu.reg_window\[631\] vssd1 vssd1 vccd1 vccd1 net2359 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07146__X _02097_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08741_ _03690_ _03691_ vssd1 vssd1 vccd1 vccd1 _03692_ sky130_fd_sc_hd__nor2_1
XFILLER_0_20_1554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1028 final_design.cpu.reg_window\[127\] vssd1 vssd1 vccd1 vccd1 net2370 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13745__CLK clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12657__B2 final_design.data_from_mem\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1039 final_design.cpu.reg_window\[401\] vssd1 vssd1 vccd1 vccd1 net2381 sky130_fd_sc_hd__dlygate4sd3_1
X_08672_ _01501_ _01505_ _01537_ _02028_ vssd1 vssd1 vccd1 vccd1 _03623_ sky130_fd_sc_hd__or4_1
XFILLER_0_75_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07623_ _01536_ _02572_ vssd1 vssd1 vccd1 vccd1 _02574_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_5_Right_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11880__A2 net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_18_clk clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_18_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_36_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13895__CLK clknet_leaf_59_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07554_ net527 _02504_ vssd1 vssd1 vccd1 vccd1 _02505_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10667__B final_design.VGA_adr\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06505_ _01454_ _01455_ vssd1 vssd1 vccd1 vccd1 _01456_ sky130_fd_sc_hd__nand2_1
XANTENNA__09381__S0 net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07485_ _02269_ _02434_ _02268_ vssd1 vssd1 vccd1 vccd1 _02436_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11632__A2 net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout334_A net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1076_A net1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09224_ _04142_ vssd1 vssd1 vccd1 vccd1 _04143_ sky130_fd_sc_hd__inv_2
X_06436_ net1051 vssd1 vssd1 vccd1 vccd1 _01391_ sky130_fd_sc_hd__inv_2
XANTENNA__13125__CLK clknet_leaf_49_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_744 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07049__C1 _01821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12374__S net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09155_ _04054_ net320 vssd1 vssd1 vccd1 vccd1 _04074_ sky130_fd_sc_hd__nand2_2
XANTENNA_fanout501_A _06264_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1243_A net1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12593__B1 net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08106_ final_design.cpu.reg_window\[908\] final_design.cpu.reg_window\[940\] net816
+ vssd1 vssd1 vccd1 vccd1 _03057_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08261__A1 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11498__B _06116_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09086_ net254 _04009_ _04010_ _04007_ vssd1 vssd1 vccd1 vccd1 _04011_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_20_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08037_ final_design.cpu.reg_window\[531\] final_design.cpu.reg_window\[563\] net822
+ vssd1 vssd1 vccd1 vccd1 _02988_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold840 final_design.reqhand.instruction\[31\] vssd1 vssd1 vccd1 vccd1 net2182 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold851 final_design.cpu.reg_window\[808\] vssd1 vssd1 vccd1 vccd1 net2193 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12345__B1 net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold862 final_design.cpu.reg_window\[381\] vssd1 vssd1 vccd1 vccd1 net2204 sky130_fd_sc_hd__dlygate4sd3_1
Xhold873 final_design.cpu.reg_window\[925\] vssd1 vssd1 vccd1 vccd1 net2215 sky130_fd_sc_hd__dlygate4sd3_1
Xhold884 final_design.cpu.reg_window\[325\] vssd1 vssd1 vccd1 vccd1 net2226 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout870_A net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold895 final_design.cpu.reg_window\[397\] vssd1 vssd1 vccd1 vccd1 net2237 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_10_Left_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout589_X net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09988_ _02737_ _04165_ vssd1 vssd1 vccd1 vccd1 _04907_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_60_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10371__A2 net1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08939_ final_design.CPU_instr_adr\[22\] net1014 _03876_ _03880_ vssd1 vssd1 vccd1
+ vccd1 _00233_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_4_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout756_X net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13343__RESET_B net1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11950_ _06151_ net291 net410 net2068 vssd1 vssd1 vccd1 vccd1 _00685_ sky130_fd_sc_hd__a22o_1
XFILLER_0_73_1717 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11320__A1 final_design.data_from_mem\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10901_ net82 net1046 vssd1 vssd1 vccd1 vccd1 _05631_ sky130_fd_sc_hd__or2_1
XANTENNA__11871__A2 net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11881_ _06115_ net290 net519 final_design.cpu.reg_window\[382\] vssd1 vssd1 vccd1
+ vccd1 _00625_ sky130_fd_sc_hd__a22o_1
XANTENNA__11453__S net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13620_ clknet_leaf_8_clk _00851_ net1154 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[608\]
+ sky130_fd_sc_hd__dfrtp_1
X_10832_ _05564_ _05565_ net1404 net1032 vssd1 vssd1 vccd1 vccd1 _00191_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_32_1403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_2961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_2972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07232__A net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13551_ clknet_leaf_39_clk _00782_ net1208 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[539\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_81_2983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10763_ _05477_ _05481_ _05498_ vssd1 vssd1 vccd1 vccd1 _05500_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_71_1496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12502_ _06164_ net343 net326 net1781 vssd1 vssd1 vccd1 vccd1 _01207_ sky130_fd_sc_hd__a22o_1
XFILLER_0_81_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10831__B1 net1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input97_A memory_size[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13482_ clknet_leaf_51_clk _00713_ net1170 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[470\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_135 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10694_ net1054 _05430_ net1001 final_design.CPU_instr_adr\[12\] vssd1 vssd1 vccd1
+ vccd1 _05434_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__14050__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12433_ net1567 net229 net335 vssd1 vssd1 vccd1 vccd1 _01140_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_179 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13618__CLK clknet_leaf_38_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11387__A1 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12584__B1 net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_2890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12364_ net1869 net231 net269 vssd1 vssd1 vccd1 vccd1 _01075_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_56_2120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_2754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14103_ clknet_leaf_24_clk _01300_ net1163 vssd1 vssd1 vccd1 vccd1 final_design.reqhand.instruction\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_56_2131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_2765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11315_ _04953_ net652 net590 _06009_ vssd1 vssd1 vccd1 vccd1 _06010_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_75_2776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_2618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12295_ net579 _06225_ net511 net370 net1965 vssd1 vssd1 vccd1 vccd1 _01010_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_71_2629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12336__B1 net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14034_ clknet_leaf_39_clk _01265_ net1207 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[1022\]
+ sky130_fd_sc_hd__dfrtp_1
X_11246_ net644 _05943_ _05948_ vssd1 vssd1 vccd1 vccd1 _05949_ sky130_fd_sc_hd__a21o_1
XANTENNA__13768__CLK clknet_leaf_40_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11177_ final_design.data_from_mem\[4\] net251 _05855_ _05887_ vssd1 vssd1 vccd1
+ vccd1 _05888_ sky130_fd_sc_hd__o211a_1
XANTENNA__10362__A2 net1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10128_ final_design.vga.v_current_state\[1\] _04997_ vssd1 vssd1 vccd1 vccd1 _05034_
+ sky130_fd_sc_hd__nand2_1
XANTENNA__13084__RESET_B net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_2547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10059_ _04571_ _04573_ _04632_ _04634_ vssd1 vssd1 vccd1 vccd1 _04978_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_69_2558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_2569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13013__RESET_B net1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12459__S net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11862__A2 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13818_ clknet_leaf_63_clk _01049_ net1121 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[806\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_1612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13148__CLK clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09807__A2 _04366_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07142__A _01468_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11614__A2 net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13749_ clknet_leaf_58_clk _00980_ net1133 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[737\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07270_ net751 _02220_ vssd1 vssd1 vccd1 vccd1 _02221_ sky130_fd_sc_hd__nor2_1
XFILLER_0_2_1334 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_14_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12194__S net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13298__CLK clknet_leaf_38_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11378__A1 _01570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11378__B2 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07677__S0 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold103 final_design.VGA_data_control.data_to_VGA\[22\] vssd1 vssd1 vccd1 vccd1 net1445
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold114 net165 vssd1 vssd1 vccd1 vccd1 net1456 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11111__B net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold125 final_design.cpu.reg_window\[197\] vssd1 vssd1 vccd1 vccd1 net1467 sky130_fd_sc_hd__dlygate4sd3_1
Xhold136 final_design.VGA_data_control.ready_data\[0\] vssd1 vssd1 vccd1 vccd1 net1478
+ sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_7_clk clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_7_clk sky130_fd_sc_hd__clkbuf_8
Xhold147 final_design.cpu.reg_window\[715\] vssd1 vssd1 vccd1 vccd1 net1489 sky130_fd_sc_hd__dlygate4sd3_1
Xhold158 net161 vssd1 vssd1 vccd1 vccd1 net1500 sky130_fd_sc_hd__dlygate4sd3_1
X_09911_ _03423_ _04148_ vssd1 vssd1 vccd1 vccd1 _04830_ sky130_fd_sc_hd__or2_1
Xhold169 final_design.VGA_data_control.ready_data\[5\] vssd1 vssd1 vccd1 vccd1 net1511
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkload21_A clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout605 net606 vssd1 vssd1 vccd1 vccd1 net605 sky130_fd_sc_hd__clkbuf_4
Xfanout616 net617 vssd1 vssd1 vccd1 vccd1 net616 sky130_fd_sc_hd__buf_2
Xfanout627 _06192_ vssd1 vssd1 vccd1 vccd1 net627 sky130_fd_sc_hd__clkbuf_4
X_09842_ _03230_ _04495_ vssd1 vssd1 vccd1 vccd1 _04761_ sky130_fd_sc_hd__or2_1
XFILLER_0_61_1687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout638 net639 vssd1 vssd1 vccd1 vccd1 net638 sky130_fd_sc_hd__buf_4
Xfanout649 net650 vssd1 vssd1 vccd1 vccd1 net649 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10353__A2 net1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08071__A1_N net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08951__C1 net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09773_ net480 _04406_ _04691_ net485 vssd1 vssd1 vccd1 vccd1 _04692_ sky130_fd_sc_hd__a211o_1
X_06985_ net763 _01935_ vssd1 vssd1 vccd1 vccd1 _01936_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout284_A _06228_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08724_ _03673_ _03674_ vssd1 vssd1 vccd1 vccd1 _03675_ sky130_fd_sc_hd__nand2_1
XANTENNA__11302__A1 final_design.data_from_mem\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08655_ _01566_ _02576_ _02604_ vssd1 vssd1 vccd1 vccd1 _03606_ sky130_fd_sc_hd__or3_1
XANTENNA__11853__A2 net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12369__S net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout451_A _04069_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1193_A net1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout549_A _01815_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07606_ net719 _02556_ vssd1 vssd1 vccd1 vccd1 _02557_ sky130_fd_sc_hd__nor2_1
XFILLER_0_37_1881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08586_ final_design.cpu.reg_window\[832\] final_design.cpu.reg_window\[864\] net835
+ vssd1 vssd1 vccd1 vccd1 _03537_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14073__CLK clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07537_ net762 _02487_ vssd1 vssd1 vccd1 vccd1 _02488_ sky130_fd_sc_hd__or2_1
XFILLER_0_7_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout337_X net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout716_A net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07468_ _02406_ _02407_ _02418_ net881 vssd1 vssd1 vccd1 vccd1 _02419_ sky130_fd_sc_hd__a22oi_4
XFILLER_0_68_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09207_ _02545_ _03608_ _04052_ _04125_ _03610_ vssd1 vssd1 vccd1 vccd1 _04126_ sky130_fd_sc_hd__o311a_1
X_06419_ final_design.reqhand.instruction\[2\] vssd1 vssd1 vccd1 vccd1 _01374_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout504_X net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07399_ final_design.cpu.reg_window\[706\] final_design.cpu.reg_window\[738\] net913
+ vssd1 vssd1 vccd1 vccd1 _02350_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11369__B2 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09138_ net542 net541 net540 net539 net459 net469 vssd1 vssd1 vccd1 vccd1 _04057_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_60_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13910__CLK clknet_leaf_59_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09069_ _02438_ net622 _03991_ net254 vssd1 vssd1 vccd1 vccd1 _03996_ sky130_fd_sc_hd__a31o_1
X_11100_ net92 _05802_ vssd1 vssd1 vccd1 vccd1 _05821_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_44_1841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12080_ net573 _05997_ net508 net395 net1829 vssd1 vssd1 vccd1 vccd1 _00805_ sky130_fd_sc_hd__a32o_1
XANTENNA__06830__S net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06891__S1 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold670 final_design.cpu.reg_window\[147\] vssd1 vssd1 vccd1 vccd1 net2012 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout873_X net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold681 final_design.cpu.reg_window\[573\] vssd1 vssd1 vccd1 vccd1 net2023 sky130_fd_sc_hd__dlygate4sd3_1
Xhold692 final_design.cpu.reg_window\[359\] vssd1 vssd1 vccd1 vccd1 net2034 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09734__A1 _04124_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11031_ _05729_ _05747_ _05752_ _05732_ vssd1 vssd1 vccd1 vccd1 _05755_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_40_1727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11675__C net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11541__A1 net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06643__S1 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12982_ net1313 _00213_ net1155 vssd1 vssd1 vccd1 vccd1 final_design.CPU_instr_adr\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input12_A DAT_I[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_2400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11933_ _06134_ net276 net408 net2084 vssd1 vssd1 vccd1 vccd1 _00668_ sky130_fd_sc_hd__a22o_1
XANTENNA__11691__B net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07233__Y _02184_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11864_ net2425 net518 _06242_ net432 vssd1 vssd1 vccd1 vccd1 _00611_ sky130_fd_sc_hd__a22o_1
XFILLER_0_19_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08058__A net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13603_ clknet_leaf_0_clk _00834_ net1061 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[591\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_32_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10815_ _05547_ _05548_ _05529_ vssd1 vssd1 vccd1 vccd1 _05549_ sky130_fd_sc_hd__o21bai_1
X_11795_ net2476 net413 _06234_ net428 vssd1 vssd1 vccd1 vccd1 _00550_ sky130_fd_sc_hd__a22o_1
XANTENNA__11911__S net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09896__S1 net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13440__CLK clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13534_ clknet_leaf_12_clk _00765_ net1088 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[522\]
+ sky130_fd_sc_hd__dfrtp_1
X_10746_ net727 _04509_ net253 _04990_ vssd1 vssd1 vccd1 vccd1 _05483_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_40_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09670__B1 net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13465_ clknet_leaf_56_clk _00696_ net1146 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[453\]
+ sky130_fd_sc_hd__dfrtp_1
X_10677_ net38 _05406_ _05414_ _05417_ vssd1 vssd1 vccd1 vccd1 _05418_ sky130_fd_sc_hd__nand4_1
XTAP_TAPCELL_ROW_77_2827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_2204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_2838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12557__B1 net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_2849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12416_ net199 net553 net500 net339 net1903 vssd1 vssd1 vccd1 vccd1 _01126_ sky130_fd_sc_hd__a32o_1
XANTENNA__12021__A2 net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13396_ clknet_leaf_9_clk _00627_ net1104 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[384\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13590__CLK clknet_leaf_62_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12347_ net2343 net361 net348 _05981_ vssd1 vssd1 vccd1 vccd1 _01059_ sky130_fd_sc_hd__a22o_1
XFILLER_0_51_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09176__X _04095_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12278_ net561 _06208_ net504 net368 net1908 vssd1 vssd1 vccd1 vccd1 _00993_ sky130_fd_sc_hd__a32o_1
X_14017_ clknet_leaf_47_clk _01248_ net1199 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[1005\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09725__A1 net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11229_ _04766_ net652 net591 _05933_ vssd1 vssd1 vccd1 vccd1 _05934_ sky130_fd_sc_hd__o211a_2
XFILLER_0_4_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_1671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12088__A2 _06053_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06770_ final_design.data_from_mem\[23\] net969 _01719_ vssd1 vssd1 vccd1 vccd1 _01721_
+ sky130_fd_sc_hd__o21ai_1
XANTENNA_clkbuf_leaf_11_clk_X clknet_leaf_11_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14096__CLK clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08387__S1 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12189__S net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08440_ _03387_ _03389_ vssd1 vssd1 vccd1 vccd1 _03391_ sky130_fd_sc_hd__or2_2
XFILLER_0_59_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08371_ net597 _03321_ vssd1 vssd1 vccd1 vccd1 _03322_ sky130_fd_sc_hd__or2_1
XANTENNA__11599__A1 net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11821__S net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07322_ final_design.cpu.reg_window\[452\] final_design.cpu.reg_window\[484\] net902
+ vssd1 vssd1 vccd1 vccd1 _02273_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08464__B2 net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07898__S0 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13933__CLK clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07253_ _02200_ _02201_ _02202_ _02203_ net764 net785 vssd1 vssd1 vccd1 vccd1 _02204_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_61_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12548__B1 net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07184_ _02131_ _02132_ _02133_ _02134_ net764 net785 vssd1 vssd1 vccd1 vccd1 _02135_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__12012__A2 net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_1885 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11220__B1 _05924_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07746__S net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09716__A1 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout402 _06257_ vssd1 vssd1 vccd1 vccd1 net402 sky130_fd_sc_hd__buf_6
XANTENNA_fanout499_A net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout413 net415 vssd1 vssd1 vccd1 vccd1 net413 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_6_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout424 _05877_ vssd1 vssd1 vccd1 vccd1 net424 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_6_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout435 net436 vssd1 vssd1 vccd1 vccd1 net435 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11523__A1 net197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08924__C1 net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout446 _04088_ vssd1 vssd1 vccd1 vccd1 net446 sky130_fd_sc_hd__clkbuf_4
XANTENNA_input4_A DAT_I[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13313__CLK clknet_leaf_49_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout457 _03551_ vssd1 vssd1 vccd1 vccd1 net457 sky130_fd_sc_hd__buf_2
X_09825_ _04737_ _04740_ _04743_ net450 vssd1 vssd1 vccd1 vccd1 _04744_ sky130_fd_sc_hd__a22o_2
Xfanout468 net469 vssd1 vssd1 vccd1 vccd1 net468 sky130_fd_sc_hd__buf_1
XANTENNA__06625__S1 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout479 net480 vssd1 vssd1 vccd1 vccd1 net479 sky130_fd_sc_hd__buf_2
XANTENNA_fanout666_A net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout287_X net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12988__RESET_B net1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09756_ _03198_ _04674_ vssd1 vssd1 vccd1 vccd1 _04675_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_74_1801 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06886__A net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06968_ final_design.cpu.reg_window\[16\] final_design.cpu.reg_window\[48\] net926
+ vssd1 vssd1 vccd1 vccd1 _01919_ sky130_fd_sc_hd__mux2_1
XANTENNA__08577__S net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11287__B1 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08707_ _03656_ _03657_ vssd1 vssd1 vccd1 vccd1 _03658_ sky130_fd_sc_hd__and2b_1
XFILLER_0_74_1845 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12099__S net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09687_ net545 net544 net542 net541 net454 net464 vssd1 vssd1 vccd1 vccd1 _04606_
+ sky130_fd_sc_hd__mux4_1
X_06899_ net882 _01831_ _01837_ _01843_ _01849_ vssd1 vssd1 vccd1 vccd1 _01850_ sky130_fd_sc_hd__o32a_4
XANTENNA_fanout833_A net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout454_X net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1196_X net1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13463__CLK clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1889 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08638_ _03586_ _03588_ vssd1 vssd1 vccd1 vccd1 _03589_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout621_X net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08569_ net595 _03514_ _03516_ _02390_ vssd1 vssd1 vccd1 vccd1 _03520_ sky130_fd_sc_hd__o211a_2
XANTENNA_fanout719_X net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10600_ _05343_ _05344_ vssd1 vssd1 vccd1 vccd1 _05345_ sky130_fd_sc_hd__or2_1
XFILLER_0_37_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11580_ net589 _06016_ net636 vssd1 vssd1 vccd1 vccd1 _06146_ sky130_fd_sc_hd__and3_1
XFILLER_0_0_1805 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10531_ _05277_ _05278_ vssd1 vssd1 vccd1 vccd1 _05279_ sky130_fd_sc_hd__and2_1
XFILLER_0_64_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_1849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12539__B1 net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13250_ clknet_leaf_3_clk _00481_ net1067 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[238\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_17_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12003__A2 net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10462_ _02540_ net592 vssd1 vssd1 vccd1 vccd1 _05215_ sky130_fd_sc_hd__nor2_1
XFILLER_0_66_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_1805 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12201_ _06129_ net498 net376 net2161 vssd1 vssd1 vccd1 vccd1 _00919_ sky130_fd_sc_hd__a22o_1
XANTENNA__14116__Q final_design.reqhand.data_from_UART\[6\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_66_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13181_ clknet_leaf_2_clk _00412_ net1064 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[169\]
+ sky130_fd_sc_hd__dfrtp_1
X_10393_ net801 net1002 _05178_ net1029 net167 vssd1 vssd1 vccd1 vccd1 _00139_ sky130_fd_sc_hd__a32o_1
XANTENNA__06769__A1 final_design.data_from_mem\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07966__B1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12132_ net241 net2361 net385 vssd1 vssd1 vccd1 vccd1 _00853_ sky130_fd_sc_hd__mux2_1
XANTENNA__09437__A net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09707__A1 _04124_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12063_ _05865_ net566 net506 net393 net1988 vssd1 vssd1 vccd1 vccd1 _00788_ sky130_fd_sc_hd__a32o_1
XANTENNA__10317__A2 net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11514__A1 net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11014_ net86 net1045 net87 vssd1 vssd1 vccd1 vccd1 _05739_ sky130_fd_sc_hd__or3b_1
XANTENNA__09183__A2 net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout980 net981 vssd1 vssd1 vccd1 vccd1 net980 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11906__S net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout991 _01413_ vssd1 vssd1 vccd1 vccd1 net991 sky130_fd_sc_hd__clkbuf_2
XANTENNA__13806__CLK clknet_leaf_45_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09172__A _03635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09566__S0 net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12965_ clknet_leaf_32_clk _00203_ net1234 vssd1 vssd1 vccd1 vccd1 net124 sky130_fd_sc_hd__dfrtp_1
X_11916_ net182 net2031 net275 vssd1 vssd1 vccd1 vccd1 _00655_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_1863 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12490__A2 net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09891__B1 net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12896_ clknet_leaf_25_clk _00134_ net1152 vssd1 vssd1 vccd1 vccd1 final_design.data_from_mem\[30\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_73_1388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13956__CLK clknet_leaf_54_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11847_ _06097_ net282 net518 final_design.cpu.reg_window\[354\] vssd1 vssd1 vccd1
+ vccd1 _00597_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_16_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_1749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_16_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11778_ net2532 net413 net280 _05905_ vssd1 vssd1 vccd1 vccd1 _00537_ sky130_fd_sc_hd__a22o_1
XFILLER_0_51_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13517_ clknet_leaf_44_clk _00748_ net1201 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[505\]
+ sky130_fd_sc_hd__dfrtp_1
X_10729_ _05465_ _05466_ _05446_ vssd1 vssd1 vccd1 vccd1 _05467_ sky130_fd_sc_hd__o21a_1
XFILLER_0_43_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07654__C1 _01566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12980__CLK clknet_leaf_19_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13448_ clknet_leaf_35_clk _00679_ net1240 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[436\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload12 clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 clkload12/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload23 clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 clkload23/Y sky130_fd_sc_hd__clkinv_16
XFILLER_0_49_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload34 clknet_leaf_43_clk vssd1 vssd1 vccd1 vccd1 clkload34/Y sky130_fd_sc_hd__inv_6
Xclkload45 clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 clkload45/Y sky130_fd_sc_hd__inv_12
XANTENNA__11202__B1 net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13379_ clknet_leaf_1_clk _00610_ net1074 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[367\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_1435 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13336__CLK clknet_leaf_63_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_53_clk_A clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11596__B net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09347__A net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09159__C1 _02423_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07940_ final_design.cpu.reg_window\[534\] final_design.cpu.reg_window\[566\] net839
+ vssd1 vssd1 vccd1 vccd1 _02891_ sky130_fd_sc_hd__mux2_1
XANTENNA__08057__S0 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07871_ _02818_ _02819_ _02820_ _02821_ net687 net705 vssd1 vssd1 vccd1 vccd1 _02822_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__06607__S1 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11816__S net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09610_ net727 _04513_ _04527_ vssd1 vssd1 vccd1 vccd1 _04529_ sky130_fd_sc_hd__or3_4
XANTENNA__13486__CLK clknet_leaf_43_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06822_ final_design.cpu.reg_window\[789\] final_design.cpu.reg_window\[821\] net938
+ vssd1 vssd1 vccd1 vccd1 _01773_ sky130_fd_sc_hd__mux2_1
XANTENNA__08397__S net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12060__X _06263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09082__A net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_3020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09541_ net481 _04459_ vssd1 vssd1 vccd1 vccd1 _04460_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_82_3031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06753_ net756 _01697_ net747 vssd1 vssd1 vccd1 vccd1 _01704_ sky130_fd_sc_hd__o21a_1
XANTENNA__11808__A2 net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_3042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_82_3053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09472_ _02609_ _04167_ _04170_ vssd1 vssd1 vccd1 vccd1 _04391_ sky130_fd_sc_hd__nand3_1
X_06684_ final_design.cpu.reg_window\[473\] final_design.cpu.reg_window\[505\] net933
+ vssd1 vssd1 vccd1 vccd1 _01635_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12481__A2 net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08423_ final_design.cpu.reg_window\[773\] final_design.cpu.reg_window\[805\] net843
+ vssd1 vssd1 vccd1 vccd1 _03374_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout247_A _04986_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06791__S0 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08354_ final_design.cpu.reg_window\[199\] final_design.cpu.reg_window\[231\] net809
+ vssd1 vssd1 vccd1 vccd1 _03305_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_28_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_24_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07330__A net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07305_ final_design.cpu.reg_window\[773\] final_design.cpu.reg_window\[805\] net923
+ vssd1 vssd1 vccd1 vccd1 _02256_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_43_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload6 clknet_leaf_64_clk vssd1 vssd1 vccd1 vccd1 clkload6/Y sky130_fd_sc_hd__inv_6
X_08285_ final_design.cpu.reg_window\[393\] final_design.cpu.reg_window\[425\] net810
+ vssd1 vssd1 vccd1 vccd1 _03236_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_43_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout414_A net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14111__CLK clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07236_ _02185_ _02186_ vssd1 vssd1 vccd1 vccd1 _02187_ sky130_fd_sc_hd__nand2_1
XFILLER_0_61_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09398__C1 _04109_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12382__S net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09937__B2 _04309_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07167_ _02114_ _02115_ _02116_ _02117_ net766 net786 vssd1 vssd1 vccd1 vccd1 _02118_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_67_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07099__S1 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07098_ final_design.cpu.reg_window\[908\] final_design.cpu.reg_window\[940\] net898
+ vssd1 vssd1 vccd1 vccd1 _02049_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout783_A net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07048__Y _01999_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout210 net211 vssd1 vssd1 vccd1 vccd1 net210 sky130_fd_sc_hd__clkbuf_2
XANTENNA__13829__CLK clknet_leaf_51_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1208 net1209 vssd1 vssd1 vccd1 vccd1 net1208 sky130_fd_sc_hd__clkbuf_4
Xfanout1219 net1221 vssd1 vssd1 vccd1 vccd1 net1219 sky130_fd_sc_hd__clkbuf_4
Xfanout221 _05921_ vssd1 vssd1 vccd1 vccd1 net221 sky130_fd_sc_hd__buf_2
Xfanout232 _05858_ vssd1 vssd1 vccd1 vccd1 net232 sky130_fd_sc_hd__clkbuf_4
Xfanout243 net244 vssd1 vssd1 vccd1 vccd1 net243 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout571_X net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout254 net255 vssd1 vssd1 vccd1 vccd1 net254 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout950_A net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07176__A1 net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout265 net267 vssd1 vssd1 vccd1 vccd1 net265 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout669_X net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout276 net277 vssd1 vssd1 vccd1 vccd1 net276 sky130_fd_sc_hd__clkbuf_4
Xfanout287 _06228_ vssd1 vssd1 vccd1 vccd1 net287 sky130_fd_sc_hd__buf_2
X_09808_ net594 _04220_ vssd1 vssd1 vccd1 vccd1 _04727_ sky130_fd_sc_hd__or2_2
Xfanout298 net299 vssd1 vssd1 vccd1 vccd1 net298 sky130_fd_sc_hd__buf_4
XANTENNA__12853__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09739_ net69 net70 _04182_ vssd1 vssd1 vccd1 vccd1 _04658_ sky130_fd_sc_hd__nand3_1
XANTENNA__13979__CLK clknet_leaf_65_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout836_X net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_3_4_0_clk_X clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12750_ _06351_ _06384_ vssd1 vssd1 vccd1 vccd1 _06388_ sky130_fd_sc_hd__xor2_1
XFILLER_0_69_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12472__A2 net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11701_ net205 net626 vssd1 vssd1 vccd1 vccd1 _06209_ sky130_fd_sc_hd__and2_1
XFILLER_0_55_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12681_ final_design.VGA_data_control.ready_data\[28\] net1021 net977 final_design.data_from_mem\[28\]
+ vssd1 vssd1 vccd1 vccd1 _06328_ sky130_fd_sc_hd__a22o_1
XANTENNA__11680__B1 net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07884__C1 _01815_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13209__CLK clknet_leaf_57_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11461__S net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11632_ net434 net578 _06173_ net300 net1525 vssd1 vssd1 vccd1 vccd1 _00448_ sky130_fd_sc_hd__a32o_1
XANTENNA__08523__S1 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11563_ net425 net560 _06137_ net302 net1887 vssd1 vssd1 vccd1 vccd1 _00415_ sky130_fd_sc_hd__a32o_1
XFILLER_0_80_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13302_ clknet_leaf_59_clk _00533_ net1138 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[290\]
+ sky130_fd_sc_hd__dfrtp_1
X_10514_ net61 _05250_ _05260_ _05262_ vssd1 vssd1 vccd1 vccd1 _05263_ sky130_fd_sc_hd__and4_1
XANTENNA__13359__CLK clknet_leaf_41_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11494_ net179 net640 vssd1 vssd1 vccd1 vccd1 _06115_ sky130_fd_sc_hd__and2_1
XANTENNA__11697__A net209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13233_ clknet_leaf_34_clk _00464_ net1242 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[221\]
+ sky130_fd_sc_hd__dfrtp_1
X_10445_ net1607 net1027 _05206_ net245 vssd1 vssd1 vccd1 vccd1 _00163_ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13164_ clknet_leaf_47_clk _00395_ net1203 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[152\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10376_ net19 net1024 net1006 final_design.data_from_mem\[25\] vssd1 vssd1 vccd1
+ vccd1 _00129_ sky130_fd_sc_hd__o22a_1
XFILLER_0_20_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output166_A net166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12115_ net1756 net198 net390 vssd1 vssd1 vccd1 vccd1 _00839_ sky130_fd_sc_hd__mux2_1
X_13095_ clknet_leaf_62_clk _00326_ net1124 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[83\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09156__A2 net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09454__X _04373_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12046_ net2039 net200 net397 vssd1 vssd1 vccd1 vccd1 _00774_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_1439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09106__S net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09539__S0 net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13997_ clknet_leaf_44_clk _01228_ net1201 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[985\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1873 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12948_ clknet_leaf_29_clk _00186_ net1194 vssd1 vssd1 vccd1 vccd1 net105 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_34_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12879_ clknet_leaf_21_clk _00117_ net1158 vssd1 vssd1 vccd1 vccd1 final_design.data_from_mem\[13\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__14134__CLK clknet_leaf_18_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1579 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_904 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07150__A net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08070_ _03015_ _03020_ net714 vssd1 vssd1 vccd1 vccd1 _03021_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07021_ final_design.cpu.reg_window\[270\] final_design.cpu.reg_window\[302\] net906
+ vssd1 vssd1 vccd1 vccd1 _01972_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_1833 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11726__A1 net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06602__B1 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08972_ net258 _03909_ net1016 vssd1 vssd1 vccd1 vccd1 _03910_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10016__A net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12876__CLK clknet_leaf_19_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09805__A net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07923_ _02870_ _02871_ _02872_ _02873_ net680 net700 vssd1 vssd1 vccd1 vccd1 _02874_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_32_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold18 net132 vssd1 vssd1 vccd1 vccd1 net1360 sky130_fd_sc_hd__dlygate4sd3_1
Xhold29 net105 vssd1 vssd1 vccd1 vccd1 net1371 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_32_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout197_A net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07854_ _01504_ _01822_ net616 vssd1 vssd1 vccd1 vccd1 _02805_ sky130_fd_sc_hd__a21o_1
XANTENNA__08450__S0 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07253__S1 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06805_ _01499_ _01503_ _01754_ vssd1 vssd1 vccd1 vccd1 _01756_ sky130_fd_sc_hd__or3b_2
X_07785_ net604 _02731_ _02707_ net552 vssd1 vssd1 vccd1 vccd1 _02736_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout364_A net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09304__C1 _02503_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09524_ net471 _04107_ _04240_ vssd1 vssd1 vccd1 vccd1 _04443_ sky130_fd_sc_hd__and3_1
X_06736_ final_design.reqhand.instruction\[24\] final_design.data_from_mem\[24\] net971
+ vssd1 vssd1 vccd1 vccd1 _01687_ sky130_fd_sc_hd__mux2_4
XANTENNA__08658__B2 _02545_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1214 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1383 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10465__A1 net68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11662__B1 net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09455_ net472 _04299_ vssd1 vssd1 vccd1 vccd1 _04374_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_49_1888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12377__S net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06667_ _01614_ _01615_ _01616_ _01617_ net775 net793 vssd1 vssd1 vccd1 vccd1 _01618_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_26_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07979__B _02929_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout629_A _06192_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06764__S0 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11134__X _05849_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08406_ net597 _03352_ _03328_ _02239_ vssd1 vssd1 vccd1 vccd1 _03357_ sky130_fd_sc_hd__o211a_1
X_09386_ _04303_ _04304_ net476 vssd1 vssd1 vccd1 vccd1 _04305_ sky130_fd_sc_hd__mux2_1
X_06598_ final_design.cpu.reg_window\[284\] final_design.cpu.reg_window\[316\] net946
+ vssd1 vssd1 vccd1 vccd1 _01549_ sky130_fd_sc_hd__mux2_1
XANTENNA__07881__A2 _02830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13501__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08337_ _02186_ net610 vssd1 vssd1 vccd1 vccd1 _03288_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout417_X net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07094__B1 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08268_ final_design.cpu.reg_window\[650\] final_design.cpu.reg_window\[682\] net815
+ vssd1 vssd1 vccd1 vccd1 _03219_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07219_ net757 _02169_ vssd1 vssd1 vccd1 vccd1 _02170_ sky130_fd_sc_hd__or2_1
X_08199_ final_design.cpu.reg_window\[974\] final_design.cpu.reg_window\[1006\] net816
+ vssd1 vssd1 vccd1 vccd1 _03150_ sky130_fd_sc_hd__mux2_1
XANTENNA__13651__CLK clknet_leaf_38_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10230_ final_design.uart.BAUD_counter\[9\] final_design.uart.BAUD_counter\[10\]
+ _05103_ final_design.uart.BAUD_counter\[11\] vssd1 vssd1 vccd1 vccd1 _05107_ sky130_fd_sc_hd__a31o_1
XFILLER_0_43_1917 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08043__C1 _01850_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06819__S1 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout786_X net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11193__A2 net251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10161_ final_design.VGA_data_control.VGA_request_address\[0\] _05054_ _05041_ vssd1
+ vssd1 vccd1 vccd1 _05056_ sky130_fd_sc_hd__a21oi_1
Xfanout1005 _05172_ vssd1 vssd1 vccd1 vccd1 net1005 sky130_fd_sc_hd__buf_4
XANTENNA__07934__S net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1016 net1017 vssd1 vssd1 vccd1 vccd1 net1016 sky130_fd_sc_hd__buf_2
XANTENNA__09138__A2 net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1027 net1028 vssd1 vssd1 vccd1 vccd1 net1027 sky130_fd_sc_hd__buf_2
XANTENNA__14007__CLK clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10092_ final_design.VGA_data_control.VGA_request_address\[1\] final_design.VGA_data_control.VGA_request_address\[0\]
+ vssd1 vssd1 vccd1 vccd1 _05008_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout953_X net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1038 _01410_ vssd1 vssd1 vccd1 vccd1 net1038 sky130_fd_sc_hd__clkbuf_4
X_14221__1279 vssd1 vssd1 vccd1 vccd1 _14221__1279/HI net1279 sky130_fd_sc_hd__conb_1
Xfanout1049 final_design.VGA_data_control.h_count\[2\] vssd1 vssd1 vccd1 vccd1 net1049
+ sky130_fd_sc_hd__clkbuf_4
X_13920_ clknet_leaf_10_clk _01151_ net1097 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[908\]
+ sky130_fd_sc_hd__dfrtp_1
X_13851_ clknet_leaf_65_clk _01082_ net1073 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[839\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13031__CLK clknet_leaf_62_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14157__CLK clknet_leaf_18_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12802_ net1392 vssd1 vssd1 vccd1 vccd1 _00243_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_2_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13782_ clknet_leaf_58_clk _01013_ net1125 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[770\]
+ sky130_fd_sc_hd__dfrtp_1
X_10994_ _05718_ _05719_ _05698_ vssd1 vssd1 vccd1 vccd1 _05720_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_2_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09846__B1 net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12733_ _06364_ _06367_ vssd1 vssd1 vccd1 vccd1 _06374_ sky130_fd_sc_hd__nand2_1
XFILLER_0_6_1833 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10017__D_N _03617_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12664_ _06319_ net1527 net979 vssd1 vssd1 vccd1 vccd1 _01334_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_1877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13181__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_2277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11615_ net224 net631 vssd1 vssd1 vccd1 vccd1 _06165_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_61_2288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_2299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12595_ net2244 net997 net983 final_design.data_from_mem\[13\] vssd1 vssd1 vccd1
+ vccd1 _01288_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09449__X _04368_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11546_ net563 net240 net634 vssd1 vssd1 vccd1 vccd1 _06129_ sky130_fd_sc_hd__and3_1
XFILLER_0_68_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07624__A2 _02570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_929 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09168__Y _04087_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11477_ net199 net2467 net307 vssd1 vssd1 vccd1 vccd1 _00358_ sky130_fd_sc_hd__mux2_1
XANTENNA__11708__A1 net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13216_ clknet_leaf_11_clk _00447_ net1086 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[204\]
+ sky130_fd_sc_hd__dfrtp_1
X_10428_ net1453 net1028 _05197_ net245 vssd1 vssd1 vccd1 vccd1 _00155_ sky130_fd_sc_hd__a22o_1
XANTENNA__09377__A2 _04223_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14196_ net1254 vssd1 vssd1 vccd1 vccd1 gpio_oeb[8] sky130_fd_sc_hd__buf_2
XANTENNA__12899__CLK clknet_leaf_62_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08585__B1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13147_ clknet_leaf_66_clk _00378_ net1063 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[135\]
+ sky130_fd_sc_hd__dfrtp_1
X_10359_ net32 net1025 net1008 final_design.data_from_mem\[8\] vssd1 vssd1 vccd1 vccd1
+ _00112_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_29_Left_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13078_ clknet_leaf_60_clk _00309_ net1139 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[66\]
+ sky130_fd_sc_hd__dfrtp_1
X_12029_ net1637 net241 net397 vssd1 vssd1 vccd1 vccd1 _00757_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10695__A1 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11892__A0 net244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07570_ net711 _02520_ vssd1 vssd1 vccd1 vccd1 _02521_ sky130_fd_sc_hd__nor2_1
XFILLER_0_53_1501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09837__B1 _04341_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06521_ final_design.data_from_mem\[0\] final_design.data_from_mem\[1\] net1039 net994
+ net991 vssd1 vssd1 vccd1 vccd1 _01472_ sky130_fd_sc_hd__a2111oi_1
XANTENNA__10447__A1 net149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13524__CLK clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11644__B1 net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10447__B2 net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_38_Left_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12197__S net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06746__S0 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09240_ _02934_ _03587_ _02932_ vssd1 vssd1 vccd1 vccd1 _04159_ sky130_fd_sc_hd__a21oi_1
X_06452_ net1053 net1057 vssd1 vssd1 vccd1 vccd1 _01406_ sky130_fd_sc_hd__nor2_1
XFILLER_0_69_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09171_ _03628_ _03650_ vssd1 vssd1 vccd1 vccd1 _04090_ sky130_fd_sc_hd__or2_1
XFILLER_0_51_1291 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13674__CLK clknet_leaf_60_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08122_ final_design.cpu.reg_window\[461\] final_design.cpu.reg_window\[493\] net851
+ vssd1 vssd1 vccd1 vccd1 _03073_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_1297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08053_ final_design.cpu.reg_window\[82\] final_design.cpu.reg_window\[114\] net844
+ vssd1 vssd1 vccd1 vccd1 _03004_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07004_ final_design.cpu.reg_window\[847\] final_design.cpu.reg_window\[879\] net900
+ vssd1 vssd1 vccd1 vccd1 _01955_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_38_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_47_Left_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12372__A1 net221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1021_A _06298_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1119_A net1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08955_ final_design.CPU_instr_adr\[20\] net1016 _03891_ _03894_ vssd1 vssd1 vccd1
+ vccd1 _00231_ sky130_fd_sc_hd__a22o_1
XANTENNA__11784__B net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout481_A net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13054__CLK clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07906_ final_design.cpu.reg_window\[727\] final_design.cpu.reg_window\[759\] net849
+ vssd1 vssd1 vccd1 vccd1 _02857_ sky130_fd_sc_hd__mux2_1
X_08886_ _01600_ _01601_ _02472_ vssd1 vssd1 vccd1 vccd1 _03833_ sky130_fd_sc_hd__nand3_1
XANTENNA__08879__A1 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07837_ final_design.cpu.reg_window\[981\] final_design.cpu.reg_window\[1013\] net858
+ vssd1 vssd1 vccd1 vccd1 _02788_ sky130_fd_sc_hd__mux2_1
XANTENNA__07551__A1 net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout746_A _01438_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout367_X net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07768_ net711 _02712_ net723 vssd1 vssd1 vccd1 vccd1 _02719_ sky130_fd_sc_hd__o21a_1
XANTENNA__12427__A2 net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09507_ _03590_ _04143_ _04157_ vssd1 vssd1 vccd1 vccd1 _04426_ sky130_fd_sc_hd__or3_1
XFILLER_0_67_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06719_ final_design.cpu.reg_window\[280\] final_design.cpu.reg_window\[312\] net944
+ vssd1 vssd1 vccd1 vccd1 _01670_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout913_A net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07303__A1 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07699_ final_design.cpu.reg_window\[91\] final_design.cpu.reg_window\[123\] net862
+ vssd1 vssd1 vccd1 vccd1 _02650_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09438_ net82 _04190_ vssd1 vssd1 vccd1 vccd1 _04357_ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09369_ _04194_ _04287_ vssd1 vssd1 vccd1 vccd1 _04288_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout701_X net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13131__RESET_B net1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11400_ net738 _03803_ _06083_ vssd1 vssd1 vccd1 vccd1 _06084_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_30_1375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12380_ net1654 net222 net269 vssd1 vssd1 vccd1 vccd1 _01091_ sky130_fd_sc_hd__mux2_1
XANTENNA__09461__D1 net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_10_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_1596 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11331_ net656 _06022_ _06023_ net590 vssd1 vssd1 vccd1 vccd1 _06024_ sky130_fd_sc_hd__o211a_2
XFILLER_0_22_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14050_ clknet_leaf_16_clk _00011_ net1093 vssd1 vssd1 vccd1 vccd1 final_design.uart.BAUD_counter\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_11262_ _02000_ net641 _05962_ net658 vssd1 vssd1 vccd1 vccd1 _05963_ sky130_fd_sc_hd__a211o_1
X_13001_ net1332 _00232_ net1196 vssd1 vssd1 vccd1 vccd1 final_design.CPU_instr_adr\[21\]
+ sky130_fd_sc_hd__dfrtp_2
X_10213_ net2518 _05094_ _05096_ vssd1 vssd1 vccd1 vccd1 _00032_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_73_2682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11193_ final_design.data_from_mem\[6\] net251 _05855_ _05901_ vssd1 vssd1 vccd1
+ vccd1 _05902_ sky130_fd_sc_hd__o211a_1
XANTENNA__10374__B1 net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_2693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07664__S net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input42_A mem_adr_start[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10144_ _01389_ _05044_ _05042_ vssd1 vssd1 vccd1 vccd1 _05045_ sky130_fd_sc_hd__o21ai_1
XANTENNA__12115__A1 net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10075_ net2553 _01372_ wb_manage.curr_state\[0\] _04992_ vssd1 vssd1 vccd1 vccd1
+ _00005_ sky130_fd_sc_hd__a22o_1
XANTENNA__08414__S0 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13547__CLK clknet_leaf_52_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13903_ clknet_leaf_42_clk _01134_ net1223 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[891\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11874__B1 net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13972__RESET_B net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09451__Y _04370_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13834_ clknet_leaf_59_clk _01065_ net1143 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[822\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08495__S net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_2486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13765_ clknet_leaf_50_clk _00996_ net1182 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[753\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11626__B1 net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10977_ final_design.CPU_instr_adr\[25\] _05703_ net1055 vssd1 vssd1 vccd1 vccd1
+ _05704_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06728__S0 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13697__CLK clknet_leaf_47_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11215__A net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12716_ final_design.VGA_data_control.v_count\[3\] _06348_ _06350_ vssd1 vssd1 vccd1
+ vccd1 _06357_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_73_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13696_ clknet_leaf_11_clk _00927_ net1086 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[684\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_1516 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12647_ final_design.VGA_data_control.ready_data\[11\] net1019 net974 final_design.data_from_mem\[11\]
+ vssd1 vssd1 vccd1 vccd1 _06311_ sky130_fd_sc_hd__a22o_1
XFILLER_0_26_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06743__S net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12578_ net1052 net35 vssd1 vssd1 vccd1 vccd1 _06294_ sky130_fd_sc_hd__and2_1
XFILLER_0_80_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11529_ net1603 net188 net523 vssd1 vssd1 vccd1 vccd1 _00396_ sky130_fd_sc_hd__mux2_1
Xhold307 final_design.cpu.reg_window\[962\] vssd1 vssd1 vccd1 vccd1 net1649 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1901 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold318 final_design.cpu.reg_window\[682\] vssd1 vssd1 vccd1 vccd1 net1660 sky130_fd_sc_hd__dlygate4sd3_1
X_14248_ net1302 vssd1 vssd1 vccd1 vccd1 gpio_out[26] sky130_fd_sc_hd__buf_2
XANTENNA__12854__RESET_B net1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold329 final_design.cpu.reg_window\[524\] vssd1 vssd1 vccd1 vccd1 net1671 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_1825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13077__CLK clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14179_ clknet_leaf_22_clk _01353_ net1164 vssd1 vssd1 vccd1 vccd1 final_design.VGA_adr\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10365__B1 net1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08530__Y _03481_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06979__A net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout809 net829 vssd1 vssd1 vccd1 vccd1 net809 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_0_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09770__A2 net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12782__13_A clknet_leaf_28_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08740_ final_design.CPU_instr_adr\[10\] _02128_ vssd1 vssd1 vccd1 vccd1 _03691_
+ sky130_fd_sc_hd__nor2_1
Xhold1007 final_design.cpu.reg_window\[95\] vssd1 vssd1 vccd1 vccd1 net2349 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1018 final_design.cpu.reg_window\[502\] vssd1 vssd1 vccd1 vccd1 net2360 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1029 final_design.cpu.reg_window\[96\] vssd1 vssd1 vccd1 vccd1 net2371 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_75_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08671_ _01568_ _01598_ _01628_ _01659_ vssd1 vssd1 vccd1 vccd1 _03622_ sky130_fd_sc_hd__or4_1
XANTENNA__11824__S net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07622_ net616 _02570_ _02571_ _01535_ vssd1 vssd1 vccd1 vccd1 _02573_ sky130_fd_sc_hd__a211oi_2
XANTENNA__12914__CLK clknet_leaf_28_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12409__A2 net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07553_ _01477_ _01497_ _01502_ vssd1 vssd1 vccd1 vccd1 _02504_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_18_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06504_ net1041 net993 net990 _01374_ vssd1 vssd1 vccd1 vccd1 _01455_ sky130_fd_sc_hd__a31o_1
XANTENNA__12290__B1 net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09381__S1 net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07484_ _02270_ _02434_ vssd1 vssd1 vccd1 vccd1 _02435_ sky130_fd_sc_hd__nand2_1
XFILLER_0_33_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09223_ _03199_ _03229_ _04136_ _04141_ vssd1 vssd1 vccd1 vccd1 _04142_ sky130_fd_sc_hd__a31o_1
X_06435_ final_design.VGA_data_control.VGA_request_address\[0\] vssd1 vssd1 vccd1
+ vccd1 _01390_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout327_A _06284_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14220__1278 vssd1 vssd1 vccd1 vccd1 _14220__1278/HI net1278 sky130_fd_sc_hd__conb_1
XANTENNA_fanout1069_A net1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07049__B1 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09154_ net497 net484 vssd1 vssd1 vccd1 vccd1 _04073_ sky130_fd_sc_hd__nor2_1
X_08105_ final_design.cpu.reg_window\[972\] final_design.cpu.reg_window\[1004\] net816
+ vssd1 vssd1 vccd1 vccd1 _03056_ sky130_fd_sc_hd__mux2_1
XANTENNA__09994__C1 net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12593__B2 final_design.data_from_mem\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09085_ _02435_ net622 _04005_ net254 vssd1 vssd1 vccd1 vccd1 _04010_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout1236_A net1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08153__B net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08036_ final_design.cpu.reg_window\[595\] final_design.cpu.reg_window\[627\] net822
+ vssd1 vssd1 vccd1 vccd1 _02987_ sky130_fd_sc_hd__mux2_1
Xinput90 memory_size[2] vssd1 vssd1 vccd1 vccd1 net90 sky130_fd_sc_hd__clkbuf_2
Xhold830 final_design.cpu.reg_window\[936\] vssd1 vssd1 vccd1 vccd1 net2172 sky130_fd_sc_hd__dlygate4sd3_1
Xhold841 final_design.cpu.reg_window\[1009\] vssd1 vssd1 vccd1 vccd1 net2183 sky130_fd_sc_hd__dlygate4sd3_1
Xhold852 final_design.cpu.reg_window\[167\] vssd1 vssd1 vccd1 vccd1 net2194 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08549__B1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout696_A net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14235__1289 vssd1 vssd1 vccd1 vccd1 _14235__1289/HI net1289 sky130_fd_sc_hd__conb_1
XFILLER_0_64_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12390__S net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold863 final_design.cpu.reg_window\[863\] vssd1 vssd1 vccd1 vccd1 net2205 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10356__B1 _05170_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold874 final_design.cpu.reg_window\[1018\] vssd1 vssd1 vccd1 vccd1 net2216 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1024_X net1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold885 final_design.cpu.reg_window\[348\] vssd1 vssd1 vccd1 vccd1 net2227 sky130_fd_sc_hd__dlygate4sd3_1
Xhold896 final_design.cpu.reg_window\[265\] vssd1 vssd1 vccd1 vccd1 net2238 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09761__A2 _04157_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09987_ _04654_ _04656_ _04905_ vssd1 vssd1 vccd1 vccd1 _04906_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout863_A net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08938_ net257 _03878_ net1014 vssd1 vssd1 vccd1 vccd1 _03880_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11305__C1 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout651_X net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08869_ net624 _03815_ vssd1 vssd1 vccd1 vccd1 _03818_ sky130_fd_sc_hd__nor2_1
XANTENNA__07524__A1 _01567_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout749_X net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11320__A2 net235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10900_ net82 net1046 vssd1 vssd1 vccd1 vccd1 _05630_ sky130_fd_sc_hd__nand2_1
XFILLER_0_73_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11880_ _06114_ net292 net519 net2204 vssd1 vssd1 vccd1 vccd1 _00624_ sky130_fd_sc_hd__a22o_1
XANTENNA__11871__A3 net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10831_ _05543_ _05562_ _05563_ net1005 vssd1 vssd1 vccd1 vccd1 _05565_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_81_2962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13550_ clknet_leaf_44_clk _00781_ net1208 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[538\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_81_2973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10762_ _05477_ _05481_ _05498_ vssd1 vssd1 vccd1 vccd1 _05499_ sky130_fd_sc_hd__or3_1
XFILLER_0_66_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12281__B1 net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_2984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_11_Right_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12501_ _06163_ net346 net326 net1713 vssd1 vssd1 vccd1 vccd1 _01206_ sky130_fd_sc_hd__a22o_1
XFILLER_0_32_1459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13481_ clknet_leaf_36_clk _00712_ net1230 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[469\]
+ sky130_fd_sc_hd__dfrtp_1
X_10693_ net965 _05432_ vssd1 vssd1 vccd1 vccd1 _05433_ sky130_fd_sc_hd__nand2_1
XANTENNA__11322__X _06016_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12432_ net1868 net231 net335 vssd1 vssd1 vccd1 vccd1 _01139_ sky130_fd_sc_hd__mux2_1
XANTENNA__11689__B net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06563__S net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11387__A2 _06070_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12363_ _06091_ net347 vssd1 vssd1 vccd1 vccd1 _06278_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_79_2891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_2110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_2121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14102_ clknet_leaf_14_clk _01299_ net1103 vssd1 vssd1 vccd1 vccd1 final_design.reqhand.instruction\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_75_2755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11314_ net643 _06007_ _06008_ vssd1 vssd1 vccd1 vccd1 _06009_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_56_2132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_2766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12294_ net577 _06224_ net510 net370 net1818 vssd1 vssd1 vccd1 vccd1 _01009_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_75_2777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_2619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14033_ clknet_leaf_34_clk _01264_ net1242 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[1021\]
+ sky130_fd_sc_hd__dfrtp_1
X_11245_ _05944_ _05945_ _05946_ _02064_ net655 vssd1 vssd1 vccd1 vccd1 _05948_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_20_Right_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07394__S net913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11176_ final_design.reqhand.data_from_UART\[4\] net251 vssd1 vssd1 vccd1 vccd1 _05887_
+ sky130_fd_sc_hd__nand2b_1
X_10127_ _01400_ _05000_ _05005_ vssd1 vssd1 vccd1 vccd1 final_design.v_out sky130_fd_sc_hd__or3b_1
XANTENNA__12937__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_2548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10058_ _04529_ _04530_ _04905_ _04975_ _04976_ vssd1 vssd1 vccd1 vccd1 _04977_ sky130_fd_sc_hd__a2111oi_1
XTAP_TAPCELL_ROW_69_2559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11847__B1 net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13817_ clknet_leaf_54_clk _01048_ net1177 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[805\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12272__B1 net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13748_ clknet_leaf_8_clk _00979_ net1153 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[736\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10784__A net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1346 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13679_ clknet_leaf_44_clk _00910_ net1208 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[667\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11232__X _05936_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06473__S net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07126__S0 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11378__A2 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08243__A2 _03192_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07677__S1 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold104 final_design.cpu.reg_window\[199\] vssd1 vssd1 vccd1 vccd1 net1446 sky130_fd_sc_hd__dlygate4sd3_1
Xhold115 net144 vssd1 vssd1 vccd1 vccd1 net1457 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09637__X _04556_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold126 final_design.VGA_data_control.ready_data\[31\] vssd1 vssd1 vccd1 vccd1 net1468
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09991__A2 net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold137 final_design.VGA_data_control.ready_data\[26\] vssd1 vssd1 vccd1 vccd1 net1479
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13712__CLK clknet_leaf_36_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold148 final_design.cpu.reg_window\[210\] vssd1 vssd1 vccd1 vccd1 net1490 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11819__S net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09910_ net90 net93 net94 vssd1 vssd1 vccd1 vccd1 _04829_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_65_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold159 final_design.cpu.reg_window\[215\] vssd1 vssd1 vccd1 vccd1 net1501 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout606 net607 vssd1 vssd1 vccd1 vccd1 net606 sky130_fd_sc_hd__buf_2
XANTENNA__10889__A1 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09841_ _04072_ _04753_ _04758_ _04759_ vssd1 vssd1 vccd1 vccd1 _04760_ sky130_fd_sc_hd__or4_1
Xfanout617 net618 vssd1 vssd1 vccd1 vccd1 net617 sky130_fd_sc_hd__clkbuf_2
XANTENNA__10889__B2 net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout628 net629 vssd1 vssd1 vccd1 vccd1 net628 sky130_fd_sc_hd__buf_4
XANTENNA_clkload14_A clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout639 _06093_ vssd1 vssd1 vccd1 vccd1 net639 sky130_fd_sc_hd__clkbuf_4
X_09772_ net474 _04645_ vssd1 vssd1 vccd1 vccd1 _04691_ sky130_fd_sc_hd__and2_1
XANTENNA__13862__CLK clknet_leaf_52_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06984_ _01931_ _01932_ _01933_ _01934_ net773 net784 vssd1 vssd1 vccd1 vccd1 _01935_
+ sky130_fd_sc_hd__mux4_1
X_08723_ final_design.CPU_instr_adr\[18\] _01881_ vssd1 vssd1 vccd1 vccd1 _03674_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_21_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout277_A net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11302__A2 net235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1415 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08654_ _01566_ _02604_ vssd1 vssd1 vccd1 vccd1 _03605_ sky130_fd_sc_hd__nor2_1
XANTENNA__10311__X final_design.pixel_data vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07605_ _02552_ _02553_ _02554_ _02555_ net687 net705 vssd1 vssd1 vccd1 vccd1 _02556_
+ sky130_fd_sc_hd__mux4_1
X_08585_ net709 _03529_ net722 vssd1 vssd1 vccd1 vccd1 _03536_ sky130_fd_sc_hd__o21a_1
XFILLER_0_77_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1186_A net1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07536_ _02483_ _02484_ _02485_ _02486_ net774 net792 vssd1 vssd1 vccd1 vccd1 _02487_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__11066__B2 _04042_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07467_ _02412_ _02417_ net750 vssd1 vssd1 vccd1 vccd1 _02418_ sky130_fd_sc_hd__mux2_1
XANTENNA__12385__S net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13242__CLK clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout232_X net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout611_A net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout709_A net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09206_ _04124_ vssd1 vssd1 vccd1 vccd1 _04125_ sky130_fd_sc_hd__inv_2
X_06418_ wb_manage.curr_state\[0\] vssd1 vssd1 vccd1 vccd1 _01373_ sky130_fd_sc_hd__inv_2
XANTENNA__12015__B1 net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07398_ _02345_ _02346_ _02347_ _02348_ net769 net782 vssd1 vssd1 vccd1 vccd1 _02349_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_31_1492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09137_ net496 _04054_ vssd1 vssd1 vccd1 vccd1 _04056_ sky130_fd_sc_hd__nand2_2
XANTENNA__11135__C_N net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09068_ _03786_ _03994_ vssd1 vssd1 vccd1 vccd1 _03995_ sky130_fd_sc_hd__nor2_1
XFILLER_0_66_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout980_A net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13392__CLK clknet_leaf_34_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12318__A1 net196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout699_X net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08019_ final_design.cpu.reg_window\[403\] final_design.cpu.reg_window\[435\] net821
+ vssd1 vssd1 vccd1 vccd1 _02970_ sky130_fd_sc_hd__mux2_1
XANTENNA__10329__B1 net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold660 final_design.cpu.reg_window\[422\] vssd1 vssd1 vccd1 vccd1 net2002 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold671 final_design.uart.working_data\[2\] vssd1 vssd1 vccd1 vccd1 net2013 sky130_fd_sc_hd__dlygate4sd3_1
X_11030_ _05693_ _05709_ vssd1 vssd1 vccd1 vccd1 _05754_ sky130_fd_sc_hd__nor2_1
Xhold682 final_design.cpu.reg_window\[77\] vssd1 vssd1 vccd1 vccd1 net2024 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09195__B1 _04113_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold693 final_design.cpu.reg_window\[464\] vssd1 vssd1 vccd1 vccd1 net2035 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_1905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08103__S net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06412__A net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11541__A2 net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12981_ clknet_leaf_20_clk _00212_ net1156 vssd1 vssd1 vccd1 vccd1 wb_manage.BUSY_O
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_77_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11932_ _06133_ net277 net408 net2484 vssd1 vssd1 vccd1 vccd1 _00667_ sky130_fd_sc_hd__a22o_1
XFILLER_0_58_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10501__B1 _04990_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_2401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11863_ net222 net554 vssd1 vssd1 vccd1 vccd1 _06242_ sky130_fd_sc_hd__and2_1
XFILLER_0_39_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10814_ net77 net1044 vssd1 vssd1 vccd1 vccd1 _05548_ sky130_fd_sc_hd__nor2_1
X_13602_ clknet_leaf_3_clk _00833_ net1067 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[590\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_36_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12254__B1 net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11794_ net648 net555 net199 vssd1 vssd1 vccd1 vccd1 _06234_ sky130_fd_sc_hd__and3_1
XANTENNA__10804__A1 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10745_ _05481_ _05482_ net1429 net1032 vssd1 vssd1 vccd1 vccd1 _00187_ sky130_fd_sc_hd__a2bb2o_1
X_13533_ clknet_leaf_2_clk _00764_ net1065 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[521\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_32_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07389__S net913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13464_ clknet_leaf_62_clk _00695_ net1119 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[452\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12006__B1 net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10676_ net961 _05416_ vssd1 vssd1 vccd1 vccd1 _05417_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_77_2828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13735__CLK clknet_leaf_63_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_2205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_2839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12415_ _06108_ net351 net339 net2119 vssd1 vssd1 vccd1 vccd1 _01125_ sky130_fd_sc_hd__a22o_1
X_13395_ clknet_leaf_40_clk _00626_ net1219 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[383\]
+ sky130_fd_sc_hd__dfrtp_1
X_12346_ net2346 net360 net342 _05973_ vssd1 vssd1 vccd1 vccd1 _01058_ sky130_fd_sc_hd__a22o_1
XFILLER_0_65_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12309__A1 net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12277_ net577 _06207_ net510 net370 net1615 vssd1 vssd1 vccd1 vccd1 _00992_ sky130_fd_sc_hd__a32o_1
XANTENNA__13885__CLK clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14016_ clknet_leaf_11_clk _01247_ net1097 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[1004\]
+ sky130_fd_sc_hd__dfrtp_1
X_11228_ net644 _05930_ _05931_ _05932_ net655 vssd1 vssd1 vccd1 vccd1 _05933_ sky130_fd_sc_hd__a221o_1
XANTENNA__09725__A2 net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08933__B1 _03655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09904__Y _04823_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11159_ final_design.reqhand.data_from_UART\[2\] net251 vssd1 vssd1 vccd1 vccd1 _05872_
+ sky130_fd_sc_hd__nand2b_1
XANTENNA__08948__S net1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12088__A3 net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12493__B1 net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13265__CLK clknet_leaf_34_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_67 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11048__A1 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12245__B1 net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08370_ _03308_ _03309_ _03320_ net874 vssd1 vssd1 vccd1 vccd1 _03321_ sky130_fd_sc_hd__a22oi_4
X_14234__1288 vssd1 vssd1 vccd1 vccd1 _14234__1288/HI net1288 sky130_fd_sc_hd__conb_1
XFILLER_0_74_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07321_ final_design.cpu.reg_window\[260\] final_design.cpu.reg_window\[292\] net903
+ vssd1 vssd1 vccd1 vccd1 _02272_ sky130_fd_sc_hd__mux2_1
XANTENNA__11599__A2 net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10032__C_N _04158_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_max_cap664_X net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07898__S1 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12260__A3 net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07299__S net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06475__A1 final_design.data_from_mem\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07252_ final_design.cpu.reg_window\[903\] final_design.cpu.reg_window\[935\] net892
+ vssd1 vssd1 vccd1 vccd1 _02203_ sky130_fd_sc_hd__mux2_1
XANTENNA__07672__B1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07183_ final_design.cpu.reg_window\[393\] final_design.cpu.reg_window\[425\] net891
+ vssd1 vssd1 vccd1 vccd1 _02134_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11220__A1 net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09808__A net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11771__A2 net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout403 _06257_ vssd1 vssd1 vccd1 vccd1 net403 sky130_fd_sc_hd__buf_2
Xfanout414 net415 vssd1 vssd1 vccd1 vccd1 net414 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_6_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout425 net426 vssd1 vssd1 vccd1 vccd1 net425 sky130_fd_sc_hd__clkbuf_4
Xfanout436 net437 vssd1 vssd1 vccd1 vccd1 net436 sky130_fd_sc_hd__buf_4
XANTENNA_fanout394_A net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout447 net449 vssd1 vssd1 vccd1 vccd1 net447 sky130_fd_sc_hd__buf_4
X_09824_ _03262_ _04742_ vssd1 vssd1 vccd1 vccd1 _04743_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout1101_A net1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout458 net459 vssd1 vssd1 vccd1 vccd1 net458 sky130_fd_sc_hd__clkbuf_4
Xfanout469 _03518_ vssd1 vssd1 vccd1 vccd1 net469 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07762__S net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14040__CLK clknet_leaf_15_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10888__A1_N net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06967_ final_design.cpu.reg_window\[80\] final_design.cpu.reg_window\[112\] net926
+ vssd1 vssd1 vccd1 vccd1 _01918_ sky130_fd_sc_hd__mux2_1
X_09755_ _03229_ _04503_ _03227_ vssd1 vssd1 vccd1 vccd1 _04674_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12079__A3 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout561_A net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout659_A _03649_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11287__A1 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13608__CLK clknet_leaf_40_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08706_ final_design.CPU_instr_adr\[30\] _01507_ vssd1 vssd1 vccd1 vccd1 _03657_
+ sky130_fd_sc_hd__or2_1
XANTENNA__12484__B1 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08688__C1 _02423_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09686_ net318 _04243_ vssd1 vssd1 vccd1 vccd1 _04605_ sky130_fd_sc_hd__nor2_1
X_06898_ net759 _01848_ net882 vssd1 vssd1 vccd1 vccd1 _01849_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_74_1857 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08637_ net613 _02961_ _02937_ _01938_ vssd1 vssd1 vccd1 vccd1 _03588_ sky130_fd_sc_hd__a211oi_2
XANTENNA_fanout826_A net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout447_X net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12957__RESET_B net1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12236__B1 net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08568_ net608 _03513_ _03515_ vssd1 vssd1 vccd1 vccd1 _03519_ sky130_fd_sc_hd__a21o_1
XFILLER_0_72_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13758__CLK clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07519_ _01661_ _02469_ vssd1 vssd1 vccd1 vccd1 _02470_ sky130_fd_sc_hd__nor2_1
XFILLER_0_65_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08499_ _03437_ _03438_ _03449_ net875 vssd1 vssd1 vccd1 vccd1 _03450_ sky130_fd_sc_hd__a22oi_4
XANTENNA__07112__C1 _01821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09652__A1 net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12251__A3 net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10530_ final_design.CPU_instr_adr\[4\] _05256_ vssd1 vssd1 vccd1 vccd1 _05278_ sky130_fd_sc_hd__or2_1
XFILLER_0_0_1817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_21_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12128__B net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10461_ net157 net1030 _05214_ net249 vssd1 vssd1 vccd1 vccd1 _00171_ sky130_fd_sc_hd__a22o_1
X_12200_ net565 _06128_ net505 net377 net1581 vssd1 vssd1 vccd1 vccd1 _00918_ sky130_fd_sc_hd__a32o_1
XANTENNA__11600__X _06156_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11211__A1 final_design.data_from_mem\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07937__S net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1817 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_3_0_0_clk_X clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13180_ clknet_leaf_3_clk _00411_ net1066 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[168\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09955__A2 _04087_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10392_ _04991_ _05176_ _04987_ vssd1 vssd1 vccd1 vccd1 _05178_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout983_X net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07966__A1 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11459__S net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12131_ net228 net2413 net385 vssd1 vssd1 vccd1 vccd1 _00852_ sky130_fd_sc_hd__mux2_1
XANTENNA__13138__CLK clknet_leaf_39_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12062_ net231 net2454 net393 vssd1 vssd1 vccd1 vccd1 _00787_ sky130_fd_sc_hd__mux2_1
Xhold490 final_design.cpu.reg_window\[460\] vssd1 vssd1 vccd1 vccd1 net1832 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11013_ _05736_ _05737_ _05719_ vssd1 vssd1 vccd1 vccd1 _05738_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_79_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout970 _01416_ vssd1 vssd1 vccd1 vccd1 net970 sky130_fd_sc_hd__clkbuf_8
Xfanout981 _06297_ vssd1 vssd1 vccd1 vccd1 net981 sky130_fd_sc_hd__clkbuf_2
Xfanout992 _01413_ vssd1 vssd1 vccd1 vccd1 net992 sky130_fd_sc_hd__clkbuf_2
XANTENNA__13288__CLK clknet_leaf_41_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11278__A1 final_design.data_from_mem\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09566__S1 net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09172__B net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12475__B1 net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12964_ clknet_leaf_32_clk _00202_ net1234 vssd1 vssd1 vccd1 vccd1 net122 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_1831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1190 final_design.cpu.reg_window\[294\] vssd1 vssd1 vccd1 vccd1 net2532 sky130_fd_sc_hd__dlygate4sd3_1
X_11915_ _06060_ _06248_ _06250_ net274 final_design.cpu.reg_window\[411\] vssd1 vssd1
+ vccd1 vccd1 _00654_ sky130_fd_sc_hd__a32o_1
X_12895_ clknet_leaf_21_clk _00133_ net1158 vssd1 vssd1 vccd1 vccd1 final_design.data_from_mem\[29\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_9_1875 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11922__S net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12227__B1 net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11846_ _06096_ net282 net518 net2141 vssd1 vssd1 vccd1 vccd1 _00596_ sky130_fd_sc_hd__a22o_1
XFILLER_0_51_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07329__S0 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11777_ net2490 net413 net283 _05898_ vssd1 vssd1 vccd1 vccd1 _00536_ sky130_fd_sc_hd__a22o_1
XANTENNA__12242__A3 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11223__A net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10728_ net73 net1043 vssd1 vssd1 vccd1 vccd1 _05466_ sky130_fd_sc_hd__nor2_1
X_13516_ clknet_leaf_46_clk _00747_ net1215 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[504\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_32_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10659_ net37 _05399_ vssd1 vssd1 vccd1 vccd1 _05401_ sky130_fd_sc_hd__or2_1
X_13447_ clknet_leaf_63_clk _00678_ net1122 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[435\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload13 clknet_leaf_12_clk vssd1 vssd1 vccd1 vccd1 clkload13/Y sky130_fd_sc_hd__clkinv_8
Xclkload24 clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 clkload24/Y sky130_fd_sc_hd__bufinv_16
Xclkload35 clknet_leaf_46_clk vssd1 vssd1 vccd1 vccd1 clkload35/Y sky130_fd_sc_hd__clkinvlp_4
XANTENNA__11202__A1 _04903_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09946__A2 _02325_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08603__C1 _02419_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13378_ clknet_leaf_10_clk _00609_ net1101 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[366\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_1414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09347__B net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12329_ _02328_ _05850_ _06260_ vssd1 vssd1 vccd1 vccd1 _06276_ sky130_fd_sc_hd__or3_1
XFILLER_0_45_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09159__B1 _01597_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07148__A net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14063__CLK clknet_leaf_15_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08057__S1 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07870_ final_design.cpu.reg_window\[916\] final_design.cpu.reg_window\[948\] net869
+ vssd1 vssd1 vccd1 vccd1 _02821_ sky130_fd_sc_hd__mux2_1
X_06821_ final_design.cpu.reg_window\[853\] final_design.cpu.reg_window\[885\] net938
+ vssd1 vssd1 vccd1 vccd1 _01772_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_30_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09540_ _04457_ _04458_ net477 vssd1 vssd1 vccd1 vccd1 _04459_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_82_3010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06752_ net763 _01702_ vssd1 vssd1 vccd1 vccd1 _01703_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_30_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_3021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12466__B1 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_3032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_3043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_3054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09471_ _04356_ _04358_ _04388_ vssd1 vssd1 vccd1 vccd1 _04390_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_56_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13900__CLK clknet_leaf_46_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06683_ final_design.cpu.reg_window\[281\] final_design.cpu.reg_window\[313\] net936
+ vssd1 vssd1 vccd1 vccd1 _01634_ sky130_fd_sc_hd__mux2_1
XANTENNA__09882__A1 net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11832__S net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08422_ final_design.cpu.reg_window\[837\] final_design.cpu.reg_window\[869\] net839
+ vssd1 vssd1 vccd1 vccd1 _03373_ sky130_fd_sc_hd__mux2_1
XANTENNA__12218__B1 net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09810__B _04087_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08353_ final_design.cpu.reg_window\[7\] final_design.cpu.reg_window\[39\] net806
+ vssd1 vssd1 vccd1 vccd1 _03304_ sky130_fd_sc_hd__mux2_1
XANTENNA__06791__S1 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12788__19 clknet_leaf_30_clk vssd1 vssd1 vccd1 vccd1 net1329 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_28_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12233__A3 net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07304_ final_design.cpu.reg_window\[837\] final_design.cpu.reg_window\[869\] net921
+ vssd1 vssd1 vccd1 vccd1 _02255_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_24_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08284_ final_design.cpu.reg_window\[457\] final_design.cpu.reg_window\[489\] net810
+ vssd1 vssd1 vccd1 vccd1 _03235_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_43_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload7 clknet_leaf_66_clk vssd1 vssd1 vccd1 vccd1 clkload7/Y sky130_fd_sc_hd__inv_12
XFILLER_0_27_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07740__S0 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11992__A2 net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07235_ net741 _01568_ net667 vssd1 vssd1 vccd1 vccd1 _02186_ sky130_fd_sc_hd__mux2_2
XFILLER_0_6_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout407_A _06255_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07757__S net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1149_A net1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09937__A2 net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07166_ final_design.cpu.reg_window\[906\] final_design.cpu.reg_window\[938\] net898
+ vssd1 vssd1 vccd1 vccd1 _02117_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07097_ final_design.cpu.reg_window\[972\] final_design.cpu.reg_window\[1004\] net897
+ vssd1 vssd1 vccd1 vccd1 _02048_ sky130_fd_sc_hd__mux2_1
XANTENNA__09257__B net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09825__X _04744_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout200 _06003_ vssd1 vssd1 vccd1 vccd1 net200 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout776_A net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1209 net1212 vssd1 vssd1 vccd1 vccd1 net1209 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout397_X net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout222 net223 vssd1 vssd1 vccd1 vccd1 net222 sky130_fd_sc_hd__buf_2
Xfanout233 _05983_ vssd1 vssd1 vccd1 vccd1 net233 sky130_fd_sc_hd__clkbuf_4
Xfanout244 _05910_ vssd1 vssd1 vccd1 vccd1 net244 sky130_fd_sc_hd__buf_2
XANTENNA__13430__CLK clknet_leaf_60_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10704__B1 net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout255 net259 vssd1 vssd1 vccd1 vccd1 net255 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_5_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09570__A0 _01626_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout266 net267 vssd1 vssd1 vccd1 vccd1 net266 sky130_fd_sc_hd__buf_6
Xfanout277 net279 vssd1 vssd1 vccd1 vccd1 net277 sky130_fd_sc_hd__buf_2
X_09807_ net482 _04366_ _04266_ vssd1 vssd1 vccd1 vccd1 _04726_ sky130_fd_sc_hd__a21oi_1
Xfanout288 net289 vssd1 vssd1 vccd1 vccd1 net288 sky130_fd_sc_hd__clkbuf_4
X_07999_ final_design.cpu.reg_window\[848\] final_design.cpu.reg_window\[880\] net843
+ vssd1 vssd1 vccd1 vccd1 _02950_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout564_X net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout943_A net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout299 _06159_ vssd1 vssd1 vccd1 vccd1 net299 sky130_fd_sc_hd__buf_4
XANTENNA__11308__A net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09738_ net728 _04639_ _04653_ _04656_ vssd1 vssd1 vccd1 vccd1 _04657_ sky130_fd_sc_hd__a31o_1
XANTENNA__09858__D1 net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13580__CLK clknet_leaf_47_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout731_X net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09669_ _02801_ net440 vssd1 vssd1 vccd1 vccd1 _04588_ sky130_fd_sc_hd__nand2_1
XFILLER_0_70_1518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout829_X net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11742__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11700_ net559 net421 _06208_ net294 net1600 vssd1 vssd1 vccd1 vccd1 _00481_ sky130_fd_sc_hd__a32o_1
X_12680_ _06327_ net1481 net979 vssd1 vssd1 vccd1 vccd1 _01342_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11680__A1 net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12209__B1 net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11631_ net209 net632 vssd1 vssd1 vccd1 vccd1 _06173_ sky130_fd_sc_hd__and2_1
XFILLER_0_77_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12224__A3 net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1403 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11562_ net212 net634 vssd1 vssd1 vccd1 vccd1 _06137_ sky130_fd_sc_hd__and2_1
XFILLER_0_64_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10513_ net964 _05261_ vssd1 vssd1 vccd1 vccd1 _05262_ sky130_fd_sc_hd__or2_1
XANTENNA__11983__A2 net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13301_ clknet_leaf_56_clk _00532_ net1144 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[289\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11493_ net181 net2514 net308 vssd1 vssd1 vccd1 vccd1 _00368_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_10_clk_X clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13232_ clknet_leaf_33_clk _00463_ net1231 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[220\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input72_A memory_size[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11697__B net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10444_ _02894_ net593 vssd1 vssd1 vccd1 vccd1 _05206_ sky130_fd_sc_hd__nor2_1
XFILLER_0_61_971 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14086__CLK clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12870__Q final_design.data_from_mem\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13163_ clknet_leaf_38_clk _00394_ net1187 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[151\]
+ sky130_fd_sc_hd__dfrtp_1
X_10375_ net18 net1025 net1008 final_design.data_from_mem\[24\] vssd1 vssd1 vccd1
+ vccd1 _00128_ sky130_fd_sc_hd__a22o_1
XANTENNA__09167__B net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08600__A2 _03550_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12114_ net1788 net200 net388 vssd1 vssd1 vccd1 vccd1 _00838_ sky130_fd_sc_hd__mux2_1
X_13094_ clknet_leaf_50_clk _00325_ net1168 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[82\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_62_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14233__1287 vssd1 vssd1 vccd1 vccd1 _14233__1287/HI net1287 sky130_fd_sc_hd__conb_1
XANTENNA__11917__S net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_25_clk_X clknet_leaf_25_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12045_ net1719 net202 net399 vssd1 vssd1 vccd1 vccd1 _00773_ sky130_fd_sc_hd__mux2_1
XANTENNA__09156__A3 _01815_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08498__S net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07798__S0 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13923__CLK clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13996_ clknet_leaf_46_clk _01227_ net1214 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[984\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09313__A0 net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12947_ clknet_leaf_29_clk _00185_ net1194 vssd1 vssd1 vccd1 vccd1 net104 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_1885 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12878_ clknet_leaf_17_clk _00116_ net1113 vssd1 vssd1 vccd1 vccd1 final_design.data_from_mem\[12\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__07431__A net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09077__C1 net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11829_ net201 net2102 net265 vssd1 vssd1 vccd1 vccd1 _00581_ sky130_fd_sc_hd__mux2_1
XANTENNA__12215__A3 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11423__A1 net209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13303__CLK clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11974__A2 net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11240__X _05943_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08533__Y _03484_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1801 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07020_ final_design.cpu.reg_window\[334\] final_design.cpu.reg_window\[366\] net906
+ vssd1 vssd1 vccd1 vccd1 _01971_ sky130_fd_sc_hd__mux2_1
XANTENNA__09358__A _03484_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_49_Right_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11187__B1 _05843_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1845 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11726__A2 net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13453__CLK clknet_leaf_44_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_1889 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06602__A1 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08971_ final_design.CPU_instr_adr\[18\] _03793_ vssd1 vssd1 vccd1 vccd1 _03909_
+ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_36_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11827__S net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07922_ final_design.cpu.reg_window\[406\] final_design.cpu.reg_window\[438\] net839
+ vssd1 vssd1 vccd1 vccd1 _02873_ sky130_fd_sc_hd__mux2_1
Xhold19 net111 vssd1 vssd1 vccd1 vccd1 net1361 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09805__B _04723_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11602__A_N _02095_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07853_ _02803_ vssd1 vssd1 vccd1 vccd1 _02804_ sky130_fd_sc_hd__inv_2
XANTENNA__07606__A net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09524__C _04240_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08450__S1 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06804_ net742 _01498_ _01504_ _01754_ vssd1 vssd1 vccd1 vccd1 _01755_ sky130_fd_sc_hd__o211a_1
XFILLER_0_78_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07784_ net552 _02733_ vssd1 vssd1 vccd1 vccd1 _02735_ sky130_fd_sc_hd__or2_2
XPHY_EDGE_ROW_58_Right_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_1805 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06735_ _01668_ _01674_ _01685_ net884 vssd1 vssd1 vccd1 vccd1 _01686_ sky130_fd_sc_hd__a22oi_4
X_09523_ _04233_ _04235_ net476 vssd1 vssd1 vccd1 vccd1 _04442_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout357_A net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09454_ _04300_ _04303_ net476 vssd1 vssd1 vccd1 vccd1 _04373_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_49_1867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1099_A net1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1226 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11662__A1 net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06656__S net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06666_ final_design.cpu.reg_window\[922\] final_design.cpu.reg_window\[954\] net943
+ vssd1 vssd1 vccd1 vccd1 _01617_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_49_1878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09032__S net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06764__S1 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08405_ _02239_ _03354_ vssd1 vssd1 vccd1 vccd1 _03356_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_4_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09385_ net535 net534 net533 net532 net457 net465 vssd1 vssd1 vccd1 vccd1 _04304_
+ sky130_fd_sc_hd__mux4_1
X_06597_ final_design.cpu.reg_window\[348\] final_design.cpu.reg_window\[380\] net946
+ vssd1 vssd1 vccd1 vccd1 _01548_ sky130_fd_sc_hd__mux2_1
XANTENNA__12206__A3 net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08336_ _03274_ _03275_ _03286_ net874 vssd1 vssd1 vccd1 vccd1 _03287_ sky130_fd_sc_hd__a22oi_4
XANTENNA__11965__A2 net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07094__A1 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12393__S net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08267_ final_design.cpu.reg_window\[714\] final_design.cpu.reg_window\[746\] net817
+ vssd1 vssd1 vccd1 vccd1 _03218_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout312_X net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_67_Right_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_1901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07218_ _02165_ _02166_ _02167_ _02168_ net765 net780 vssd1 vssd1 vccd1 vccd1 _02169_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_15_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08198_ final_design.cpu.reg_window\[782\] final_design.cpu.reg_window\[814\] net825
+ vssd1 vssd1 vccd1 vccd1 _03149_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07149_ _02099_ vssd1 vssd1 vccd1 vccd1 _02100_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_1475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1355 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09791__A0 net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10160_ _05042_ _05054_ _05055_ vssd1 vssd1 vccd1 vccd1 final_design.vga.h_next_count\[5\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_63_1388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout681_X net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13946__CLK clknet_leaf_63_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1006 _05171_ vssd1 vssd1 vccd1 vccd1 net1006 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11737__S net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout779_X net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09138__A3 net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10091_ _05000_ _05005_ _05004_ vssd1 vssd1 vccd1 vccd1 _05007_ sky130_fd_sc_hd__a21oi_1
Xfanout1017 _01411_ vssd1 vssd1 vccd1 vccd1 net1017 sky130_fd_sc_hd__buf_4
Xfanout1028 net1029 vssd1 vssd1 vccd1 vccd1 net1028 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout1039 _01394_ vssd1 vssd1 vccd1 vccd1 net1039 sky130_fd_sc_hd__buf_2
XANTENNA__07075__X _02026_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11350__B1 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_76_Right_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13850_ clknet_leaf_58_clk _01081_ net1125 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[838\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12972__RESET_B net1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12970__CLK clknet_leaf_15_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10993_ net86 net1045 vssd1 vssd1 vccd1 vccd1 _05719_ sky130_fd_sc_hd__or2_1
X_13781_ clknet_leaf_57_clk _01012_ net1145 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[769\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11472__S net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12732_ _06372_ vssd1 vssd1 vccd1 vccd1 _06373_ sky130_fd_sc_hd__inv_2
XFILLER_0_70_1326 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06566__S net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13326__CLK clknet_leaf_43_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1845 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_52_clk_A clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12663_ final_design.VGA_data_control.ready_data\[19\] net1021 net976 final_design.data_from_mem\[19\]
+ vssd1 vssd1 vccd1 vccd1 _06319_ sky130_fd_sc_hd__a22o_1
XFILLER_0_2_1709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_1889 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_2278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11614_ net563 net421 _06164_ net298 net1488 vssd1 vssd1 vccd1 vccd1 _00439_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_61_2289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12594_ final_design.reqhand.instruction\[12\] net997 net983 final_design.data_from_mem\[12\]
+ vssd1 vssd1 vccd1 vccd1 _01287_ sky130_fd_sc_hd__a22o_1
XFILLER_0_4_1591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11545_ net427 net563 _06128_ net302 net1622 vssd1 vssd1 vccd1 vccd1 _00406_ sky130_fd_sc_hd__a32o_1
XFILLER_0_0_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13476__CLK clknet_leaf_54_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11501__A net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11476_ net201 net2440 net309 vssd1 vssd1 vccd1 vccd1 _00357_ sky130_fd_sc_hd__mux2_1
XANTENNA__11708__A2 net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10427_ _03160_ _05190_ vssd1 vssd1 vccd1 vccd1 _05197_ sky130_fd_sc_hd__nor2_1
X_13215_ clknet_leaf_8_clk _00446_ net1134 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[203\]
+ sky130_fd_sc_hd__dfrtp_1
X_14195_ net1253 vssd1 vssd1 vccd1 vccd1 gpio_oeb[7] sky130_fd_sc_hd__buf_2
XANTENNA__13007__RESET_B net1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08585__A1 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13146_ clknet_leaf_6_clk _00377_ net1128 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[134\]
+ sky130_fd_sc_hd__dfrtp_1
X_10358_ net31 net1023 net1007 net2546 vssd1 vssd1 vccd1 vccd1 _00111_ sky130_fd_sc_hd__o22a_1
XANTENNA__06691__S0 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13077_ clknet_leaf_7_clk _00308_ net1145 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[65\]
+ sky130_fd_sc_hd__dfrtp_1
X_10289_ net1533 net1039 vssd1 vssd1 vccd1 vccd1 _00000_ sky130_fd_sc_hd__and2_1
XFILLER_0_57_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12028_ net2001 net228 net397 vssd1 vssd1 vccd1 vccd1 _00756_ sky130_fd_sc_hd__mux2_1
XANTENNA__11341__B1 net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14101__CLK clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06899__A1 net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13979_ clknet_leaf_65_clk _01210_ net1070 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[967\]
+ sky130_fd_sc_hd__dfrtp_1
X_06520_ net1039 net994 net991 _01470_ vssd1 vssd1 vccd1 vccd1 _01471_ sky130_fd_sc_hd__o31a_1
XANTENNA__11644__A1 net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10447__A2 net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06746__S1 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06451_ _01397_ _01400_ _01403_ _01404_ net1039 vssd1 vssd1 vccd1 vccd1 _01405_ sky130_fd_sc_hd__a221o_2
XTAP_TAPCELL_ROW_44_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13819__CLK clknet_leaf_65_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09170_ _03628_ _03650_ vssd1 vssd1 vccd1 vccd1 _04089_ sky130_fd_sc_hd__nor2_1
XFILLER_0_43_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08121_ _02030_ net600 vssd1 vssd1 vccd1 vccd1 _03072_ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11947__A2 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08052_ _02999_ _03000_ _03001_ _03002_ net682 net693 vssd1 vssd1 vccd1 vccd1 _03003_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_3_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_1328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12843__CLK clknet_leaf_15_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload44_A clknet_leaf_36_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07003_ net749 _01947_ net745 vssd1 vssd1 vccd1 vccd1 _01954_ sky130_fd_sc_hd__o21a_1
XANTENNA__13969__CLK clknet_leaf_34_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11130__B _05843_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_1041 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06587__B1 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08954_ _03655_ _03893_ net1038 vssd1 vssd1 vccd1 vccd1 _03894_ sky130_fd_sc_hd__o21a_1
XANTENNA__11784__C net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1014_A net1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07905_ _02852_ _02853_ _02854_ _02855_ net683 net693 vssd1 vssd1 vccd1 vccd1 _02856_
+ sky130_fd_sc_hd__mux4_1
X_08885_ _03773_ _03831_ vssd1 vssd1 vccd1 vccd1 _03832_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout474_A _03485_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07836_ final_design.cpu.reg_window\[789\] final_design.cpu.reg_window\[821\] net858
+ vssd1 vssd1 vccd1 vccd1 _02787_ sky130_fd_sc_hd__mux2_1
XANTENNA__07770__S net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13349__CLK clknet_leaf_52_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout641_A _05946_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07767_ net719 _02717_ vssd1 vssd1 vccd1 vccd1 _02718_ sky130_fd_sc_hd__or2_1
XANTENNA__12388__S net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09506_ _04385_ _04387_ vssd1 vssd1 vccd1 vccd1 _04425_ sky130_fd_sc_hd__or2_1
XFILLER_0_39_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06718_ final_design.cpu.reg_window\[344\] final_design.cpu.reg_window\[376\] net944
+ vssd1 vssd1 vccd1 vccd1 _01669_ sky130_fd_sc_hd__mux2_1
X_07698_ net711 _02648_ vssd1 vssd1 vccd1 vccd1 _02649_ sky130_fd_sc_hd__nor2_1
XFILLER_0_67_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06649_ _01596_ _01599_ vssd1 vssd1 vccd1 vccd1 _01600_ sky130_fd_sc_hd__nand2_1
XFILLER_0_36_1799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09437_ net727 _04333_ _04355_ vssd1 vssd1 vccd1 vccd1 _04356_ sky130_fd_sc_hd__or3_2
XANTENNA__13499__CLK clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout906_A net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout527_X net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14232__1286 vssd1 vssd1 vccd1 vccd1 _14232__1286/HI net1286 sky130_fd_sc_hd__conb_1
X_09368_ net86 _04193_ net87 vssd1 vssd1 vccd1 vccd1 _04287_ sky130_fd_sc_hd__o21ai_1
XANTENNA__09687__S0 net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11399__B1 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08319_ final_design.cpu.reg_window\[8\] final_design.cpu.reg_window\[40\] net812
+ vssd1 vssd1 vccd1 vccd1 _03270_ sky130_fd_sc_hd__mux2_1
XANTENNA__10636__S net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09299_ _02503_ _03419_ vssd1 vssd1 vccd1 vccd1 _04218_ sky130_fd_sc_hd__nor2_1
XFILLER_0_65_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11330_ _04333_ _04355_ net656 vssd1 vssd1 vccd1 vccd1 _06023_ sky130_fd_sc_hd__o21ai_1
X_11261_ net736 _03940_ _05961_ vssd1 vssd1 vccd1 vccd1 _05962_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_28_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13000_ net1331 _00231_ net1196 vssd1 vssd1 vccd1 vccd1 final_design.CPU_instr_adr\[20\]
+ sky130_fd_sc_hd__dfrtp_4
X_10212_ final_design.uart.BAUD_counter\[4\] _05094_ net800 vssd1 vssd1 vccd1 vccd1
+ _05096_ sky130_fd_sc_hd__o21ai_1
XANTENNA__11020__C1 net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11192_ final_design.reqhand.data_from_UART\[6\] net251 vssd1 vssd1 vccd1 vccd1 _05901_
+ sky130_fd_sc_hd__nand2b_1
XFILLER_0_63_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10374__B2 final_design.data_from_mem\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_2683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11571__B1 net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_2060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_1196 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_2694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11467__S net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10143_ final_design.vga.h_current_state\[1\] _05011_ _05043_ vssd1 vssd1 vccd1 vccd1
+ _05044_ sky130_fd_sc_hd__or3_1
XANTENNA__14124__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06673__S0 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input35_A gpio_in[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10074_ net668 _04991_ vssd1 vssd1 vccd1 vccd1 _04992_ sky130_fd_sc_hd__nor2_1
XFILLER_0_27_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08414__S1 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13902_ clknet_leaf_43_clk _01133_ net1216 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[890\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_1535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_1568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07680__S net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13833_ clknet_leaf_33_clk _01064_ net1231 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[821\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12298__S net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_2487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_2498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11626__A1 net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13764_ clknet_leaf_54_clk _00995_ net1179 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[752\]
+ sky130_fd_sc_hd__dfrtp_1
X_10976_ _05701_ _05702_ vssd1 vssd1 vccd1 vccd1 _05703_ sky130_fd_sc_hd__nor2_1
XFILLER_0_54_1877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06728__S1 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12715_ _06348_ _06352_ vssd1 vssd1 vccd1 vccd1 _06356_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_35_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13695_ clknet_leaf_8_clk _00926_ net1130 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[683\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1528 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12646_ _06310_ net1414 net978 vssd1 vssd1 vccd1 vccd1 _01325_ sky130_fd_sc_hd__mux2_1
XANTENNA__12866__CLK clknet_leaf_25_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11929__A2 net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09452__C1 _04370_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12577_ net2423 _06293_ _06286_ vssd1 vssd1 vccd1 vccd1 _01273_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11528_ net1960 net190 net523 vssd1 vssd1 vccd1 vccd1 _00395_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold308 final_design.VGA_data_control.ready_data\[8\] vssd1 vssd1 vccd1 vccd1 net1650
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold319 final_design.cpu.reg_window\[451\] vssd1 vssd1 vccd1 vccd1 net1661 sky130_fd_sc_hd__dlygate4sd3_1
X_14247_ net1301 vssd1 vssd1 vccd1 vccd1 gpio_out[25] sky130_fd_sc_hd__buf_2
XFILLER_0_26_1913 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11459_ net243 net2173 net306 vssd1 vssd1 vccd1 vccd1 _00346_ sky130_fd_sc_hd__mux2_1
XANTENNA__12354__A2 net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14178_ clknet_leaf_22_clk _01352_ net1164 vssd1 vssd1 vccd1 vccd1 final_design.VGA_adr\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10365__B2 final_design.data_from_mem\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13129_ clknet_leaf_36_clk _00360_ net1236 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[117\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07156__A net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1008 final_design.cpu.reg_window\[351\] vssd1 vssd1 vccd1 vccd1 net2350 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1019 final_design.cpu.reg_window\[610\] vssd1 vssd1 vccd1 vccd1 net2361 sky130_fd_sc_hd__dlygate4sd3_1
X_08670_ _01481_ _01487_ _03620_ vssd1 vssd1 vccd1 vccd1 _03621_ sky130_fd_sc_hd__o21ai_1
XANTENNA__10668__A2 final_design.VGA_adr\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07621_ net605 _02570_ _02546_ vssd1 vssd1 vccd1 vccd1 _02572_ sky130_fd_sc_hd__o21ai_2
X_07552_ net885 _02495_ _02501_ _02488_ _02489_ vssd1 vssd1 vccd1 vccd1 _02503_ sky130_fd_sc_hd__a32o_4
XANTENNA__11406__A net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13641__CLK clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1917 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06503_ _01375_ net1039 net994 net991 vssd1 vssd1 vccd1 vccd1 _01454_ sky130_fd_sc_hd__or4_2
XFILLER_0_48_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07483_ _02300_ _02433_ _02298_ vssd1 vssd1 vccd1 vccd1 _02434_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_9_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11840__S net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06434_ final_design.vga.h_current_state\[0\] vssd1 vssd1 vccd1 vccd1 _01389_ sky130_fd_sc_hd__inv_2
XFILLER_0_75_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09222_ _04136_ _04140_ _04139_ _03133_ vssd1 vssd1 vccd1 vccd1 _04141_ sky130_fd_sc_hd__a211o_1
XFILLER_0_33_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13791__CLK clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09153_ _03652_ net447 vssd1 vssd1 vccd1 vccd1 _04072_ sky130_fd_sc_hd__nand2_4
XANTENNA__07049__A1 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07049__B2 _01999_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout222_A net223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08104_ final_design.cpu.reg_window\[780\] final_design.cpu.reg_window\[812\] net816
+ vssd1 vssd1 vccd1 vccd1 _03055_ sky130_fd_sc_hd__mux2_1
XANTENNA__12593__A2 net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09084_ _03785_ _04008_ vssd1 vssd1 vccd1 vccd1 _04009_ sky130_fd_sc_hd__or2_1
XFILLER_0_47_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08035_ final_design.cpu.reg_window\[659\] final_design.cpu.reg_window\[691\] net821
+ vssd1 vssd1 vccd1 vccd1 _02986_ sky130_fd_sc_hd__mux2_1
XANTENNA__13021__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput80 memory_size[20] vssd1 vssd1 vccd1 vccd1 net80 sky130_fd_sc_hd__clkbuf_2
XANTENNA__14147__CLK clknet_leaf_19_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10980__A net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold820 final_design.cpu.reg_window\[70\] vssd1 vssd1 vccd1 vccd1 net2162 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_47_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput91 memory_size[30] vssd1 vssd1 vccd1 vccd1 net91 sky130_fd_sc_hd__buf_1
XANTENNA_fanout1131_A net1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold831 final_design.cpu.reg_window\[103\] vssd1 vssd1 vccd1 vccd1 net2173 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08549__A1 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07765__S net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold842 final_design.cpu.reg_window\[521\] vssd1 vssd1 vccd1 vccd1 net2184 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12345__A2 net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09746__B1 _04341_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold853 final_design.cpu.reg_window\[443\] vssd1 vssd1 vccd1 vccd1 net2195 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09546__A net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold864 final_design.cpu.reg_window\[144\] vssd1 vssd1 vccd1 vccd1 net2206 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10356__A1 net29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold875 final_design.cpu.reg_window\[1006\] vssd1 vssd1 vccd1 vccd1 net2217 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout689_A net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold886 final_design.cpu.reg_window\[232\] vssd1 vssd1 vccd1 vccd1 net2228 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold897 final_design.cpu.reg_window\[830\] vssd1 vssd1 vccd1 vccd1 net2239 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06655__S0 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09986_ _04887_ _04904_ vssd1 vssd1 vccd1 vccd1 _04905_ sky130_fd_sc_hd__xnor2_2
XANTENNA_fanout1017_X net1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13171__CLK clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08937_ _03878_ vssd1 vssd1 vccd1 vccd1 _03879_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout856_A net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout477_X net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08868_ _02475_ _03816_ vssd1 vssd1 vccd1 vccd1 _03817_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07524__A2 _01570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08182__C1 net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07819_ _02769_ vssd1 vssd1 vccd1 vccd1 _02770_ sky130_fd_sc_hd__inv_2
XFILLER_0_54_1118 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08799_ _03676_ _03749_ vssd1 vssd1 vccd1 vccd1 _03750_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout644_X net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11316__A net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10830_ _05543_ _05563_ _05562_ vssd1 vssd1 vccd1 vccd1 _05564_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11608__B2 net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12889__CLK clknet_leaf_17_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07005__S net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_2963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_2340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10761_ _05496_ _05497_ vssd1 vssd1 vccd1 vccd1 _05498_ sky130_fd_sc_hd__nor2_1
XANTENNA__12281__A1 net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_2974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_2985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11750__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout909_X net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12500_ _06162_ net349 net327 net1649 vssd1 vssd1 vccd1 vccd1 _01205_ sky130_fd_sc_hd__a22o_1
XFILLER_0_48_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10692_ net960 _05430_ _05431_ _04042_ vssd1 vssd1 vccd1 vccd1 _05432_ sky130_fd_sc_hd__a22o_1
X_13480_ clknet_leaf_41_clk _00711_ net1224 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[468\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_48_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12431_ _06246_ _06260_ vssd1 vssd1 vccd1 vccd1 _06282_ sky130_fd_sc_hd__nor2_1
XFILLER_0_63_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06416__Y _01371_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12584__A2 net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12362_ net2452 net362 net354 _06090_ vssd1 vssd1 vccd1 vccd1 _01074_ sky130_fd_sc_hd__a22o_1
XANTENNA__10595__A1 net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_2892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_2111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10595__B2 net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11792__B1 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14101_ clknet_leaf_9_clk _01298_ net1103 vssd1 vssd1 vccd1 vccd1 final_design.reqhand.instruction\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_11313_ _01823_ net642 _06005_ _06006_ net656 vssd1 vssd1 vccd1 vccd1 _06008_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_56_2122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_2756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12293_ net584 _06223_ net513 net370 net2153 vssd1 vssd1 vccd1 vccd1 _01008_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_56_2133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_2767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_2778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12336__A2 net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14032_ clknet_leaf_33_clk _01263_ net1238 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[1020\]
+ sky130_fd_sc_hd__dfrtp_1
X_11244_ net744 _01480_ vssd1 vssd1 vccd1 vccd1 _05947_ sky130_fd_sc_hd__nand2_2
XANTENNA__13514__CLK clknet_leaf_60_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11175_ net735 _04016_ _05885_ vssd1 vssd1 vccd1 vccd1 _05886_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_78_1619 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10126_ _04999_ _05033_ vssd1 vssd1 vccd1 vccd1 final_design.vga.v_next_count\[8\]
+ sky130_fd_sc_hd__and2_1
XANTENNA__14140__RESET_B net1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_66_Left_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08399__S0 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10057_ net68 _04940_ _04954_ _04956_ _04657_ vssd1 vssd1 vccd1 vccd1 _04976_ sky130_fd_sc_hd__o221ai_2
XANTENNA__13664__CLK clknet_leaf_11_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_2549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07704__A net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06723__B1 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkload0_A clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13816_ clknet_leaf_65_clk _01047_ net1073 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[804\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13747_ clknet_leaf_39_clk _00978_ net1206 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[735\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07142__C net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10959_ net1055 _05683_ net1000 final_design.CPU_instr_adr\[24\] vssd1 vssd1 vccd1
+ vccd1 _05687_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_35_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_1461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06754__S net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13678_ clknet_leaf_44_clk _00909_ net1208 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[666\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_75_Left_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_1358 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12629_ final_design.VGA_data_control.ready_data\[2\] net1022 net976 final_design.data_from_mem\[2\]
+ vssd1 vssd1 vccd1 vccd1 _06302_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_14_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13044__CLK clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1382 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07126__S1 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold105 final_design.VGA_data_control.data_to_VGA\[9\] vssd1 vssd1 vccd1 vccd1 net1447
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold116 final_design.reqhand.instruction\[25\] vssd1 vssd1 vccd1 vccd1 net1458 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06885__S0 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold127 final_design.cpu.reg_window\[202\] vssd1 vssd1 vccd1 vccd1 net1469 sky130_fd_sc_hd__dlygate4sd3_1
Xhold138 final_design.reqhand.instruction\[19\] vssd1 vssd1 vccd1 vccd1 net1480 sky130_fd_sc_hd__dlygate4sd3_1
Xhold149 final_design.cpu.reg_window\[734\] vssd1 vssd1 vccd1 vccd1 net1491 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13194__CLK clknet_leaf_61_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10338__B2 final_design.data_from_mem\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06637__S0 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09840_ _04517_ _04524_ net495 vssd1 vssd1 vccd1 vccd1 _04759_ sky130_fd_sc_hd__a21oi_2
Xfanout607 _02514_ vssd1 vssd1 vccd1 vccd1 net607 sky130_fd_sc_hd__buf_2
Xfanout618 _02513_ vssd1 vssd1 vccd1 vccd1 net618 sky130_fd_sc_hd__clkbuf_2
Xfanout629 _06192_ vssd1 vssd1 vccd1 vccd1 net629 sky130_fd_sc_hd__buf_4
XFILLER_0_0_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14231__1285 vssd1 vssd1 vccd1 vccd1 _14231__1285/HI net1285 sky130_fd_sc_hd__conb_1
XANTENNA__08951__B2 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09771_ _04642_ _04644_ net480 vssd1 vssd1 vccd1 vccd1 _04690_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06983_ final_design.cpu.reg_window\[528\] final_design.cpu.reg_window\[560\] net923
+ vssd1 vssd1 vccd1 vccd1 _01934_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11835__S net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08722_ final_design.CPU_instr_adr\[18\] _01881_ vssd1 vssd1 vccd1 vccd1 _03673_
+ sky130_fd_sc_hd__nand2_1
XANTENNA__09900__B1 net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07062__S0 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08653_ _02610_ _02642_ _03603_ vssd1 vssd1 vccd1 vccd1 _03604_ sky130_fd_sc_hd__and3_1
XANTENNA__10510__A1 net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10510__B2 net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07604_ final_design.cpu.reg_window\[157\] final_design.cpu.reg_window\[189\] net870
+ vssd1 vssd1 vccd1 vccd1 _02555_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08584_ net717 _03534_ vssd1 vssd1 vccd1 vccd1 _03535_ sky130_fd_sc_hd__or2_1
XFILLER_0_72_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07535_ final_design.cpu.reg_window\[159\] final_design.cpu.reg_window\[191\] net937
+ vssd1 vssd1 vccd1 vccd1 _02486_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout1081_A net1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout437_A _05847_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07466_ _02413_ _02414_ _02415_ _02416_ net768 net781 vssd1 vssd1 vccd1 vccd1 _02417_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__06517__X _01468_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06664__S net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06417_ net1 vssd1 vssd1 vccd1 vccd1 _01372_ sky130_fd_sc_hd__inv_2
X_09205_ _03631_ _04053_ vssd1 vssd1 vccd1 vccd1 _04124_ sky130_fd_sc_hd__or2_4
XFILLER_0_63_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07397_ final_design.cpu.reg_window\[770\] final_design.cpu.reg_window\[802\] net914
+ vssd1 vssd1 vccd1 vccd1 _02348_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09136_ _03629_ _04053_ vssd1 vssd1 vccd1 vccd1 _04055_ sky130_fd_sc_hd__or2_2
XFILLER_0_32_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10577__A1 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13537__CLK clknet_leaf_47_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10577__B2 net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12776__7 clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 net1317 sky130_fd_sc_hd__inv_2
X_09067_ final_design.CPU_instr_adr\[6\] _03785_ final_design.CPU_instr_adr\[7\] vssd1
+ vssd1 vccd1 vccd1 _03994_ sky130_fd_sc_hd__a21oi_1
X_08018_ final_design.cpu.reg_window\[467\] final_design.cpu.reg_window\[499\] net830
+ vssd1 vssd1 vccd1 vccd1 _02969_ sky130_fd_sc_hd__mux2_1
XANTENNA__10411__A1_N net250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold650 final_design.cpu.reg_window\[537\] vssd1 vssd1 vccd1 vccd1 net1992 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10329__B2 final_design.data_from_mem\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold661 final_design.cpu.reg_window\[918\] vssd1 vssd1 vccd1 vccd1 net2003 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout594_X net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout973_A _01415_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold672 final_design.cpu.reg_window\[570\] vssd1 vssd1 vccd1 vccd1 net2014 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold683 final_design.cpu.reg_window\[953\] vssd1 vssd1 vccd1 vccd1 net2025 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09195__B2 net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold694 final_design.cpu.reg_window\[333\] vssd1 vssd1 vccd1 vccd1 net2036 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13687__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1917 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout761_X net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09969_ _03324_ net441 net438 _03326_ vssd1 vssd1 vccd1 vccd1 _04888_ sky130_fd_sc_hd__o22a_1
XANTENNA__11745__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12980_ clknet_leaf_19_clk _00005_ net1156 vssd1 vssd1 vccd1 vccd1 wb_manage.curr_state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_11931_ net2468 net408 _06254_ net426 vssd1 vssd1 vccd1 vccd1 _00666_ sky130_fd_sc_hd__a22o_1
XANTENNA__10501__A1 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_2402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1901 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11862_ _06107_ net277 net517 net2018 vssd1 vssd1 vccd1 vccd1 _00610_ sky130_fd_sc_hd__a22o_1
XFILLER_0_24_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13601_ clknet_leaf_47_clk _00832_ net1203 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[589\]
+ sky130_fd_sc_hd__dfrtp_1
X_10813_ net77 net1044 vssd1 vssd1 vccd1 vccd1 _05547_ sky130_fd_sc_hd__and2_1
XANTENNA__12254__A1 net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13067__CLK clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11793_ net2442 net413 net283 _05997_ vssd1 vssd1 vccd1 vccd1 _00549_ sky130_fd_sc_hd__a22o_1
XANTENNA__11480__S net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13532_ clknet_leaf_3_clk _00763_ net1066 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[520\]
+ sky130_fd_sc_hd__dfrtp_1
X_10744_ _05478_ _05480_ net1004 vssd1 vssd1 vccd1 vccd1 _05482_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_39_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09670__A2 net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14255__1309 vssd1 vssd1 vccd1 vccd1 _14255__1309/HI net1309 sky130_fd_sc_hd__conb_1
X_13463_ clknet_leaf_6_clk _00694_ net1130 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[451\]
+ sky130_fd_sc_hd__dfrtp_1
X_10675_ net958 _05412_ _05415_ net955 vssd1 vssd1 vccd1 vccd1 _05416_ sky130_fd_sc_hd__o22a_1
XFILLER_0_10_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_77_2818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_2829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12414_ _06243_ net501 net340 net2040 vssd1 vssd1 vccd1 vccd1 _01124_ sky130_fd_sc_hd__a22o_1
XANTENNA__12557__A2 net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13394_ clknet_leaf_39_clk _00625_ net1208 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[382\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08642__X _03593_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1191 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12345_ _06233_ net498 net360 net2104 vssd1 vssd1 vccd1 vccd1 _01057_ sky130_fd_sc_hd__a22o_1
XANTENNA__12904__CLK clknet_leaf_61_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12276_ net561 _06206_ net503 net368 net1867 vssd1 vssd1 vccd1 vccd1 _00991_ sky130_fd_sc_hd__a32o_1
XFILLER_0_23_1905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14015_ clknet_leaf_7_clk _01246_ net1134 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[1003\]
+ sky130_fd_sc_hd__dfrtp_1
X_11227_ net732 _03968_ vssd1 vssd1 vccd1 vccd1 _05932_ sky130_fd_sc_hd__or2_1
XANTENNA__09725__A3 _01815_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09281__S1 net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08933__A1 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11158_ net1018 net734 _05870_ vssd1 vssd1 vccd1 vccd1 _05871_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_21_1640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10109_ final_design.VGA_data_control.v_count\[2\] _05019_ _05022_ vssd1 vssd1 vccd1
+ vccd1 final_design.vga.v_next_count\[2\] sky130_fd_sc_hd__a21oi_1
X_11089_ final_design.CPU_instr_adr\[30\] net1000 _05807_ net1056 vssd1 vssd1 vccd1
+ vccd1 _05811_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_76_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12493__A1 _06153_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11296__A2 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08249__B net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_79 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09646__C1 _04113_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07320_ final_design.cpu.reg_window\[324\] final_design.cpu.reg_window\[356\] net903
+ vssd1 vssd1 vccd1 vccd1 _02271_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09110__A1 final_design.CPU_instr_adr\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07251_ final_design.cpu.reg_window\[967\] final_design.cpu.reg_window\[999\] net892
+ vssd1 vssd1 vccd1 vccd1 _02202_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07672__A1 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12548__A2 net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07182_ final_design.cpu.reg_window\[457\] final_design.cpu.reg_window\[489\] net891
+ vssd1 vssd1 vccd1 vccd1 _02133_ sky130_fd_sc_hd__mux2_1
XANTENNA__11756__A0 net197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10019__B net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10734__S net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08712__B _01630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout404 net405 vssd1 vssd1 vccd1 vccd1 net404 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_6_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10035__A net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout415 _06227_ vssd1 vssd1 vccd1 vccd1 net415 sky130_fd_sc_hd__clkbuf_8
XANTENNA__08924__A1 _02507_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout426 net431 vssd1 vssd1 vccd1 vccd1 net426 sky130_fd_sc_hd__buf_2
Xfanout437 _05847_ vssd1 vssd1 vccd1 vccd1 net437 sky130_fd_sc_hd__buf_2
X_09823_ _03293_ _04153_ _04154_ _03290_ vssd1 vssd1 vccd1 vccd1 _04742_ sky130_fd_sc_hd__a31o_1
Xfanout448 net449 vssd1 vssd1 vccd1 vccd1 net448 sky130_fd_sc_hd__buf_4
Xfanout459 _03551_ vssd1 vssd1 vccd1 vccd1 net459 sky130_fd_sc_hd__buf_4
XANTENNA_fanout387_A _06266_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09754_ _03229_ _04503_ vssd1 vssd1 vccd1 vccd1 _04673_ sky130_fd_sc_hd__nand2_1
XANTENNA__06659__S net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06966_ _01913_ _01914_ _01915_ _01916_ net773 net791 vssd1 vssd1 vccd1 vccd1 _01917_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__09035__S net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08705_ final_design.CPU_instr_adr\[30\] _01507_ vssd1 vssd1 vccd1 vccd1 _03656_
+ sky130_fd_sc_hd__and2_1
XANTENNA__08688__B1 _02419_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09685_ net496 _04603_ _04602_ _04072_ vssd1 vssd1 vccd1 vccd1 _04604_ sky130_fd_sc_hd__a211o_1
XFILLER_0_55_1213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout554_A _06238_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06897_ _01844_ _01845_ _01846_ _01847_ net768 net781 vssd1 vssd1 vccd1 vccd1 _01848_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__10495__B1 net58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08636_ net603 _02961_ _02962_ _01938_ vssd1 vssd1 vccd1 vccd1 _03587_ sky130_fd_sc_hd__o211ai_4
XANTENNA__12236__A1 net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout342_X net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08567_ net608 _03513_ _03515_ vssd1 vssd1 vccd1 vccd1 _03518_ sky130_fd_sc_hd__a21oi_2
XANTENNA_fanout721_A _01720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout819_A net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07518_ _01686_ _01690_ _02468_ vssd1 vssd1 vccd1 vccd1 _02469_ sky130_fd_sc_hd__o21a_1
XFILLER_0_65_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08498_ _03443_ _03448_ net709 vssd1 vssd1 vccd1 vccd1 _03449_ sky130_fd_sc_hd__mux2_1
XANTENNA__11995__B1 net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12997__RESET_B net1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07449_ _02396_ _02397_ _02398_ _02399_ net768 net787 vssd1 vssd1 vccd1 vccd1 _02400_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_21_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout607_X net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12927__CLK clknet_leaf_47_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_1864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12539__A2 net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10460_ _02635_ net592 vssd1 vssd1 vccd1 vccd1 _05214_ sky130_fd_sc_hd__nor2_2
XANTENNA__06871__C1 _01821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12798__29_A clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11747__A0 net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09119_ net964 _04037_ vssd1 vssd1 vccd1 vccd1 _04038_ sky130_fd_sc_hd__nor2_1
X_10391_ _05176_ vssd1 vssd1 vccd1 vccd1 _05177_ sky130_fd_sc_hd__inv_2
XFILLER_0_81_1829 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12130_ _06094_ _06268_ _06267_ vssd1 vssd1 vccd1 vccd1 _00851_ sky130_fd_sc_hd__a21o_1
X_12061_ net804 _05839_ _05841_ vssd1 vssd1 vccd1 vccd1 _06264_ sky130_fd_sc_hd__and3_4
Xhold480 final_design.cpu.reg_window\[856\] vssd1 vssd1 vccd1 vccd1 net1822 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold491 final_design.cpu.reg_window\[86\] vssd1 vssd1 vccd1 vccd1 net1833 sky130_fd_sc_hd__dlygate4sd3_1
X_11012_ net87 net1045 vssd1 vssd1 vccd1 vccd1 _05737_ sky130_fd_sc_hd__nor2_1
XFILLER_0_25_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout960 _04040_ vssd1 vssd1 vccd1 vccd1 net960 sky130_fd_sc_hd__buf_4
XANTENNA__11328__X _06021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout971 _01415_ vssd1 vssd1 vccd1 vccd1 net971 sky130_fd_sc_hd__clkbuf_4
Xfanout982 net983 vssd1 vssd1 vccd1 vccd1 net982 sky130_fd_sc_hd__buf_2
Xfanout993 _01409_ vssd1 vssd1 vccd1 vccd1 net993 sky130_fd_sc_hd__buf_2
X_12963_ clknet_leaf_32_clk _00201_ net1234 vssd1 vssd1 vccd1 vccd1 net121 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1180 final_design.cpu.reg_window\[445\] vssd1 vssd1 vccd1 vccd1 net2522 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1191 final_design.cpu.reg_window\[311\] vssd1 vssd1 vccd1 vccd1 net2533 sky130_fd_sc_hd__dlygate4sd3_1
X_11914_ final_design.cpu.reg_window\[411\] _05845_ vssd1 vssd1 vccd1 vccd1 _06250_
+ sky130_fd_sc_hd__or2_1
X_12894_ clknet_leaf_21_clk _00132_ net1158 vssd1 vssd1 vccd1 vccd1 final_design.data_from_mem\[28\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_34_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13702__CLK clknet_leaf_51_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12227__A1 net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1887 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11845_ net231 net2339 net517 vssd1 vssd1 vccd1 vccd1 _00595_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07329__S1 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_16_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07260__Y _02211_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11776_ net2399 net412 net280 _05891_ vssd1 vssd1 vccd1 vccd1 _00535_ sky130_fd_sc_hd__a22o_1
XANTENNA__08085__A _01785_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09643__A2 _04559_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11986__B1 net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13515_ clknet_leaf_38_clk _00746_ net1188 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[503\]
+ sky130_fd_sc_hd__dfrtp_1
X_10727_ net73 net1043 vssd1 vssd1 vccd1 vccd1 _05465_ sky130_fd_sc_hd__and2_1
X_14230__1284 vssd1 vssd1 vccd1 vccd1 _14230__1284/HI net1284 sky130_fd_sc_hd__conb_1
XFILLER_0_71_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13852__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13446_ clknet_leaf_51_clk _00677_ net1170 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[434\]
+ sky130_fd_sc_hd__dfrtp_1
X_10658_ net37 _05399_ vssd1 vssd1 vccd1 vccd1 _05400_ sky130_fd_sc_hd__nand2_1
XANTENNA__11738__A0 net242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload14 clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 clkload14/X sky130_fd_sc_hd__clkbuf_4
Xclkload25 clknet_leaf_25_clk vssd1 vssd1 vccd1 vccd1 clkload25/Y sky130_fd_sc_hd__bufinv_16
Xclkload36 clknet_leaf_48_clk vssd1 vssd1 vccd1 vccd1 clkload36/Y sky130_fd_sc_hd__clkinvlp_4
XANTENNA__08603__B1 _03524_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11202__A2 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13377_ clknet_leaf_47_clk _00608_ net1202 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[365\]
+ sky130_fd_sc_hd__dfrtp_1
X_10589_ _05311_ _05333_ vssd1 vssd1 vccd1 vccd1 _05334_ sky130_fd_sc_hd__nor2_1
XFILLER_0_80_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12328_ net1862 net177 net366 vssd1 vssd1 vccd1 vccd1 _01042_ sky130_fd_sc_hd__mux2_1
X_12259_ net584 _06188_ net512 net374 net1549 vssd1 vssd1 vccd1 vccd1 _00975_ sky130_fd_sc_hd__a32o_1
XANTENNA__06917__B1 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11910__B1 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13232__CLK clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06820_ net754 _01770_ net748 vssd1 vssd1 vccd1 vccd1 _01771_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_30_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_3000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_3011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06751_ _01698_ _01699_ _01700_ _01701_ net772 net791 vssd1 vssd1 vccd1 vccd1 _01702_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_30_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_3022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_3033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_3044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_3055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09470_ _04356_ _04358_ vssd1 vssd1 vccd1 vccd1 _04389_ sky130_fd_sc_hd__nand2_1
X_06682_ final_design.cpu.reg_window\[345\] final_design.cpu.reg_window\[377\] net936
+ vssd1 vssd1 vccd1 vccd1 _01633_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_1408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13382__CLK clknet_leaf_52_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08421_ net715 _03365_ net724 vssd1 vssd1 vccd1 vccd1 _03372_ sky130_fd_sc_hd__o21a_1
XFILLER_0_59_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08352_ final_design.cpu.reg_window\[71\] final_design.cpu.reg_window\[103\] net806
+ vssd1 vssd1 vccd1 vccd1 _03303_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_1905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11977__B1 net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07303_ net752 _02253_ net746 vssd1 vssd1 vccd1 vccd1 _02254_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_24_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08283_ final_design.cpu.reg_window\[265\] final_design.cpu.reg_window\[297\] net810
+ vssd1 vssd1 vccd1 vccd1 _03234_ sky130_fd_sc_hd__mux2_1
Xclkload8 clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 clkload8/Y sky130_fd_sc_hd__clkinvlp_4
XANTENNA__07740__S1 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07234_ net881 _02177_ _02183_ _02170_ _02171_ vssd1 vssd1 vccd1 vccd1 _02185_ sky130_fd_sc_hd__a32o_4
XFILLER_0_41_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07165_ final_design.cpu.reg_window\[970\] final_design.cpu.reg_window\[1002\] net898
+ vssd1 vssd1 vccd1 vccd1 _02116_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout302_A net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1044_A final_design.VGA_adr\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07948__A2 _02894_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07096_ final_design.cpu.reg_window\[780\] final_design.cpu.reg_window\[812\] net897
+ vssd1 vssd1 vccd1 vccd1 _02047_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1211_A net1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout201 _05996_ vssd1 vssd1 vccd1 vccd1 net201 sky130_fd_sc_hd__clkbuf_2
Xfanout212 net213 vssd1 vssd1 vccd1 vccd1 net212 sky130_fd_sc_hd__clkbuf_2
Xfanout223 _05980_ vssd1 vssd1 vccd1 vccd1 net223 sky130_fd_sc_hd__clkbuf_2
XANTENNA__10704__A1 net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout234 _05983_ vssd1 vssd1 vccd1 vccd1 net234 sky130_fd_sc_hd__buf_1
XANTENNA_fanout671_A net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11901__A0 net223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout245 net247 vssd1 vssd1 vccd1 vccd1 net245 sky130_fd_sc_hd__buf_4
XANTENNA_fanout292_X net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout769_A net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout256 net257 vssd1 vssd1 vccd1 vccd1 net256 sky130_fd_sc_hd__clkbuf_4
X_09806_ _04704_ _04724_ vssd1 vssd1 vccd1 vccd1 _04725_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09570__A1 _01657_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08373__A2 _03321_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout267 _06237_ vssd1 vssd1 vccd1 vccd1 net267 sky130_fd_sc_hd__buf_6
XFILLER_0_5_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout278 net279 vssd1 vssd1 vccd1 vccd1 net278 sky130_fd_sc_hd__clkbuf_4
X_14254__1308 vssd1 vssd1 vccd1 vccd1 _14254__1308/HI net1308 sky130_fd_sc_hd__conb_1
X_07998_ net714 _02942_ net723 vssd1 vssd1 vccd1 vccd1 _02949_ sky130_fd_sc_hd__o21a_1
Xfanout289 net290 vssd1 vssd1 vccd1 vccd1 net289 sky130_fd_sc_hd__clkbuf_2
X_09737_ _04184_ _04655_ vssd1 vssd1 vccd1 vccd1 _04656_ sky130_fd_sc_hd__and2_1
XANTENNA__07008__S0 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11308__B net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12457__A1 net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13725__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06949_ final_design.cpu.reg_window\[913\] final_design.cpu.reg_window\[945\] net925
+ vssd1 vssd1 vccd1 vccd1 _01900_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout936_A net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_66_clk clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_66_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__09322__A1 net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09668_ _04583_ _04584_ _04586_ _04342_ vssd1 vssd1 vccd1 vccd1 _04587_ sky130_fd_sc_hd__o22a_1
XFILLER_0_74_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08619_ net538 _03194_ vssd1 vssd1 vccd1 vccd1 _03570_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout724_X net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11680__A2 net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09599_ net478 _04200_ vssd1 vssd1 vccd1 vccd1 _04518_ sky130_fd_sc_hd__and2_1
XFILLER_0_38_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11324__A net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13875__CLK clknet_leaf_36_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11630_ net425 net560 _06172_ net298 net1683 vssd1 vssd1 vccd1 vccd1 _00447_ sky130_fd_sc_hd__a32o_1
XANTENNA__08145__A1_N net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11968__B1 net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11561_ net429 net568 _06136_ net303 net1644 vssd1 vssd1 vccd1 vccd1 _00414_ sky130_fd_sc_hd__a32o_1
XFILLER_0_68_1415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_939 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13300_ clknet_leaf_9_clk _00531_ net1104 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[288\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_64_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10512_ final_design.CPU_instr_adr\[3\] net1001 _05255_ net1042 vssd1 vssd1 vccd1
+ vccd1 _05261_ sky130_fd_sc_hd__o22a_1
XANTENNA__06852__S net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13105__CLK clknet_leaf_34_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11492_ net181 _06093_ vssd1 vssd1 vccd1 vccd1 _06114_ sky130_fd_sc_hd__and2_1
X_13231_ clknet_leaf_43_clk _00462_ net1218 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[219\]
+ sky130_fd_sc_hd__dfrtp_1
X_10443_ net1459 net1035 _05205_ net248 vssd1 vssd1 vccd1 vccd1 _00162_ sky130_fd_sc_hd__a22o_1
XFILLER_0_33_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09448__B _04366_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input65_A mem_adr_start[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13162_ clknet_leaf_61_clk _00393_ net1140 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[150\]
+ sky130_fd_sc_hd__dfrtp_1
X_10374_ net17 net1024 net1006 final_design.data_from_mem\[23\] vssd1 vssd1 vccd1
+ vccd1 _00127_ sky130_fd_sc_hd__o22a_1
XFILLER_0_62_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12113_ net1859 net202 net391 vssd1 vssd1 vccd1 vccd1 _00837_ sky130_fd_sc_hd__mux2_1
XANTENNA__13255__CLK clknet_leaf_62_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13093_ clknet_leaf_49_clk _00324_ net1184 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[81\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07683__S net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07247__S0 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12044_ net1676 net203 net399 vssd1 vssd1 vccd1 vccd1 _00772_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07798__S1 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout790 _01418_ vssd1 vssd1 vccd1 vccd1 net790 sky130_fd_sc_hd__buf_4
X_13995_ clknet_leaf_53_clk _01226_ net1188 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[983\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_57_clk clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_57_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__09313__A1 net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08116__A2 _03065_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12946_ clknet_leaf_29_clk _00184_ net1193 vssd1 vssd1 vccd1 vccd1 net103 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_62_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12877_ clknet_leaf_17_clk _00115_ net1108 vssd1 vssd1 vccd1 vccd1 final_design.data_from_mem\[11\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_73_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11234__A net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11828_ net204 net2134 net266 vssd1 vssd1 vccd1 vccd1 _00580_ sky130_fd_sc_hd__mux2_1
XANTENNA__08019__S net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10306__S0 net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11959__B1 net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12620__A1 final_design.reqhand.data_from_UART\[6\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_3_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11759_ net193 net2055 net418 vssd1 vssd1 vccd1 vccd1 _00522_ sky130_fd_sc_hd__mux2_1
XANTENNA__10792__B net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14030__CLK clknet_leaf_43_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13429_ clknet_leaf_56_clk _00660_ net1149 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[417\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_64_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09475__S1 net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1857 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xmax_cap968 _01472_ vssd1 vssd1 vccd1 vccd1 net968 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_80_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08970_ _02458_ net625 _03905_ _03907_ net258 vssd1 vssd1 vccd1 vccd1 _03908_ sky130_fd_sc_hd__a311o_1
XANTENNA__14180__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_36_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07921_ final_design.cpu.reg_window\[470\] final_design.cpu.reg_window\[502\] net839
+ vssd1 vssd1 vccd1 vccd1 _02872_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_36_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13748__CLK clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09001__B1 net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12687__B2 final_design.data_from_mem\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07852_ _02800_ _02801_ vssd1 vssd1 vccd1 vccd1 _02803_ sky130_fd_sc_hd__nor2_2
XANTENNA_wire525_X net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06803_ net742 _01752_ vssd1 vssd1 vccd1 vccd1 _01754_ sky130_fd_sc_hd__nand2_1
XANTENNA__12439__A1 net244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput1 ACK_I vssd1 vssd1 vccd1 vccd1 net1 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_39_1038 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07783_ net615 _02731_ _02732_ _01686_ vssd1 vssd1 vccd1 vccd1 _02734_ sky130_fd_sc_hd__a211oi_1
Xclkbuf_leaf_48_clk clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_48_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_79_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09522_ _04084_ _04440_ vssd1 vssd1 vccd1 vccd1 _04441_ sky130_fd_sc_hd__and2_1
X_06734_ _01679_ _01684_ net753 vssd1 vssd1 vccd1 vccd1 _01685_ sky130_fd_sc_hd__mux2_1
XANTENNA__13898__CLK clknet_leaf_59_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1817 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09453_ net493 _04342_ _04368_ _04371_ vssd1 vssd1 vccd1 vccd1 _04372_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_49_1868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06665_ final_design.cpu.reg_window\[986\] final_design.cpu.reg_window\[1018\] net943
+ vssd1 vssd1 vccd1 vccd1 _01616_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_49_1879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11662__A2 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout252_A net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_26_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08404_ net610 _03352_ _03353_ _02239_ vssd1 vssd1 vccd1 vccd1 _03355_ sky130_fd_sc_hd__a211oi_2
X_09384_ net540 net539 _02091_ net537 net457 net466 vssd1 vssd1 vccd1 vccd1 _04303_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__13128__CLK clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06596_ net761 _01546_ vssd1 vssd1 vccd1 vccd1 _01547_ sky130_fd_sc_hd__or2_1
X_08335_ _03280_ _03285_ net707 vssd1 vssd1 vccd1 vccd1 _03286_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout1161_A net1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12611__B2 final_design.data_from_mem\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout517_A net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08266_ _03213_ _03214_ _03215_ _03216_ net676 net697 vssd1 vssd1 vccd1 vccd1 _03217_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_62_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07217_ final_design.cpu.reg_window\[8\] final_design.cpu.reg_window\[40\] net893
+ vssd1 vssd1 vccd1 vccd1 _02168_ sky130_fd_sc_hd__mux2_1
XANTENNA__13278__CLK clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout305_X net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08197_ final_design.cpu.reg_window\[846\] final_design.cpu.reg_window\[878\] net825
+ vssd1 vssd1 vccd1 vccd1 _03148_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07148_ net538 _02098_ vssd1 vssd1 vccd1 vccd1 _02099_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout886_A _01437_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07079_ _01851_ _02029_ _01821_ vssd1 vssd1 vccd1 vccd1 _02030_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_30_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10090_ _05004_ _05005_ vssd1 vssd1 vccd1 vccd1 _05006_ sky130_fd_sc_hd__nor2_1
Xfanout1007 _05171_ vssd1 vssd1 vccd1 vccd1 net1007 sky130_fd_sc_hd__buf_2
Xfanout1018 final_design.CPU_instr_adr\[2\] vssd1 vssd1 vccd1 vccd1 net1018 sky130_fd_sc_hd__clkbuf_4
Xfanout1029 net1036 vssd1 vssd1 vccd1 vccd1 net1029 sky130_fd_sc_hd__buf_4
XANTENNA_fanout674_X net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09543__A1 net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11350__A1 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout841_X net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11753__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_39_clk clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_39_clk sky130_fd_sc_hd__clkbuf_8
X_13780_ clknet_leaf_9_clk _01011_ net1152 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[768\]
+ sky130_fd_sc_hd__dfrtp_1
X_10992_ net86 net1045 vssd1 vssd1 vccd1 vccd1 _05718_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_2_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10877__B net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12731_ _06368_ _06371_ vssd1 vssd1 vccd1 vccd1 _06372_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_70_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_1857 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12941__RESET_B net1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12662_ _06318_ net1466 net979 vssd1 vssd1 vccd1 vccd1 _01333_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14053__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14165__RESET_B net1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11613_ net239 net631 vssd1 vssd1 vccd1 vccd1 _06164_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_61_2279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12602__B2 final_design.data_from_mem\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12593_ net1528 net998 net984 final_design.data_from_mem\[11\] vssd1 vssd1 vccd1
+ vccd1 _01286_ sky130_fd_sc_hd__a22o_1
X_11544_ net226 net635 vssd1 vssd1 vccd1 vccd1 _06128_ sky130_fd_sc_hd__and2_1
XFILLER_0_80_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12881__Q final_design.data_from_mem\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11475_ net202 net639 vssd1 vssd1 vccd1 vccd1 _06108_ sky130_fd_sc_hd__and2_1
X_13214_ clknet_leaf_13_clk _00445_ net1089 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[202\]
+ sky130_fd_sc_hd__dfrtp_1
X_10426_ net1460 net1030 _05196_ net249 vssd1 vssd1 vccd1 vccd1 _00154_ sky130_fd_sc_hd__a22o_1
X_14194_ net1252 vssd1 vssd1 vccd1 vccd1 gpio_oeb[6] sky130_fd_sc_hd__buf_2
XANTENNA_input68_X net68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13145_ clknet_leaf_57_clk _00376_ net1142 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[133\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_1418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10357_ net30 net1023 net1007 final_design.data_from_mem\[6\] vssd1 vssd1 vccd1 vccd1
+ _00110_ sky130_fd_sc_hd__o22a_1
XFILLER_0_57_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08810__B _01788_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09194__A net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13076_ clknet_leaf_13_clk _00307_ net1089 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[64\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12669__B2 final_design.data_from_mem\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06691__S1 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10288_ _01487_ net725 _02094_ net654 vssd1 vssd1 vccd1 vccd1 final_design.cpu.Error
+ sky130_fd_sc_hd__and4_1
XFILLER_0_40_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_1330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12027_ net1891 net230 net396 vssd1 vssd1 vccd1 vccd1 _00755_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11341__A1 net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09922__A _04341_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07145__C _02095_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13978_ clknet_leaf_58_clk _01209_ net1121 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[966\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06757__S net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12929_ clknet_leaf_47_clk _00167_ net1198 vssd1 vssd1 vccd1 vccd1 net152 sky130_fd_sc_hd__dfrtp_1
XANTENNA__11644__A2 net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06450_ final_design.vga.v_current_state\[0\] final_design.vga.v_current_state\[1\]
+ vssd1 vssd1 vccd1 vccd1 _01404_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_44_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13420__CLK clknet_leaf_45_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11251__X _05953_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08120_ _03070_ vssd1 vssd1 vccd1 vccd1 _03071_ sky130_fd_sc_hd__inv_2
XANTENNA__06492__S net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14253__1307 vssd1 vssd1 vccd1 vccd1 _14253__1307/HI net1307 sky130_fd_sc_hd__conb_1
X_08051_ final_design.cpu.reg_window\[274\] final_design.cpu.reg_window\[306\] net844
+ vssd1 vssd1 vccd1 vccd1 _03002_ sky130_fd_sc_hd__mux2_1
XANTENNA__12357__B1 net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07002_ net757 _01952_ vssd1 vssd1 vccd1 vccd1 _01953_ sky130_fd_sc_hd__or2_1
XFILLER_0_12_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13570__CLK clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload37_A clknet_leaf_27_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11838__S net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07176__X _02127_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08953_ _03795_ _03892_ vssd1 vssd1 vccd1 vccd1 _03893_ sky130_fd_sc_hd__nor2_1
XANTENNA__10314__Y _05167_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07904_ final_design.cpu.reg_window\[791\] final_design.cpu.reg_window\[823\] net849
+ vssd1 vssd1 vccd1 vccd1 _02855_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09525__B2 net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08884_ _03660_ _03661_ vssd1 vssd1 vccd1 vccd1 _03831_ sky130_fd_sc_hd__and2b_1
XFILLER_0_47_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07835_ final_design.cpu.reg_window\[853\] final_design.cpu.reg_window\[885\] net858
+ vssd1 vssd1 vccd1 vccd1 _02786_ sky130_fd_sc_hd__mux2_1
XANTENNA__07631__S0 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09289__A0 _01566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07766_ _02713_ _02714_ _02715_ _02716_ net686 net704 vssd1 vssd1 vccd1 vccd1 _02717_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_75_1761 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14076__CLK clknet_leaf_15_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09505_ _04421_ _04423_ vssd1 vssd1 vccd1 vccd1 _04424_ sky130_fd_sc_hd__xor2_1
XFILLER_0_71_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06717_ net761 _01667_ vssd1 vssd1 vccd1 vccd1 _01668_ sky130_fd_sc_hd__or2_1
XFILLER_0_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07697_ _02644_ _02645_ _02646_ _02647_ net688 net705 vssd1 vssd1 vccd1 vccd1 _02648_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout634_A net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout255_X net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09436_ net321 _04354_ _04349_ _04347_ vssd1 vssd1 vccd1 vccd1 _04355_ sky130_fd_sc_hd__o211a_1
X_06648_ net743 _01598_ net665 vssd1 vssd1 vccd1 vccd1 _01599_ sky130_fd_sc_hd__a21oi_4
XANTENNA_fanout801_A net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_24_clk_X clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09367_ net730 _04280_ _04285_ vssd1 vssd1 vccd1 vccd1 _04286_ sky130_fd_sc_hd__nand3_1
XANTENNA_fanout422_X net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06579_ final_design.cpu.reg_window\[669\] final_design.cpu.reg_window\[701\] net949
+ vssd1 vssd1 vccd1 vccd1 _01530_ sky130_fd_sc_hd__mux2_1
XANTENNA__11399__A1 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12596__B1 net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09687__S1 net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08318_ final_design.cpu.reg_window\[72\] final_design.cpu.reg_window\[104\] net812
+ vssd1 vssd1 vccd1 vccd1 _03269_ sky130_fd_sc_hd__mux2_1
X_09298_ _04119_ _04215_ _04216_ _04212_ vssd1 vssd1 vccd1 vccd1 _04217_ sky130_fd_sc_hd__o211a_1
XFILLER_0_7_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13913__CLK clknet_leaf_54_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08249_ _02128_ net599 vssd1 vssd1 vccd1 vccd1 _03200_ sky130_fd_sc_hd__nand2_1
XFILLER_0_82_1721 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12348__B1 net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_39_clk_X clknet_leaf_39_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11260_ net663 _03938_ net736 vssd1 vssd1 vccd1 vccd1 _05961_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout791_X net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10211_ _05094_ _05095_ net799 vssd1 vssd1 vccd1 vccd1 _00031_ sky130_fd_sc_hd__and3b_1
XANTENNA__11748__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11191_ net732 _04002_ _05899_ vssd1 vssd1 vccd1 vccd1 _05900_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_54_2050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10374__A2 net1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_2684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11571__A1 net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_2061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10142_ net1050 final_design.VGA_data_control.h_count\[3\] net1049 final_design.VGA_data_control.h_count\[4\]
+ vssd1 vssd1 vccd1 vccd1 _05043_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_73_2695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08122__S net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06673__S1 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13140__RESET_B net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10073_ _01481_ net725 net251 vssd1 vssd1 vccd1 vccd1 _04991_ sky130_fd_sc_hd__or3_2
XANTENNA__12520__B1 net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13901_ clknet_leaf_44_clk _01132_ net1205 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[889\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input28_A DAT_I[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11874__A2 net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11336__X _06028_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11369__A2_N _05947_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13832_ clknet_leaf_41_clk _01063_ net1224 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[820\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12876__Q final_design.data_from_mem\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_2488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13763_ clknet_leaf_1_clk _00994_ net1062 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[751\]
+ sky130_fd_sc_hd__dfrtp_1
X_10975_ _05679_ _05681_ _05699_ _05700_ vssd1 vssd1 vccd1 vccd1 _05702_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_67_2499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10400__B _05181_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13443__CLK clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12714_ final_design.VGA_data_control.v_count\[2\] _06354_ vssd1 vssd1 vccd1 vccd1
+ _06355_ sky130_fd_sc_hd__or2_1
XFILLER_0_54_1889 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06502__A1 net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11215__C net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13694_ clknet_leaf_11_clk _00925_ net1087 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[682\]
+ sky130_fd_sc_hd__dfrtp_1
X_12645_ final_design.VGA_data_control.ready_data\[10\] net1019 net974 final_design.data_from_mem\[10\]
+ vssd1 vssd1 vccd1 vccd1 _06310_ sky130_fd_sc_hd__a22o_1
XANTENNA__12587__B1 net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08805__B _01722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12576_ net1052 final_design.uart.working_data\[8\] vssd1 vssd1 vccd1 vccd1 _06293_
+ sky130_fd_sc_hd__and2_1
XANTENNA__13593__CLK clknet_leaf_52_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11527_ net2286 net192 net523 vssd1 vssd1 vccd1 vccd1 _00394_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12339__B1 net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14246_ net1300 vssd1 vssd1 vccd1 vccd1 gpio_out[24] sky130_fd_sc_hd__buf_2
Xhold309 final_design.VGA_data_control.ready_data\[17\] vssd1 vssd1 vccd1 vccd1 net1651
+ sky130_fd_sc_hd__dlygate4sd3_1
X_11458_ net244 net638 vssd1 vssd1 vccd1 vccd1 _06102_ sky130_fd_sc_hd__and2_1
XFILLER_0_7_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10409_ net1500 net1030 _05187_ net246 vssd1 vssd1 vccd1 vccd1 _00146_ sky130_fd_sc_hd__a22o_1
XFILLER_0_46_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14177_ clknet_leaf_21_clk _01351_ net1161 vssd1 vssd1 vccd1 vccd1 final_design.VGA_adr\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11389_ net649 net180 vssd1 vssd1 vccd1 vccd1 _06075_ sky130_fd_sc_hd__and2_1
XANTENNA__10365__A2 net1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07437__A net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1248 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13128_ clknet_leaf_35_clk _00359_ net1240 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[116\]
+ sky130_fd_sc_hd__dfrtp_1
X_13059_ clknet_leaf_0_clk _00290_ net1062 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[47\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1009 final_design.cpu.reg_window\[104\] vssd1 vssd1 vccd1 vccd1 net2351 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11314__A1 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14099__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12511__B1 net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07620_ _01539_ net616 vssd1 vssd1 vccd1 vccd1 _02571_ sky130_fd_sc_hd__nor2_1
XFILLER_0_72_1901 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07551_ net885 _02495_ _02501_ _02488_ _02489_ vssd1 vssd1 vccd1 vccd1 _02502_ sky130_fd_sc_hd__a32oi_4
X_06502_ net885 _01445_ _01451_ _01439_ _01436_ vssd1 vssd1 vccd1 vccd1 _01453_ sky130_fd_sc_hd__a32o_2
XFILLER_0_75_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07482_ _02332_ _02431_ _02331_ vssd1 vssd1 vccd1 vccd1 _02433_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_5_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09221_ _02126_ _03195_ _03226_ _03197_ vssd1 vssd1 vccd1 vccd1 _04140_ sky130_fd_sc_hd__o31ai_2
X_06433_ net57 vssd1 vssd1 vccd1 vccd1 _01388_ sky130_fd_sc_hd__inv_2
XANTENNA__13936__CLK clknet_leaf_34_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08715__B _01660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09152_ _03645_ _03651_ net450 vssd1 vssd1 vccd1 vccd1 _04071_ sky130_fd_sc_hd__a21oi_2
XANTENNA__07049__A2 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10053__A1 _04954_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08103_ final_design.cpu.reg_window\[844\] final_design.cpu.reg_window\[876\] net825
+ vssd1 vssd1 vccd1 vccd1 _03054_ sky130_fd_sc_hd__mux2_1
XANTENNA__10053__B2 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09994__A1 net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11250__B1 net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09083_ final_design.CPU_instr_adr\[5\] _03784_ vssd1 vssd1 vccd1 vccd1 _04008_ sky130_fd_sc_hd__nor2_1
XANTENNA__10038__A _04954_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout215_A _05941_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08034_ final_design.cpu.reg_window\[723\] final_design.cpu.reg_window\[755\] net830
+ vssd1 vssd1 vccd1 vccd1 _02985_ sky130_fd_sc_hd__mux2_1
Xinput70 memory_size[11] vssd1 vssd1 vccd1 vccd1 net70 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput81 memory_size[21] vssd1 vssd1 vccd1 vccd1 net81 sky130_fd_sc_hd__buf_1
Xhold810 final_design.cpu.reg_window\[997\] vssd1 vssd1 vccd1 vccd1 net2152 sky130_fd_sc_hd__dlygate4sd3_1
Xhold821 final_design.cpu.reg_window\[516\] vssd1 vssd1 vccd1 vccd1 net2163 sky130_fd_sc_hd__dlygate4sd3_1
Xinput92 memory_size[31] vssd1 vssd1 vccd1 vccd1 net92 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold832 final_design.cpu.reg_window\[790\] vssd1 vssd1 vccd1 vccd1 net2174 sky130_fd_sc_hd__dlygate4sd3_1
Xhold843 final_design.cpu.reg_window\[35\] vssd1 vssd1 vccd1 vccd1 net2185 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09546__B _04368_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold854 final_design.cpu.reg_window\[988\] vssd1 vssd1 vccd1 vccd1 net2196 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold865 final_design.cpu.reg_window\[324\] vssd1 vssd1 vccd1 vccd1 net2207 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1124_A net1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold876 final_design.cpu.reg_window\[123\] vssd1 vssd1 vccd1 vccd1 net2218 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11553__B2 net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold887 final_design.cpu.reg_window\[661\] vssd1 vssd1 vccd1 vccd1 net2229 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07347__A _02294_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_51_clk_A clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold898 final_design.cpu.reg_window\[303\] vssd1 vssd1 vccd1 vccd1 net2240 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13316__CLK clknet_leaf_52_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06655__S1 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09985_ net728 _04898_ _04901_ vssd1 vssd1 vccd1 vccd1 _04904_ sky130_fd_sc_hd__and3_1
XFILLER_0_60_1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout584_A net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08936_ _03796_ _03877_ vssd1 vssd1 vccd1 vccd1 _03878_ sky130_fd_sc_hd__or2_1
XANTENNA__12502__B1 net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08867_ _01540_ _01541_ vssd1 vssd1 vccd1 vccd1 _03816_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout751_A net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout372_X net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_66_clk_A clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13466__CLK clknet_leaf_58_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07818_ _02766_ _02767_ vssd1 vssd1 vccd1 vccd1 _02769_ sky130_fd_sc_hd__nor2_2
XFILLER_0_58_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08798_ _03677_ _03678_ _03747_ vssd1 vssd1 vccd1 vccd1 _03749_ sky130_fd_sc_hd__nor3_1
XANTENNA__07082__A _02026_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11608__A2 net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07749_ net604 _02698_ _02674_ vssd1 vssd1 vccd1 vccd1 _02700_ sky130_fd_sc_hd__o21a_1
XANTENNA__11316__B net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout637_X net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10760_ net42 _05483_ _05493_ _05495_ vssd1 vssd1 vccd1 vccd1 _05497_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_62_2330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_2964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_2341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_2975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1805 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_2986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09419_ _04336_ _04337_ net472 vssd1 vssd1 vccd1 vccd1 _04338_ sky130_fd_sc_hd__mux2_1
X_10691_ _01365_ _03957_ net1058 vssd1 vssd1 vccd1 vccd1 _05431_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_1849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11332__A net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12430_ net177 net640 net354 _06281_ vssd1 vssd1 vccd1 vccd1 _01138_ sky130_fd_sc_hd__a31o_1
XFILLER_0_35_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06426__A final_design.data_from_mem\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07021__S net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12361_ net2239 net362 net353 _06082_ vssd1 vssd1 vccd1 vccd1 _01073_ sky130_fd_sc_hd__a22o_1
XANTENNA__11241__B1 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06799__A1 net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_2893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14100_ clknet_leaf_9_clk _01297_ net1104 vssd1 vssd1 vccd1 vccd1 final_design.reqhand.instruction\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_11312_ final_design.data_from_mem\[20\] net236 net234 vssd1 vssd1 vccd1 vccd1 _06007_
+ sky130_fd_sc_hd__a21o_2
XTAP_TAPCELL_ROW_56_2112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_2123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12292_ net584 _06222_ net512 net370 net2175 vssd1 vssd1 vccd1 vccd1 _01007_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_75_2757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_2134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_2768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_2779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14031_ clknet_leaf_42_clk _01262_ net1223 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[1019\]
+ sky130_fd_sc_hd__dfrtp_1
X_11243_ net741 _01481_ vssd1 vssd1 vccd1 vccd1 _05946_ sky130_fd_sc_hd__nor2_2
XANTENNA_clkbuf_leaf_19_clk_A clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11174_ net662 _04014_ net735 vssd1 vssd1 vccd1 vccd1 _05885_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_60_1871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10125_ final_design.VGA_data_control.v_count\[8\] _05017_ _05032_ vssd1 vssd1 vccd1
+ vccd1 _05033_ sky130_fd_sc_hd__mux2_1
XANTENNA__13809__CLK clknet_leaf_34_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08399__S1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10056_ _04970_ _04972_ _04973_ _04974_ vssd1 vssd1 vccd1 vccd1 _04975_ sky130_fd_sc_hd__or4_1
XANTENNA__11847__A2 net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14252__1306 vssd1 vssd1 vccd1 vccd1 _14252__1306/HI net1306 sky130_fd_sc_hd__conb_1
XFILLER_0_76_1344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12102__S net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06723__A1 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13959__CLK clknet_leaf_61_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13815_ clknet_leaf_58_clk _01046_ net1132 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[803\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13746_ clknet_leaf_39_clk _00977_ net1205 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[734\]
+ sky130_fd_sc_hd__dfrtp_1
X_10958_ net967 _05685_ vssd1 vssd1 vccd1 vccd1 _05686_ sky130_fd_sc_hd__nand2_1
XFILLER_0_70_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08020__S0 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11480__A0 _06017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_1096 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13677_ clknet_leaf_48_clk _00908_ net1186 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[665\]
+ sky130_fd_sc_hd__dfrtp_1
X_10889_ net669 _05608_ _05619_ net966 _05618_ vssd1 vssd1 vccd1 vccd1 _05620_ sky130_fd_sc_hd__o221a_1
XANTENNA__06582__S0 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11242__A net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12628_ _06301_ net1448 net980 vssd1 vssd1 vccd1 vccd1 _01316_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_14_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_1394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_14_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12559_ _06222_ net357 net324 net2450 vssd1 vssd1 vccd1 vccd1 _01263_ sky130_fd_sc_hd__a22o_1
XFILLER_0_48_1435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold106 final_design.VGA_data_control.data_to_VGA\[1\] vssd1 vssd1 vccd1 vccd1 net1448
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06885__S1 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold117 net147 vssd1 vssd1 vccd1 vccd1 net1459 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_9_Right_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold128 net112 vssd1 vssd1 vccd1 vccd1 net1470 sky130_fd_sc_hd__dlygate4sd3_1
X_14229_ net1283 vssd1 vssd1 vccd1 vccd1 gpio_out[7] sky130_fd_sc_hd__buf_2
Xhold139 final_design.VGA_data_control.data_to_VGA\[27\] vssd1 vssd1 vccd1 vccd1 net1481
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_65_1793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11535__A1 net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout608 net609 vssd1 vssd1 vccd1 vccd1 net608 sky130_fd_sc_hd__buf_2
XANTENNA__06637__S1 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout619 net620 vssd1 vssd1 vccd1 vccd1 net619 sky130_fd_sc_hd__buf_2
XFILLER_0_42_1067 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13489__CLK clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09770_ _03590_ net446 _04687_ _04688_ net261 vssd1 vssd1 vccd1 vccd1 _04689_ sky130_fd_sc_hd__o2111a_1
X_06982_ final_design.cpu.reg_window\[592\] final_design.cpu.reg_window\[624\] net923
+ vssd1 vssd1 vccd1 vccd1 _01933_ sky130_fd_sc_hd__mux2_1
X_08721_ final_design.CPU_instr_adr\[19\] _01853_ vssd1 vssd1 vccd1 vccd1 _03672_
+ sky130_fd_sc_hd__nand2_1
XANTENNA__07454__X _02405_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11299__B1 net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1190 net1191 vssd1 vssd1 vccd1 vccd1 net1190 sky130_fd_sc_hd__clkbuf_4
X_08652_ _02706_ _03600_ _03602_ _02673_ _03601_ vssd1 vssd1 vccd1 vccd1 _03603_ sky130_fd_sc_hd__a221o_1
XANTENNA__07062__S1 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07603_ final_design.cpu.reg_window\[221\] final_design.cpu.reg_window\[253\] net870
+ vssd1 vssd1 vccd1 vccd1 _02554_ sky130_fd_sc_hd__mux2_1
X_08583_ _03530_ _03531_ _03532_ _03533_ net675 net697 vssd1 vssd1 vccd1 vccd1 _03534_
+ sky130_fd_sc_hd__mux4_2
X_07534_ final_design.cpu.reg_window\[223\] final_design.cpu.reg_window\[255\] net937
+ vssd1 vssd1 vccd1 vccd1 _02485_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09664__B1 _04117_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_14_Left_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07465_ final_design.cpu.reg_window\[512\] final_design.cpu.reg_window\[544\] net906
+ vssd1 vssd1 vccd1 vccd1 _02416_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout332_A net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14114__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09204_ net487 _04077_ _04117_ _04122_ _04068_ vssd1 vssd1 vccd1 vccd1 _04123_ sky130_fd_sc_hd__o311a_1
X_06416_ net1053 vssd1 vssd1 vccd1 vccd1 _01371_ sky130_fd_sc_hd__inv_2
XANTENNA__12015__A2 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07396_ final_design.cpu.reg_window\[834\] final_design.cpu.reg_window\[866\] net913
+ vssd1 vssd1 vccd1 vccd1 _02347_ sky130_fd_sc_hd__mux2_1
XANTENNA__09416__B1 _04234_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10026__A1 net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10026__B2 net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09135_ _03629_ _04053_ vssd1 vssd1 vccd1 vccd1 _04054_ sky130_fd_sc_hd__nor2_2
XANTENNA__12682__S net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1241_A net1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07776__S net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11386__A1_N net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09066_ net622 _03992_ vssd1 vssd1 vccd1 vccd1 _03993_ sky130_fd_sc_hd__nor2_1
XFILLER_0_4_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08017_ final_design.cpu.reg_window\[275\] final_design.cpu.reg_window\[307\] net830
+ vssd1 vssd1 vccd1 vccd1 _02968_ sky130_fd_sc_hd__mux2_1
Xhold640 final_design.cpu.reg_window\[743\] vssd1 vssd1 vccd1 vccd1 net1982 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10329__A2 net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold651 final_design.cpu.reg_window\[694\] vssd1 vssd1 vccd1 vccd1 net1993 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08180__B net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_2610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold662 final_design.cpu.reg_window\[339\] vssd1 vssd1 vccd1 vccd1 net2004 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1127_X net1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold673 final_design.cpu.reg_window\[889\] vssd1 vssd1 vccd1 vccd1 net2015 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09195__A2 net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold684 final_design.cpu.reg_window\[738\] vssd1 vssd1 vccd1 vccd1 net2026 sky130_fd_sc_hd__dlygate4sd3_1
Xhold695 final_design.cpu.reg_window\[944\] vssd1 vssd1 vccd1 vccd1 net2037 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout966_A net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout587_X net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09968_ _04180_ _04886_ vssd1 vssd1 vccd1 vccd1 _04887_ sky130_fd_sc_hd__or2_1
XANTENNA__10930__S net1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12856__CLK clknet_leaf_17_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08919_ _03758_ _03861_ vssd1 vssd1 vccd1 vccd1 _03862_ sky130_fd_sc_hd__and2_1
XANTENNA__08400__S net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09899_ net490 _04664_ vssd1 vssd1 vccd1 vccd1 _04818_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout754_X net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11930_ net555 net244 net634 vssd1 vssd1 vccd1 vccd1 _06254_ sky130_fd_sc_hd__and3_1
XANTENNA__10501__A2 _04825_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_2403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11861_ net427 _05965_ net553 net517 net1775 vssd1 vssd1 vccd1 vccd1 _00609_ sky130_fd_sc_hd__a32o_1
XFILLER_0_68_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1913 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11761__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13600_ clknet_leaf_11_clk _00831_ net1086 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[588\]
+ sky130_fd_sc_hd__dfrtp_1
X_10812_ _04452_ net252 vssd1 vssd1 vccd1 vccd1 _05546_ sky130_fd_sc_hd__nor2_1
XFILLER_0_39_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06708__X _01659_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11792_ net2455 net414 net285 _05990_ vssd1 vssd1 vccd1 vccd1 _00548_ sky130_fd_sc_hd__a22o_1
XANTENNA__06855__S net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13531_ clknet_leaf_66_clk _00762_ net1063 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[519\]
+ sky130_fd_sc_hd__dfrtp_1
X_10743_ _05478_ _05480_ vssd1 vssd1 vccd1 vccd1 _05481_ sky130_fd_sc_hd__and2_1
XFILLER_0_32_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06564__S0 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13462_ clknet_leaf_59_clk _00693_ net1139 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[450\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input95_A memory_size[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10674_ final_design.CPU_instr_adr\[11\] _03965_ net1058 vssd1 vssd1 vccd1 vccd1
+ _05415_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_11_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_2819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12413_ _06242_ net501 net339 net1924 vssd1 vssd1 vccd1 vccd1 _01123_ sky130_fd_sc_hd__a22o_1
XFILLER_0_36_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13393_ clknet_leaf_35_clk _00624_ net1241 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[381\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12344_ net2278 net363 net353 _05959_ vssd1 vssd1 vccd1 vccd1 _01056_ sky130_fd_sc_hd__a22o_1
XFILLER_0_49_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08069__S0 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12275_ net568 _06205_ net506 net368 net1970 vssd1 vssd1 vccd1 vccd1 _00990_ sky130_fd_sc_hd__a32o_1
XANTENNA__10406__A _03415_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08090__B net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13631__CLK clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1332 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14014_ clknet_leaf_13_clk _01245_ net1099 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[1002\]
+ sky130_fd_sc_hd__dfrtp_1
X_11226_ net660 _03971_ net732 vssd1 vssd1 vccd1 vccd1 _05931_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_23_1917 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12190__A1 net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10840__S net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11157_ net662 _04025_ net734 vssd1 vssd1 vccd1 vccd1 _05870_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_65_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10108_ final_design.VGA_data_control.v_count\[2\] _05019_ _05006_ vssd1 vssd1 vccd1
+ vccd1 _05022_ sky130_fd_sc_hd__o21ai_1
X_11088_ net966 _05809_ vssd1 vssd1 vccd1 vccd1 _05810_ sky130_fd_sc_hd__nand2_1
XANTENNA__13781__CLK clknet_leaf_57_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11237__A net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10039_ _04614_ _04615_ _04941_ _04942_ _04957_ vssd1 vssd1 vccd1 vccd1 _04958_ sky130_fd_sc_hd__o2111a_1
XANTENNA__12493__A2 net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14137__CLK clknet_leaf_17_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11243__Y _05946_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13729_ clknet_leaf_47_clk _00960_ net1198 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[717\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07250_ final_design.cpu.reg_window\[775\] final_design.cpu.reg_window\[807\] net892
+ vssd1 vssd1 vccd1 vccd1 _02201_ sky130_fd_sc_hd__mux2_1
XANTENNA__11403__C _06086_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13161__CLK clknet_leaf_36_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07181_ final_design.cpu.reg_window\[265\] final_design.cpu.reg_window\[297\] net891
+ vssd1 vssd1 vccd1 vccd1 _02132_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_41_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1276 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06632__B1 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12879__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout405 _06255_ vssd1 vssd1 vccd1 vccd1 net405 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_6_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout416 net417 vssd1 vssd1 vccd1 vccd1 net416 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_6_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout427 net431 vssd1 vssd1 vccd1 vccd1 net427 sky130_fd_sc_hd__clkbuf_4
X_09822_ _03293_ _04153_ _04154_ vssd1 vssd1 vccd1 vccd1 _04741_ sky130_fd_sc_hd__and3_1
XFILLER_0_22_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout438 _04095_ vssd1 vssd1 vccd1 vccd1 net438 sky130_fd_sc_hd__buf_4
XANTENNA__08480__S0 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout449 _04070_ vssd1 vssd1 vccd1 vccd1 net449 sky130_fd_sc_hd__buf_4
X_09753_ _04660_ _04661_ _04671_ vssd1 vssd1 vccd1 vccd1 _04672_ sky130_fd_sc_hd__a21oi_1
X_06965_ final_design.cpu.reg_window\[400\] final_design.cpu.reg_window\[432\] net926
+ vssd1 vssd1 vccd1 vccd1 _01916_ sky130_fd_sc_hd__mux2_1
XANTENNA__08220__S net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout282_A net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08704_ net256 vssd1 vssd1 vccd1 vccd1 _03655_ sky130_fd_sc_hd__clkinv_4
X_09684_ _04097_ _04205_ _04229_ vssd1 vssd1 vccd1 vccd1 _04603_ sky130_fd_sc_hd__o21ai_1
XANTENNA__12484__A2 net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06896_ final_design.cpu.reg_window\[531\] final_design.cpu.reg_window\[563\] net903
+ vssd1 vssd1 vccd1 vccd1 _01847_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08635_ net603 _02961_ _02962_ _01938_ vssd1 vssd1 vccd1 vccd1 _03586_ sky130_fd_sc_hd__o211a_1
XANTENNA__11692__B1 net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10986__A net1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1191_A net1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout547_A _01880_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1269 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08566_ _02394_ net595 vssd1 vssd1 vccd1 vccd1 _03517_ sky130_fd_sc_hd__nand2_1
XANTENNA__12974__Q final_design.reqhand.current_client\[3\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__07360__A net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13504__CLK clknet_leaf_11_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07517_ _01725_ _02465_ _01692_ _01724_ vssd1 vssd1 vccd1 vccd1 _02468_ sky130_fd_sc_hd__a211o_1
XFILLER_0_65_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08497_ _03444_ _03445_ _03446_ _03447_ net678 net692 vssd1 vssd1 vccd1 vccd1 _03448_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__07112__A1 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout714_A net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout335_X net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07112__B2 _02061_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07448_ final_design.cpu.reg_window\[384\] final_design.cpu.reg_window\[416\] net907
+ vssd1 vssd1 vccd1 vccd1 _02399_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_21_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout502_X net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07379_ _01496_ net710 net672 _01484_ vssd1 vssd1 vccd1 vccd1 _02330_ sky130_fd_sc_hd__a2bb2o_2
XANTENNA_fanout1244_X net1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13654__CLK clknet_leaf_61_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09118_ net1053 final_design.reqhand.current_client\[1\] vssd1 vssd1 vccd1 vccd1
+ _04037_ sky130_fd_sc_hd__or2_1
XFILLER_0_44_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09287__A net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14251__1305 vssd1 vssd1 vccd1 vccd1 _14251__1305/HI net1305 sky130_fd_sc_hd__conb_1
X_10390_ _02028_ _03624_ _03613_ vssd1 vssd1 vccd1 vccd1 _05176_ sky130_fd_sc_hd__o21a_1
XANTENNA__07078__Y _02029_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09049_ _02158_ _02159_ vssd1 vssd1 vccd1 vccd1 _03978_ sky130_fd_sc_hd__or2_1
XFILLER_0_60_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12966__RESET_B net1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12060_ net671 _05850_ _06262_ vssd1 vssd1 vccd1 vccd1 _06263_ sky130_fd_sc_hd__or3_4
Xhold470 final_design.uart.BAUD_counter\[25\] vssd1 vssd1 vccd1 vccd1 net1812 sky130_fd_sc_hd__dlygate4sd3_1
Xhold481 final_design.cpu.reg_window\[695\] vssd1 vssd1 vccd1 vccd1 net1823 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout871_X net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12172__A1 net221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11011_ net87 net1045 vssd1 vssd1 vccd1 vccd1 _05736_ sky130_fd_sc_hd__and2_1
Xhold492 final_design.cpu.reg_window\[983\] vssd1 vssd1 vccd1 vccd1 net1834 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11756__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11380__C1 net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout950 net951 vssd1 vssd1 vccd1 vccd1 net950 sky130_fd_sc_hd__buf_4
Xfanout961 _04036_ vssd1 vssd1 vccd1 vccd1 net961 sky130_fd_sc_hd__clkbuf_4
Xfanout972 _01415_ vssd1 vssd1 vccd1 vccd1 net972 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout983 net985 vssd1 vssd1 vccd1 vccd1 net983 sky130_fd_sc_hd__clkbuf_4
Xfanout994 _01408_ vssd1 vssd1 vccd1 vccd1 net994 sky130_fd_sc_hd__clkbuf_2
XANTENNA__13034__CLK clknet_leaf_60_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12962_ clknet_leaf_32_clk _00200_ net1234 vssd1 vssd1 vccd1 vccd1 net120 sky130_fd_sc_hd__dfrtp_1
XANTENNA__12475__A2 net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1170 final_design.cpu.reg_window\[843\] vssd1 vssd1 vccd1 vccd1 net2512 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_input10_A DAT_I[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11913_ net187 net2274 net274 vssd1 vssd1 vccd1 vccd1 _00653_ sky130_fd_sc_hd__mux2_1
Xhold1181 final_design.cpu.reg_window\[942\] vssd1 vssd1 vccd1 vccd1 net2523 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1192 final_design.cpu.reg_window\[806\] vssd1 vssd1 vccd1 vccd1 net2534 sky130_fd_sc_hd__dlygate4sd3_1
X_12893_ clknet_leaf_17_clk _00131_ net1113 vssd1 vssd1 vccd1 vccd1 final_design.data_from_mem\[27\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__11491__S net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06785__S0 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11344__X _06035_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11844_ net804 _05842_ net553 vssd1 vssd1 vccd1 vccd1 _06239_ sky130_fd_sc_hd__or3b_1
XFILLER_0_9_1899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07270__A net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12884__Q final_design.data_from_mem\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09723__S0 net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11775_ net2415 net413 _06230_ net428 vssd1 vssd1 vccd1 vccd1 _00534_ sky130_fd_sc_hd__a22o_1
XFILLER_0_51_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10726_ _05427_ _05449_ _05463_ _05447_ vssd1 vssd1 vccd1 vccd1 _05464_ sky130_fd_sc_hd__o211a_1
X_13514_ clknet_leaf_60_clk _00745_ net1143 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[502\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07654__A2 _02602_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13445_ clknet_leaf_48_clk _00676_ net1182 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[433\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_64_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10657_ net668 _05388_ _05398_ net964 _05397_ vssd1 vssd1 vccd1 vccd1 _05399_ sky130_fd_sc_hd__o221a_1
Xclkload15 clknet_leaf_15_clk vssd1 vssd1 vccd1 vccd1 clkload15/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_24_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09197__A net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload26 clknet_leaf_26_clk vssd1 vssd1 vccd1 vccd1 clkload26/Y sky130_fd_sc_hd__inv_16
Xclkload37 clknet_leaf_27_clk vssd1 vssd1 vccd1 vccd1 clkload37/Y sky130_fd_sc_hd__clkinv_8
XFILLER_0_3_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13376_ clknet_leaf_10_clk _00607_ net1101 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[364\]
+ sky130_fd_sc_hd__dfrtp_1
X_10588_ _05331_ _05332_ vssd1 vssd1 vccd1 vccd1 _05333_ sky130_fd_sc_hd__nand2_1
XANTENNA__06614__A net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12327_ net1892 net179 net366 vssd1 vssd1 vccd1 vccd1 _01041_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09159__A2 _03550_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12258_ net581 _06187_ net514 net374 net1550 vssd1 vssd1 vccd1 vccd1 _00974_ sky130_fd_sc_hd__a32o_1
X_11209_ net735 _03987_ _05915_ vssd1 vssd1 vccd1 vccd1 _05916_ sky130_fd_sc_hd__a21oi_2
X_12189_ net1710 net188 net382 vssd1 vssd1 vccd1 vccd1 _00908_ sky130_fd_sc_hd__mux2_1
XANTENNA__08462__S0 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1195 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06917__A1 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_34_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06750_ final_design.cpu.reg_window\[151\] final_design.cpu.reg_window\[183\] net929
+ vssd1 vssd1 vccd1 vccd1 _01701_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_82_3001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_3012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12466__A2 net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_3023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_3034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13527__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_3045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11674__B1 net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06681_ _01627_ _01630_ vssd1 vssd1 vccd1 vccd1 _01632_ sky130_fd_sc_hd__or2_1
XFILLER_0_25_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08420_ net718 _03370_ vssd1 vssd1 vccd1 vccd1 _03371_ sky130_fd_sc_hd__or2_1
XFILLER_0_8_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08351_ _03298_ _03299_ _03300_ _03301_ net676 net696 vssd1 vssd1 vccd1 vccd1 _03302_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_28_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13677__CLK clknet_leaf_48_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07302_ _02249_ _02250_ _02251_ _02252_ net770 net789 vssd1 vssd1 vccd1 vccd1 _02253_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_28_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_1917 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08282_ final_design.cpu.reg_window\[329\] final_design.cpu.reg_window\[361\] net820
+ vssd1 vssd1 vccd1 vccd1 _03233_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_24_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload9 clknet_leaf_56_clk vssd1 vssd1 vccd1 vccd1 clkload9/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_50_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07233_ net881 _02177_ _02183_ _02170_ _02171_ vssd1 vssd1 vccd1 vccd1 _02184_ sky130_fd_sc_hd__a32oi_4
XFILLER_0_70_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07164_ final_design.cpu.reg_window\[778\] final_design.cpu.reg_window\[810\] net898
+ vssd1 vssd1 vccd1 vccd1 _02115_ sky130_fd_sc_hd__mux2_1
XFILLER_0_41_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10401__B2 net246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07095_ final_design.cpu.reg_window\[844\] final_design.cpu.reg_window\[876\] net906
+ vssd1 vssd1 vccd1 vccd1 _02046_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout1037_A _01410_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08358__B1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout202 _05996_ vssd1 vssd1 vccd1 vccd1 net202 sky130_fd_sc_hd__clkbuf_2
XANTENNA__13057__CLK clknet_leaf_49_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout497_A _03418_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09555__C1 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout213 _05951_ vssd1 vssd1 vccd1 vccd1 net213 sky130_fd_sc_hd__clkbuf_2
Xfanout224 _05897_ vssd1 vssd1 vccd1 vccd1 net224 sky130_fd_sc_hd__buf_2
XANTENNA_fanout1204_A net1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout235 _05982_ vssd1 vssd1 vccd1 vccd1 net235 sky130_fd_sc_hd__buf_2
Xfanout246 net247 vssd1 vssd1 vccd1 vccd1 net246 sky130_fd_sc_hd__buf_4
X_09805_ net728 _04723_ vssd1 vssd1 vccd1 vccd1 _04724_ sky130_fd_sc_hd__nand2_1
Xfanout257 net258 vssd1 vssd1 vccd1 vccd1 net257 sky130_fd_sc_hd__buf_2
XANTENNA_input2_A DAT_I[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09570__A2 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11148__Y _05862_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout268 net269 vssd1 vssd1 vccd1 vccd1 net268 sky130_fd_sc_hd__buf_4
X_07997_ net721 _02947_ vssd1 vssd1 vccd1 vccd1 _02948_ sky130_fd_sc_hd__or2_1
Xfanout279 net284 vssd1 vssd1 vccd1 vccd1 net279 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout285_X net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09736_ net71 _04183_ vssd1 vssd1 vccd1 vccd1 _04655_ sky130_fd_sc_hd__nand2_1
X_06948_ final_design.cpu.reg_window\[977\] final_design.cpu.reg_window\[1009\] net928
+ vssd1 vssd1 vccd1 vccd1 _01899_ sky130_fd_sc_hd__mux2_1
XANTENNA__07008__S1 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10468__A1 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09322__A2 _04240_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09667_ net486 _04578_ _04579_ _04585_ vssd1 vssd1 vccd1 vccd1 _04586_ sky130_fd_sc_hd__a31o_1
X_06879_ _01826_ _01827_ _01828_ _01829_ net769 net790 vssd1 vssd1 vccd1 vccd1 _01830_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout831_A net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout929_A net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08618_ _03426_ _03561_ _03567_ vssd1 vssd1 vccd1 vccd1 _03569_ sky130_fd_sc_hd__a21o_1
XFILLER_0_74_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09598_ _04097_ _04437_ vssd1 vssd1 vccd1 vccd1 _04517_ sky130_fd_sc_hd__or2_1
XANTENNA__07884__A2 _02830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08549_ net710 _03493_ net722 vssd1 vssd1 vccd1 vccd1 _03500_ sky130_fd_sc_hd__o21a_1
XANTENNA__11324__B net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout717_X net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11560_ net214 net635 vssd1 vssd1 vccd1 vccd1 _06136_ sky130_fd_sc_hd__and2_2
XANTENNA__12090__B1 net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10511_ net961 _05259_ vssd1 vssd1 vccd1 vccd1 _05260_ sky130_fd_sc_hd__or2_1
XFILLER_0_0_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11491_ net182 net2519 net309 vssd1 vssd1 vccd1 vccd1 _00367_ sky130_fd_sc_hd__mux2_1
XANTENNA__11340__A net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13230_ clknet_leaf_43_clk _00461_ net1218 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[218\]
+ sky130_fd_sc_hd__dfrtp_1
X_10442_ _02797_ net592 vssd1 vssd1 vccd1 vccd1 _05205_ sky130_fd_sc_hd__nor2_1
XFILLER_0_32_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13161_ clknet_leaf_36_clk _00392_ net1228 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[149\]
+ sky130_fd_sc_hd__dfrtp_1
X_10373_ net16 net1024 net1006 final_design.data_from_mem\[22\] vssd1 vssd1 vccd1
+ vccd1 _00126_ sky130_fd_sc_hd__o22a_1
XFILLER_0_81_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12112_ net1669 net203 net391 vssd1 vssd1 vccd1 vccd1 _00836_ sky130_fd_sc_hd__mux2_1
XANTENNA_input58_A mem_adr_start[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13092_ clknet_leaf_53_clk _00323_ net1187 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[80\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_44_1460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12043_ net1564 net222 net399 vssd1 vssd1 vccd1 vccd1 _00771_ sky130_fd_sc_hd__mux2_1
XANTENNA__11339__X _06031_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07247__S1 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11353__C1 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12879__Q final_design.data_from_mem\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout780 net782 vssd1 vssd1 vccd1 vccd1 net780 sky130_fd_sc_hd__clkbuf_4
Xfanout791 net795 vssd1 vssd1 vccd1 vccd1 net791 sky130_fd_sc_hd__buf_4
X_13994_ clknet_leaf_60_clk _01225_ net1142 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[982\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07552__X _02503_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input13_X net13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09313__A2 net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10459__B2 net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11656__B1 net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12945_ clknet_leaf_29_clk _00183_ net1193 vssd1 vssd1 vccd1 vccd1 net102 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06758__S0 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12110__S net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_49 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12876_ clknet_leaf_19_clk _00114_ net1111 vssd1 vssd1 vccd1 vccd1 final_design.data_from_mem\[10\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_51_1420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09077__A1 net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11827_ net222 net1932 net265 vssd1 vssd1 vccd1 vccd1 _00579_ sky130_fd_sc_hd__mux2_1
XANTENNA__10306__S1 net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12081__B1 net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11758_ net195 net2029 net417 vssd1 vssd1 vccd1 vccd1 _00521_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_1486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10709_ net71 net1043 net72 vssd1 vssd1 vccd1 vccd1 _05448_ sky130_fd_sc_hd__or3b_1
XANTENNA__09198__Y _04117_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11689_ net218 net626 vssd1 vssd1 vccd1 vccd1 _06203_ sky130_fd_sc_hd__and2_1
XANTENNA__06615__Y _01566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12793__24 clknet_leaf_31_clk vssd1 vssd1 vccd1 vccd1 net1334 sky130_fd_sc_hd__inv_2
XANTENNA__08035__S net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13428_ clknet_leaf_10_clk _00659_ net1103 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[416\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12384__A1 net197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11187__A2 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13359_ clknet_leaf_41_clk _00590_ net1225 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[347\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_64_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10395__B1 net1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07874__S net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07920_ final_design.cpu.reg_window\[278\] final_design.cpu.reg_window\[310\] net839
+ vssd1 vssd1 vccd1 vccd1 _02871_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_36_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11249__X _05952_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11895__A0 net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07851_ net550 _02799_ vssd1 vssd1 vccd1 vccd1 _02802_ sky130_fd_sc_hd__or2_1
XANTENNA__11409__B net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06802_ final_design.data_from_mem\[22\] net969 _01751_ vssd1 vssd1 vccd1 vccd1 _01753_
+ sky130_fd_sc_hd__o21ai_2
XANTENNA__12917__CLK clknet_leaf_62_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput2 DAT_I[0] vssd1 vssd1 vccd1 vccd1 net2 sky130_fd_sc_hd__dlymetal6s2s_1
X_07782_ net604 _02731_ _02707_ vssd1 vssd1 vccd1 vccd1 _02733_ sky130_fd_sc_hd__o21a_1
XFILLER_0_78_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09521_ _04201_ _04232_ net479 vssd1 vssd1 vccd1 vccd1 _04440_ sky130_fd_sc_hd__mux2_1
X_06733_ _01680_ _01681_ _01682_ _01683_ net775 net793 vssd1 vssd1 vccd1 vccd1 _01684_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_36_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14250__1304 vssd1 vssd1 vccd1 vccd1 _14250__1304/HI net1304 sky130_fd_sc_hd__conb_1
XANTENNA__07315__B2 net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_1829 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09452_ _02768_ net439 _04369_ _02766_ _04370_ vssd1 vssd1 vccd1 vccd1 _04371_ sky130_fd_sc_hd__o221a_1
XFILLER_0_17_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06664_ final_design.cpu.reg_window\[794\] final_design.cpu.reg_window\[826\] net945
+ vssd1 vssd1 vccd1 vccd1 _01615_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_49_1869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08403_ net597 _03352_ _03328_ vssd1 vssd1 vccd1 vccd1 _03354_ sky130_fd_sc_hd__o21ai_1
X_09383_ _01657_ net552 _01717_ net551 net458 net467 vssd1 vssd1 vccd1 vccd1 _04302_
+ sky130_fd_sc_hd__mux4_1
X_06595_ _01542_ _01543_ _01544_ _01545_ net776 net783 vssd1 vssd1 vccd1 vccd1 _01546_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout245_A net247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08334_ _03281_ _03282_ _03283_ _03284_ net674 net691 vssd1 vssd1 vccd1 vccd1 _03285_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__07079__B1 _01821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12072__B1 net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08276__C1 net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08265_ final_design.cpu.reg_window\[906\] final_design.cpu.reg_window\[938\] net817
+ vssd1 vssd1 vccd1 vccd1 _03216_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout412_A net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06525__Y _01476_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1154_A net1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07216_ final_design.cpu.reg_window\[72\] final_design.cpu.reg_window\[104\] net893
+ vssd1 vssd1 vccd1 vccd1 _02167_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08196_ net716 _03146_ vssd1 vssd1 vccd1 vccd1 _03147_ sky130_fd_sc_hd__nor2_1
XFILLER_0_14_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07147_ _02097_ vssd1 vssd1 vccd1 vccd1 _02098_ sky130_fd_sc_hd__inv_2
XANTENNA__08043__A2 _02991_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07078_ final_design.data_from_mem\[13\] net970 _02027_ vssd1 vssd1 vccd1 vccd1 _02029_
+ sky130_fd_sc_hd__o21ai_4
XANTENNA_fanout781_A net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout879_A _01687_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08426__S0 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1008 _05170_ vssd1 vssd1 vccd1 vccd1 net1008 sky130_fd_sc_hd__clkbuf_4
Xfanout1019 _06298_ vssd1 vssd1 vccd1 vccd1 net1019 sky130_fd_sc_hd__buf_2
XANTENNA__07003__B1 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout667_X net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13842__CLK clknet_leaf_44_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08468__X _03419_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07813__A _01660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11638__B1 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09719_ _03070_ _04504_ vssd1 vssd1 vccd1 vccd1 _04638_ sky130_fd_sc_hd__or2_1
X_10991_ _05681_ _05700_ _05716_ vssd1 vssd1 vccd1 vccd1 _05717_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout834_X net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12730_ _06364_ _06370_ final_design.VGA_data_control.v_count\[0\] vssd1 vssd1 vccd1
+ vccd1 _06371_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_2_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12661_ final_design.VGA_data_control.ready_data\[18\] net1020 net975 final_design.data_from_mem\[18\]
+ vssd1 vssd1 vccd1 vccd1 _06318_ sky130_fd_sc_hd__a22o_1
XANTENNA__13992__CLK clknet_leaf_42_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11612_ net427 net564 _06163_ net298 net2303 vssd1 vssd1 vccd1 vccd1 _00438_ sky130_fd_sc_hd__a32o_1
XFILLER_0_13_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12063__B1 net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12592_ net2473 net997 net983 final_design.data_from_mem\[10\] vssd1 vssd1 vccd1
+ vccd1 _01285_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11543_ net430 net569 _06127_ net303 net1653 vssd1 vssd1 vccd1 vccd1 _00405_ sky130_fd_sc_hd__a32o_1
XANTENNA__13222__CLK clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11474_ net204 net2416 net309 vssd1 vssd1 vccd1 vccd1 _00356_ sky130_fd_sc_hd__mux2_1
XANTENNA__09178__C net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12366__A1 net242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_2_Left_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13213_ clknet_leaf_2_clk _00444_ net1064 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[201\]
+ sky130_fd_sc_hd__dfrtp_1
X_10425_ _03096_ _05190_ vssd1 vssd1 vccd1 vccd1 _05196_ sky130_fd_sc_hd__nor2_1
X_14193_ net1310 vssd1 vssd1 vccd1 vccd1 gpio_oeb[5] sky130_fd_sc_hd__buf_2
XANTENNA__10377__B1 net1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13144_ clknet_leaf_65_clk _00375_ net1073 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[132\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13372__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10356_ net29 net1026 _05170_ final_design.data_from_mem\[5\] vssd1 vssd1 vccd1 vccd1
+ _00109_ sky130_fd_sc_hd__a22o_1
XFILLER_0_57_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13075_ clknet_leaf_40_clk _00306_ net1210 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[63\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12105__S net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10287_ net744 net734 _01494_ vssd1 vssd1 vccd1 vccd1 _05143_ sky130_fd_sc_hd__or3_4
X_12026_ _05839_ _06260_ vssd1 vssd1 vccd1 vccd1 _06261_ sky130_fd_sc_hd__nor2_2
XANTENNA__11877__B1 net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11341__A2 net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07723__A _01630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13087__RESET_B net1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09298__A1 _04119_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13977_ clknet_leaf_56_clk _01208_ net1147 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[965\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_17_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12928_ clknet_leaf_47_clk _00166_ net1198 vssd1 vssd1 vccd1 vccd1 net151 sky130_fd_sc_hd__dfrtp_1
XANTENNA__07848__A2 _02797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12859_ clknet_leaf_17_clk _00097_ net1108 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.ready_data\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_44_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1879 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11801__B1 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08050_ final_design.cpu.reg_window\[338\] final_design.cpu.reg_window\[370\] net844
+ vssd1 vssd1 vccd1 vccd1 _03001_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07001_ _01948_ _01949_ _01950_ _01951_ net764 net785 vssd1 vssd1 vccd1 vccd1 _01952_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__13715__CLK clknet_leaf_40_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12357__B2 _06053_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09758__C1 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10368__B1 _05170_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09773__A2 _04406_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12109__A1 net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06587__A2 _01537_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08952_ final_design.CPU_instr_adr\[20\] _03794_ vssd1 vssd1 vccd1 vccd1 _03892_
+ sky130_fd_sc_hd__nor2_1
XANTENNA__13865__CLK clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07903_ final_design.cpu.reg_window\[855\] final_design.cpu.reg_window\[887\] net852
+ vssd1 vssd1 vccd1 vccd1 _02854_ sky130_fd_sc_hd__mux2_1
X_08883_ final_design.CPU_instr_adr\[28\] net1015 _03827_ _03830_ vssd1 vssd1 vccd1
+ vccd1 _00239_ sky130_fd_sc_hd__a22o_1
XANTENNA__11868__B1 net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout195_A _06024_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07834_ net720 _02778_ net723 vssd1 vssd1 vccd1 vccd1 _02785_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_47_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07631__S1 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07765_ final_design.cpu.reg_window\[152\] final_design.cpu.reg_window\[184\] net862
+ vssd1 vssd1 vccd1 vccd1 _02716_ sky130_fd_sc_hd__mux2_1
XANTENNA__09289__A1 _01596_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout362_A net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1773 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09504_ _04195_ _04422_ vssd1 vssd1 vccd1 vccd1 _04423_ sky130_fd_sc_hd__nand2_2
X_06716_ _01663_ _01664_ _01665_ _01666_ net775 net793 vssd1 vssd1 vccd1 vccd1 _01667_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__09384__S1 net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12293__B1 net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07696_ final_design.cpu.reg_window\[411\] final_design.cpu.reg_window\[443\] net868
+ vssd1 vssd1 vccd1 vccd1 _02647_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09435_ _02900_ _04353_ vssd1 vssd1 vccd1 vccd1 _04354_ sky130_fd_sc_hd__xnor2_1
X_06647_ final_design.reqhand.instruction\[27\] final_design.data_from_mem\[27\] net973
+ vssd1 vssd1 vccd1 vccd1 _01598_ sky130_fd_sc_hd__mux2_4
XANTENNA__10843__B2 net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13245__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout248_X net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout627_A _06192_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11442__X _06093_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07779__S net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09366_ _04283_ _04284_ vssd1 vssd1 vccd1 vccd1 _04285_ sky130_fd_sc_hd__or2_1
X_06578_ final_design.cpu.reg_window\[733\] final_design.cpu.reg_window\[765\] net949
+ vssd1 vssd1 vccd1 vccd1 _01529_ sky130_fd_sc_hd__mux2_1
X_08317_ _03264_ _03265_ _03266_ _03267_ net676 net698 vssd1 vssd1 vccd1 vccd1 _03268_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__12596__B2 final_design.data_from_mem\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09297_ net487 net318 _04202_ vssd1 vssd1 vccd1 vccd1 _04216_ sky130_fd_sc_hd__or3_1
XFILLER_0_62_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout415_X net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08248_ _03198_ vssd1 vssd1 vccd1 vccd1 _03199_ sky130_fd_sc_hd__inv_2
XANTENNA__13395__CLK clknet_leaf_40_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout996_A net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08179_ net600 net526 vssd1 vssd1 vccd1 vccd1 _03130_ sky130_fd_sc_hd__nor2_1
XANTENNA__10359__B1 net1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10210_ final_design.uart.BAUD_counter\[3\] _05093_ vssd1 vssd1 vccd1 vccd1 _05095_
+ sky130_fd_sc_hd__or2_1
XANTENNA__11020__A1 _04040_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1777 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11020__B2 _04042_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11190_ net662 _03723_ _04000_ net735 vssd1 vssd1 vccd1 vccd1 _05899_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_54_2040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout784_X net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11571__A2 net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_2051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10141_ _05041_ final_design.h_out vssd1 vssd1 vccd1 vccd1 _05042_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_73_2685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_2062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10072_ net973 _04038_ vssd1 vssd1 vccd1 vccd1 _04990_ sky130_fd_sc_hd__or2_4
XANTENNA_fanout951_X net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11764__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13900_ clknet_leaf_46_clk _01131_ net1216 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[888\]
+ sky130_fd_sc_hd__dfrtp_1
X_13831_ clknet_leaf_59_clk _01062_ net1125 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[819\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14020__CLK clknet_leaf_54_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10886__A1_N net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_67_2478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10974_ _05699_ _05700_ _05679_ _05681_ vssd1 vssd1 vccd1 vccd1 _05701_ sky130_fd_sc_hd__a211oi_1
XANTENNA__11087__B2 net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_2489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12284__B1 net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13762_ clknet_leaf_4_clk _00993_ net1079 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[750\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07386__S0 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12713_ _06352_ _06353_ vssd1 vssd1 vccd1 vccd1 _06354_ sky130_fd_sc_hd__nand2_1
XFILLER_0_6_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13693_ clknet_leaf_2_clk _00924_ net1064 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[681\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_1655 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14170__CLK clknet_leaf_18_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11352__X _06042_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12644_ _06309_ net1447 net978 vssd1 vssd1 vccd1 vccd1 _01324_ sky130_fd_sc_hd__mux2_1
XANTENNA__06593__S net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07138__S0 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12892__Q final_design.data_from_mem\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13738__CLK clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12575_ final_design.uart.working_data\[6\] _06292_ _06286_ vssd1 vssd1 vccd1 vccd1
+ _01272_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11526_ net1758 net194 net522 vssd1 vssd1 vccd1 vccd1 _00393_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14245_ net1299 vssd1 vssd1 vccd1 vccd1 gpio_out[23] sky130_fd_sc_hd__buf_2
X_11457_ net237 net2405 net306 vssd1 vssd1 vccd1 vccd1 _00345_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13888__CLK clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10408_ _03384_ _05181_ vssd1 vssd1 vccd1 vccd1 _05187_ sky130_fd_sc_hd__nor2_1
X_14176_ clknet_leaf_22_clk _01350_ net1164 vssd1 vssd1 vccd1 vccd1 final_design.VGA_adr\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07718__A _01599_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11388_ _04324_ net656 _06073_ vssd1 vssd1 vccd1 vccd1 _06074_ sky130_fd_sc_hd__a21oi_4
XANTENNA__10415__Y _05191_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10339_ net1517 net1010 net987 final_design.data_from_mem\[24\] vssd1 vssd1 vccd1
+ vccd1 _00096_ sky130_fd_sc_hd__a22o_1
X_13127_ clknet_leaf_62_clk _00358_ net1124 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[115\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13118__CLK clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09492__X _04411_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13058_ clknet_leaf_3_clk _00289_ net1066 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[46\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07518__A1 _01686_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11314__A2 _06007_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12009_ _06211_ net285 net402 net2471 vssd1 vssd1 vccd1 vccd1 _00740_ sky130_fd_sc_hd__a22o_1
XANTENNA__10431__X _05199_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_1047 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13268__CLK clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1913 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07550_ net762 _02500_ vssd1 vssd1 vccd1 vccd1 _02501_ sky130_fd_sc_hd__or2_1
XANTENNA__12275__B1 net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06501_ net885 _01445_ _01451_ _01439_ _01436_ vssd1 vssd1 vccd1 vccd1 _01452_ sky130_fd_sc_hd__a32oi_4
XFILLER_0_53_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07481_ _02332_ _02431_ vssd1 vssd1 vccd1 vccd1 _02432_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12290__A3 net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07599__S net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09220_ _03134_ _03164_ _04137_ _04138_ vssd1 vssd1 vccd1 vccd1 _04139_ sky130_fd_sc_hd__a31o_1
X_06432_ net56 vssd1 vssd1 vccd1 vccd1 _01387_ sky130_fd_sc_hd__inv_2
XFILLER_0_53_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_884 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09151_ _03628_ _04053_ vssd1 vssd1 vccd1 vccd1 _04070_ sky130_fd_sc_hd__or2_1
XANTENNA__09099__B net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08102_ net708 _03046_ net722 vssd1 vssd1 vccd1 vccd1 _03053_ sky130_fd_sc_hd__o21a_1
XANTENNA__09667__X _04586_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09082_ net622 _04006_ vssd1 vssd1 vccd1 vccd1 _04007_ sky130_fd_sc_hd__nor2_1
XANTENNA__11250__A1 net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09994__A2 _04411_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08033_ net710 _02983_ vssd1 vssd1 vccd1 vccd1 _02984_ sky130_fd_sc_hd__nor2_1
Xinput60 mem_adr_start[31] vssd1 vssd1 vccd1 vccd1 net60 sky130_fd_sc_hd__clkbuf_1
Xhold800 final_design.cpu.reg_window\[890\] vssd1 vssd1 vccd1 vccd1 net2142 sky130_fd_sc_hd__dlygate4sd3_1
Xinput71 memory_size[12] vssd1 vssd1 vccd1 vccd1 net71 sky130_fd_sc_hd__buf_1
Xhold811 final_design.cpu.reg_window\[765\] vssd1 vssd1 vccd1 vccd1 net2153 sky130_fd_sc_hd__dlygate4sd3_1
Xinput82 memory_size[22] vssd1 vssd1 vccd1 vccd1 net82 sky130_fd_sc_hd__buf_1
XFILLER_0_64_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout208_A _05965_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput93 memory_size[3] vssd1 vssd1 vccd1 vccd1 net93 sky130_fd_sc_hd__clkbuf_2
XANTENNA__11002__A1 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold822 final_design.cpu.reg_window\[740\] vssd1 vssd1 vccd1 vccd1 net2164 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11002__B2 net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09746__A2 _04559_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold833 final_design.cpu.reg_window\[764\] vssd1 vssd1 vccd1 vccd1 net2175 sky130_fd_sc_hd__dlygate4sd3_1
Xhold844 final_design.cpu.reg_window\[784\] vssd1 vssd1 vccd1 vccd1 net2186 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08223__S net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold855 final_design.cpu.reg_window\[853\] vssd1 vssd1 vccd1 vccd1 net2197 sky130_fd_sc_hd__dlygate4sd3_1
Xhold866 final_design.cpu.reg_window\[634\] vssd1 vssd1 vccd1 vccd1 net2208 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08954__B1 net1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11553__A2 net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold877 final_design.cpu.reg_window\[340\] vssd1 vssd1 vccd1 vccd1 net2219 sky130_fd_sc_hd__dlygate4sd3_1
Xhold888 final_design.cpu.reg_window\[157\] vssd1 vssd1 vccd1 vccd1 net2230 sky130_fd_sc_hd__dlygate4sd3_1
Xhold899 final_design.cpu.reg_window\[827\] vssd1 vssd1 vccd1 vccd1 net2241 sky130_fd_sc_hd__dlygate4sd3_1
X_09984_ _04902_ vssd1 vssd1 vccd1 vccd1 _04903_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout1117_A net1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14043__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08935_ final_design.CPU_instr_adr\[21\] _03795_ final_design.CPU_instr_adr\[22\]
+ vssd1 vssd1 vccd1 vccd1 _03877_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_23_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13620__RESET_B net1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11305__A2 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout577_A net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout198_X net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09903__C1 _04120_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08866_ _03776_ _03814_ vssd1 vssd1 vccd1 vccd1 _03815_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_4_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08182__A1 net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07817_ _01657_ _02765_ vssd1 vssd1 vccd1 vccd1 _02768_ sky130_fd_sc_hd__or2_1
X_08797_ _03678_ _03747_ vssd1 vssd1 vccd1 vccd1 _03748_ sky130_fd_sc_hd__nor2_1
XFILLER_0_79_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout365_X net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout744_A _01476_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12266__B1 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07748_ _01630_ net615 vssd1 vssd1 vccd1 vccd1 _02699_ sky130_fd_sc_hd__nor2_1
XANTENNA__11316__C net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_2320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_2954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout911_A net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07679_ final_design.cpu.reg_window\[670\] final_design.cpu.reg_window\[702\] net851
+ vssd1 vssd1 vccd1 vccd1 _02630_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_62_2331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_2965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_2976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1817 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_2987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12018__B1 net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09418_ _01657_ net552 _01717_ net551 net453 net462 vssd1 vssd1 vccd1 vccd1 _04337_
+ sky130_fd_sc_hd__mux4_1
X_10690_ _05425_ _05429_ vssd1 vssd1 vccd1 vccd1 _05430_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_48_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09349_ _04267_ vssd1 vssd1 vccd1 vccd1 _04268_ sky130_fd_sc_hd__inv_2
XFILLER_0_69_1330 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12360_ net2526 net362 net357 _06075_ vssd1 vssd1 vccd1 vccd1 _01072_ sky130_fd_sc_hd__a22o_1
XANTENNA__11241__A1 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11311_ net733 _03893_ vssd1 vssd1 vccd1 vccd1 _06006_ sky130_fd_sc_hd__or2_1
XANTENNA__11759__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_2894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11792__A2 net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12291_ net581 _06221_ net514 net370 net1690 vssd1 vssd1 vccd1 vccd1 _01006_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_56_2113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_2124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_2758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_2135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_2769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14030_ clknet_leaf_43_clk _01261_ net1221 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[1018\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_31_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11242_ net736 _03957_ vssd1 vssd1 vccd1 vccd1 _05945_ sky130_fd_sc_hd__nand2_1
XANTENNA__12741__B2 _05039_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11173_ net2185 net314 net421 _05884_ vssd1 vssd1 vccd1 vccd1 _00278_ sky130_fd_sc_hd__a22o_1
XFILLER_0_38_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input40_A mem_adr_start[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10124_ final_design.VGA_data_control.v_count\[1\] _04998_ _05031_ vssd1 vssd1 vccd1
+ vccd1 _05032_ sky130_fd_sc_hd__and3_1
XANTENNA__11347__X _06038_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10055_ _04701_ _04725_ _04768_ _04884_ vssd1 vssd1 vccd1 vccd1 _04974_ sky130_fd_sc_hd__nand4_1
XANTENNA__13410__CLK clknet_leaf_11_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12887__Q final_design.data_from_mem\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13814_ clknet_leaf_59_clk _01045_ net1138 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[802\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12257__B1 net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07359__S0 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1031 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13560__CLK clknet_leaf_65_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13745_ clknet_leaf_35_clk _00976_ net1240 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[733\]
+ sky130_fd_sc_hd__dfrtp_1
X_10957_ _04040_ _05683_ _05684_ _04042_ vssd1 vssd1 vccd1 vccd1 _05685_ sky130_fd_sc_hd__a22o_1
XANTENNA__08020__S1 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12272__A3 net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12009__B1 net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_851 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13676_ clknet_leaf_45_clk _00907_ net1214 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[664\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10888_ net1055 _05615_ net1000 final_design.CPU_instr_adr\[21\] vssd1 vssd1 vccd1
+ vccd1 _05619_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_6_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07212__S net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06582__S1 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12627_ final_design.VGA_data_control.ready_data\[1\] net1021 net976 final_design.data_from_mem\[1\]
+ vssd1 vssd1 vccd1 vccd1 _06301_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_14_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09487__X _04406_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11232__A1 final_design.data_from_mem\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1051 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12558_ _06221_ net355 net324 net1956 vssd1 vssd1 vccd1 vccd1 _01262_ sky130_fd_sc_hd__a22o_1
XFILLER_0_48_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07531__S0 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11783__A2 net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11509_ net1547 net243 net521 vssd1 vssd1 vccd1 vccd1 _00378_ sky130_fd_sc_hd__mux2_1
Xhold107 net102 vssd1 vssd1 vccd1 vccd1 net1449 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12489_ _06149_ net356 net333 net2140 vssd1 vssd1 vccd1 vccd1 _01195_ sky130_fd_sc_hd__a22o_1
Xhold118 net138 vssd1 vssd1 vccd1 vccd1 net1460 sky130_fd_sc_hd__dlygate4sd3_1
Xhold129 final_design.VGA_data_control.data_to_VGA\[12\] vssd1 vssd1 vccd1 vccd1 net1471
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_65_1761 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14228_ net1282 vssd1 vssd1 vccd1 vccd1 gpio_out[6] sky130_fd_sc_hd__buf_2
XANTENNA__14066__CLK clknet_leaf_15_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14159_ clknet_leaf_14_clk _01333_ net1106 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.data_to_VGA\[18\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout609 net612 vssd1 vssd1 vccd1 vccd1 net609 sky130_fd_sc_hd__buf_2
XFILLER_0_10_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06981_ final_design.cpu.reg_window\[656\] final_design.cpu.reg_window\[688\] net923
+ vssd1 vssd1 vccd1 vccd1 _01932_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11257__X _05959_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13090__CLK clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08720_ final_design.CPU_instr_adr\[19\] _01853_ vssd1 vssd1 vccd1 vccd1 _03671_
+ sky130_fd_sc_hd__or2_1
XANTENNA__06498__S net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12496__B1 net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1180 net1192 vssd1 vssd1 vccd1 vccd1 net1180 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09361__B1 _04279_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1191 net1192 vssd1 vssd1 vccd1 vccd1 net1191 sky130_fd_sc_hd__clkbuf_2
X_08651_ _01627_ _02700_ vssd1 vssd1 vccd1 vccd1 _03602_ sky130_fd_sc_hd__and2_1
XANTENNA__09900__A2 _04087_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08703__A3 _03635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13903__CLK clknet_leaf_42_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07602_ final_design.cpu.reg_window\[29\] final_design.cpu.reg_window\[61\] net871
+ vssd1 vssd1 vccd1 vccd1 _02553_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12248__B1 net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08582_ final_design.cpu.reg_window\[128\] final_design.cpu.reg_window\[160\] net814
+ vssd1 vssd1 vccd1 vccd1 _03533_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_1721 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_38_clk_X clknet_leaf_38_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07533_ final_design.cpu.reg_window\[31\] final_design.cpu.reg_window\[63\] net937
+ vssd1 vssd1 vccd1 vccd1 _02484_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_1765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08467__A2 _03415_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07464_ final_design.cpu.reg_window\[576\] final_design.cpu.reg_window\[608\] net909
+ vssd1 vssd1 vccd1 vccd1 _02415_ sky130_fd_sc_hd__mux2_1
XANTENNA__08218__S net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06415_ final_design.VGA_data_control.v_count\[6\] vssd1 vssd1 vccd1 vccd1 _01370_
+ sky130_fd_sc_hd__inv_2
X_09203_ _04106_ _04110_ _04119_ _04121_ _04115_ vssd1 vssd1 vccd1 vccd1 _04122_ sky130_fd_sc_hd__o311a_1
X_07395_ final_design.cpu.reg_window\[898\] final_design.cpu.reg_window\[930\] net913
+ vssd1 vssd1 vccd1 vccd1 _02346_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout325_A _06285_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09416__B2 _04073_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1067_A net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09134_ _03647_ net659 vssd1 vssd1 vccd1 vccd1 _04053_ sky130_fd_sc_hd__nand2b_4
XANTENNA__12420__B1 net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09065_ _03699_ _03724_ vssd1 vssd1 vccd1 vccd1 _03992_ sky130_fd_sc_hd__xor2_1
XFILLER_0_60_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1234_A net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08016_ final_design.cpu.reg_window\[339\] final_design.cpu.reg_window\[371\] net830
+ vssd1 vssd1 vccd1 vccd1 _02967_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold630 final_design.cpu.reg_window\[75\] vssd1 vssd1 vccd1 vccd1 net1972 sky130_fd_sc_hd__dlygate4sd3_1
Xhold641 final_design.cpu.reg_window\[38\] vssd1 vssd1 vccd1 vccd1 net1983 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout694_A net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_2600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold652 final_design.cpu.reg_window\[350\] vssd1 vssd1 vccd1 vccd1 net1994 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_70_2611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold663 final_design.cpu.reg_window\[130\] vssd1 vssd1 vccd1 vccd1 net2005 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13119__RESET_B net1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13433__CLK clknet_leaf_56_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold674 final_design.cpu.reg_window\[227\] vssd1 vssd1 vccd1 vccd1 net2016 sky130_fd_sc_hd__dlygate4sd3_1
Xhold685 final_design.cpu.reg_window\[181\] vssd1 vssd1 vccd1 vccd1 net2027 sky130_fd_sc_hd__dlygate4sd3_1
X_14189__1248 vssd1 vssd1 vccd1 vccd1 _14189__1248/HI net1248 sky130_fd_sc_hd__conb_1
XFILLER_0_44_1889 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07792__S net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold696 final_design.cpu.reg_window\[41\] vssd1 vssd1 vccd1 vccd1 net2038 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09967_ net96 _04179_ net97 vssd1 vssd1 vccd1 vccd1 _04886_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout861_A net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout482_X net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout959_A _04041_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08918_ _03753_ _03765_ _03761_ vssd1 vssd1 vccd1 vccd1 _03861_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_77_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12487__B1 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09898_ net475 _04814_ _04816_ vssd1 vssd1 vccd1 vccd1 _04817_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_58_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09352__B1 net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07093__A net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13583__CLK clknet_leaf_42_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08849_ final_design.CPU_instr_adr\[28\] final_design.CPU_instr_adr\[27\] _03799_
+ vssd1 vssd1 vccd1 vccd1 _03800_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_68_2540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout747_X net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10501__A3 net250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_2404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12239__B1 net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11860_ _06106_ net290 net520 net2552 vssd1 vssd1 vccd1 vccd1 _00608_ sky130_fd_sc_hd__a22o_1
XFILLER_0_79_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10811_ _05541_ _05543_ _05545_ net1032 net1357 vssd1 vssd1 vccd1 vccd1 _00190_ sky130_fd_sc_hd__a32o_1
XFILLER_0_16_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11791_ net2401 net414 net287 _05981_ vssd1 vssd1 vccd1 vccd1 _00547_ sky130_fd_sc_hd__a22o_1
XFILLER_0_39_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06469__A1 final_design.data_from_mem\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13530_ clknet_leaf_64_clk _00761_ net1075 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[518\]
+ sky130_fd_sc_hd__dfrtp_1
X_10742_ _05458_ _05479_ vssd1 vssd1 vccd1 vccd1 _05480_ sky130_fd_sc_hd__nand2_1
XANTENNA__06437__A net35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07032__S net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07761__S0 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06564__S1 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10673_ net1054 _05412_ _05413_ vssd1 vssd1 vccd1 vccd1 _05414_ sky130_fd_sc_hd__a21o_1
X_13461_ clknet_leaf_57_clk _00692_ net1144 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[449\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_11_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12412_ _06107_ net343 net338 net1735 vssd1 vssd1 vccd1 vccd1 _01122_ sky130_fd_sc_hd__a22o_1
XANTENNA__12411__B1 net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input88_A memory_size[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13392_ clknet_leaf_34_clk _00623_ net1238 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[380\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14089__CLK clknet_leaf_25_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11489__S net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12343_ net2418 net360 net344 _05952_ vssd1 vssd1 vccd1 vccd1 _01055_ sky130_fd_sc_hd__a22o_1
XANTENNA__08371__B _03321_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_1901 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12274_ net561 _06204_ net503 net368 net1831 vssd1 vssd1 vccd1 vccd1 _00989_ sky130_fd_sc_hd__a32o_1
XANTENNA__09186__C net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08069__S1 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10406__B _05181_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11225_ final_design.data_from_mem\[10\] _05914_ _05917_ vssd1 vssd1 vccd1 vccd1
+ _05930_ sky130_fd_sc_hd__a21o_1
X_14013_ clknet_leaf_1_clk _01244_ net1077 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[1001\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07555__X _02506_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11156_ net429 _05865_ net567 net315 net2096 vssd1 vssd1 vccd1 vccd1 _00276_ sky130_fd_sc_hd__a32o_1
XANTENNA__13926__CLK clknet_leaf_51_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10107_ _05007_ _05020_ _05021_ vssd1 vssd1 vccd1 vccd1 final_design.vga.v_next_count\[1\]
+ sky130_fd_sc_hd__and3_1
XFILLER_0_65_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_8_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11518__A net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11087_ net956 _05808_ _05807_ net960 vssd1 vssd1 vccd1 vccd1 _05809_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__12478__B1 net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12113__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10038_ _04954_ _04955_ vssd1 vssd1 vccd1 vccd1 _04957_ sky130_fd_sc_hd__xnor2_1
XANTENNA__11150__B1 _05843_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12950__CLK clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12245__A3 net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11989_ _06191_ net288 net407 net1749 vssd1 vssd1 vccd1 vccd1 _00722_ sky130_fd_sc_hd__a22o_1
XANTENNA__11253__A net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13728_ clknet_leaf_11_clk _00959_ net1087 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[716\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_50_clk_A clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13306__CLK clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1135 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13659_ clknet_leaf_66_clk _00890_ net1063 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[647\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10008__A2 _04045_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07180_ final_design.cpu.reg_window\[329\] final_design.cpu.reg_window\[361\] net901
+ vssd1 vssd1 vccd1 vccd1 _02131_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_26_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12402__B1 net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_65_clk_A clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13456__CLK clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08281__B net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06632__A1 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07178__A _02127_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1119 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_6_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout406 _06255_ vssd1 vssd1 vccd1 vccd1 net406 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_26_1586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout417 net419 vssd1 vssd1 vccd1 vccd1 net417 sky130_fd_sc_hd__buf_4
X_09821_ _03262_ _03574_ _04738_ _04739_ vssd1 vssd1 vccd1 vccd1 _04740_ sky130_fd_sc_hd__a31o_1
Xfanout428 net429 vssd1 vssd1 vccd1 vccd1 net428 sky130_fd_sc_hd__clkbuf_4
XANTENNA_clkload12_A clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout439 _04095_ vssd1 vssd1 vccd1 vccd1 net439 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08480__S1 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07593__C1 net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12469__B1 net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09752_ _04072_ _04662_ _04666_ _04670_ vssd1 vssd1 vccd1 vccd1 _04671_ sky130_fd_sc_hd__or4b_1
X_06964_ final_design.cpu.reg_window\[464\] final_design.cpu.reg_window\[496\] net926
+ vssd1 vssd1 vccd1 vccd1 _01915_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08703_ _02510_ _03611_ _03635_ _03653_ _03634_ vssd1 vssd1 vccd1 vccd1 _03654_ sky130_fd_sc_hd__o311a_1
X_06895_ final_design.cpu.reg_window\[595\] final_design.cpu.reg_window\[627\] net903
+ vssd1 vssd1 vccd1 vccd1 _01846_ sky130_fd_sc_hd__mux2_1
X_09683_ _03164_ _04087_ net440 _03162_ _04601_ vssd1 vssd1 vccd1 vccd1 _04602_ sky130_fd_sc_hd__a221o_1
XANTENNA__08688__A2 _03550_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07912__Y _02863_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08634_ _03296_ _03569_ _03578_ _03584_ vssd1 vssd1 vccd1 vccd1 _03585_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_55_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11692__A1 net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06956__S net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07991__S0 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09637__A1 net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08565_ _02394_ net608 vssd1 vssd1 vccd1 vccd1 _03516_ sky130_fd_sc_hd__or2_1
XANTENNA__12236__A3 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09637__B2 net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout442_A net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1901 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11163__A net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07516_ _01725_ _02465_ _01724_ vssd1 vssd1 vccd1 vccd1 _02467_ sky130_fd_sc_hd__a21o_1
XANTENNA_clkbuf_leaf_18_clk_A clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08496_ final_design.cpu.reg_window\[515\] final_design.cpu.reg_window\[547\] net825
+ vssd1 vssd1 vccd1 vccd1 _03447_ sky130_fd_sc_hd__mux2_1
X_12799__30 clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 net1340 sky130_fd_sc_hd__inv_2
XANTENNA__07112__A2 _01498_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11995__A2 net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07447_ final_design.cpu.reg_window\[448\] final_design.cpu.reg_window\[480\] net907
+ vssd1 vssd1 vccd1 vccd1 _02398_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout707_A net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout328_X net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_21_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07378_ final_design.reqhand.instruction\[10\] net972 _02327_ vssd1 vssd1 vccd1 vccd1
+ _02329_ sky130_fd_sc_hd__o21a_1
XANTENNA_clkbuf_3_5_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09117_ net995 net992 net1040 vssd1 vssd1 vccd1 vccd1 _04036_ sky130_fd_sc_hd__a21o_2
XANTENNA__09287__B _04097_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11102__S net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09048_ net622 _03976_ vssd1 vssd1 vccd1 vccd1 _03977_ sky130_fd_sc_hd__nor2_1
XANTENNA__13949__CLK clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout697_X net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold460 final_design.cpu.reg_window\[775\] vssd1 vssd1 vccd1 vccd1 net1802 sky130_fd_sc_hd__dlygate4sd3_1
Xhold471 final_design.reqhand.instruction\[3\] vssd1 vssd1 vccd1 vccd1 net1813 sky130_fd_sc_hd__dlygate4sd3_1
X_11010_ _04286_ net252 _04990_ vssd1 vssd1 vccd1 vccd1 _05735_ sky130_fd_sc_hd__o21a_1
Xhold482 final_design.cpu.reg_window\[791\] vssd1 vssd1 vccd1 vccd1 net1824 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07375__X _02326_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold493 final_design.cpu.reg_window\[862\] vssd1 vssd1 vccd1 vccd1 net1835 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_1705 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout864_X net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout940 net952 vssd1 vssd1 vccd1 vccd1 net940 sky130_fd_sc_hd__buf_2
XFILLER_0_79_1749 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout951 net952 vssd1 vssd1 vccd1 vccd1 net951 sky130_fd_sc_hd__clkbuf_2
Xfanout962 _04036_ vssd1 vssd1 vccd1 vccd1 net962 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12935__RESET_B net1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout973 _01415_ vssd1 vssd1 vccd1 vccd1 net973 sky130_fd_sc_hd__buf_4
Xfanout984 net985 vssd1 vssd1 vccd1 vccd1 net984 sky130_fd_sc_hd__clkbuf_4
Xfanout995 _01408_ vssd1 vssd1 vccd1 vccd1 net995 sky130_fd_sc_hd__buf_2
X_12961_ clknet_leaf_32_clk _00199_ net1233 vssd1 vssd1 vccd1 vccd1 net119 sky130_fd_sc_hd__dfrtp_1
Xhold1160 final_design.cpu.reg_window\[821\] vssd1 vssd1 vccd1 vccd1 net2502 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_73_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1171 final_design.CPU_instr_adr\[19\] vssd1 vssd1 vccd1 vccd1 net2513 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1182 final_design.CPU_instr_adr\[13\] vssd1 vssd1 vccd1 vccd1 net2524 sky130_fd_sc_hd__dlygate4sd3_1
X_11912_ net189 net2077 net275 vssd1 vssd1 vccd1 vccd1 _00652_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12892_ clknet_leaf_15_clk _00130_ net1107 vssd1 vssd1 vccd1 vccd1 final_design.data_from_mem\[26\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__08647__A _01658_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1193 final_design.cpu.reg_window\[828\] vssd1 vssd1 vccd1 vccd1 net2535 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_9_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13329__CLK clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06785__S1 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11843_ net672 net638 vssd1 vssd1 vccd1 vccd1 _06238_ sky130_fd_sc_hd__and2_2
XFILLER_0_5_1709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12227__A3 net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11073__A _05172_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11774_ net648 net555 net227 vssd1 vssd1 vccd1 vccd1 _06230_ sky130_fd_sc_hd__and3_1
XANTENNA__09723__S1 net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13513_ clknet_leaf_36_clk _00744_ net1230 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[501\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11986__A2 net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10725_ _05425_ _05429_ _05448_ vssd1 vssd1 vccd1 vccd1 _05463_ sky130_fd_sc_hd__or3b_1
XFILLER_0_82_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13479__CLK clknet_leaf_63_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11360__X _06049_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13444_ clknet_leaf_54_clk _00675_ net1180 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[432\]
+ sky130_fd_sc_hd__dfrtp_1
X_10656_ net1054 _05394_ net1001 final_design.CPU_instr_adr\[10\] vssd1 vssd1 vccd1
+ vccd1 _05398_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_42_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkload16 clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 clkload16/X sky130_fd_sc_hd__clkbuf_8
X_10587_ net97 final_design.VGA_adr\[5\] vssd1 vssd1 vccd1 vccd1 _05332_ sky130_fd_sc_hd__or2_1
XANTENNA__12108__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload27 clknet_leaf_38_clk vssd1 vssd1 vccd1 vccd1 clkload27/X sky130_fd_sc_hd__clkbuf_8
X_13375_ clknet_leaf_7_clk _00606_ net1134 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[363\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08603__A2 _03550_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload38 clknet_leaf_28_clk vssd1 vssd1 vccd1 vccd1 clkload38/X sky130_fd_sc_hd__clkbuf_8
XANTENNA__10417__A _03257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06929__A1_N net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12326_ net2247 net181 net366 vssd1 vssd1 vccd1 vccd1 _01040_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_1742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12257_ net581 _06186_ net514 net374 net1921 vssd1 vssd1 vccd1 vccd1 _00973_ sky130_fd_sc_hd__a32o_1
XANTENNA__09564__B1 net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11208_ net660 _03983_ net732 vssd1 vssd1 vccd1 vccd1 _05915_ sky130_fd_sc_hd__o21a_1
X_12188_ net1752 net191 net383 vssd1 vssd1 vccd1 vccd1 _00907_ sky130_fd_sc_hd__mux2_1
XANTENNA__10423__Y _05195_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08462__S1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11371__B1 _05143_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11910__A2 _06248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11248__A net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11139_ _01395_ _04037_ vssd1 vssd1 vccd1 vccd1 _05854_ sky130_fd_sc_hd__nor2_1
XANTENNA__14104__CLK clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_3002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09867__A1 _04125_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_3013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_3024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_3035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11674__A1 net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07878__B1 net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06680_ _01627_ _01630_ vssd1 vssd1 vccd1 vccd1 _01631_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_82_3046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12218__A3 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08350_ final_design.cpu.reg_window\[391\] final_design.cpu.reg_window\[423\] net811
+ vssd1 vssd1 vccd1 vccd1 _03301_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11426__A1 net223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12791__22_A clknet_leaf_30_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09095__A2 net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07301_ final_design.cpu.reg_window\[389\] final_design.cpu.reg_window\[421\] net919
+ vssd1 vssd1 vccd1 vccd1 _02252_ sky130_fd_sc_hd__mux2_1
X_14188__1247 vssd1 vssd1 vccd1 vccd1 _14188__1247/HI net1247 sky130_fd_sc_hd__conb_1
XANTENNA__11977__A2 net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08281_ _02157_ net612 vssd1 vssd1 vccd1 vccd1 _03232_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_24_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11270__X _05970_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_24_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11711__A net197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07232_ net749 _02182_ vssd1 vssd1 vccd1 vccd1 _02183_ sky130_fd_sc_hd__or2_1
XFILLER_0_15_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12846__CLK clknet_leaf_17_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07400__S net913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07163_ final_design.cpu.reg_window\[842\] final_design.cpu.reg_window\[874\] net907
+ vssd1 vssd1 vccd1 vccd1 _02114_ sky130_fd_sc_hd__mux2_1
X_07094_ net750 _02038_ net745 vssd1 vssd1 vccd1 vccd1 _02045_ sky130_fd_sc_hd__o21a_1
XFILLER_0_67_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08358__A1 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout203 _05989_ vssd1 vssd1 vccd1 vccd1 net203 sky130_fd_sc_hd__buf_2
Xfanout214 net215 vssd1 vssd1 vccd1 vccd1 net214 sky130_fd_sc_hd__buf_2
XFILLER_0_5_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout225 _05897_ vssd1 vssd1 vccd1 vccd1 net225 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout392_A net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout236 _05982_ vssd1 vssd1 vccd1 vccd1 net236 sky130_fd_sc_hd__buf_1
Xfanout247 _04986_ vssd1 vssd1 vccd1 vccd1 net247 sky130_fd_sc_hd__clkbuf_4
X_09804_ net447 _04707_ _04717_ _04722_ vssd1 vssd1 vccd1 vccd1 _04723_ sky130_fd_sc_hd__o22a_2
Xfanout258 net259 vssd1 vssd1 vccd1 vccd1 net258 sky130_fd_sc_hd__clkbuf_4
Xfanout269 net271 vssd1 vssd1 vccd1 vccd1 net269 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_66_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07996_ _02943_ _02944_ _02945_ _02946_ net682 net702 vssd1 vssd1 vccd1 vccd1 _02947_
+ sky130_fd_sc_hd__mux4_1
X_09735_ net728 _04639_ _04653_ vssd1 vssd1 vccd1 vccd1 _04654_ sky130_fd_sc_hd__and3_1
XANTENNA__12688__S net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06947_ final_design.cpu.reg_window\[785\] final_design.cpu.reg_window\[817\] net926
+ vssd1 vssd1 vccd1 vccd1 _01898_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout657_A net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09666_ net472 _04297_ net486 vssd1 vssd1 vccd1 vccd1 _04585_ sky130_fd_sc_hd__a21oi_1
X_06878_ final_design.cpu.reg_window\[403\] final_design.cpu.reg_window\[435\] net902
+ vssd1 vssd1 vccd1 vccd1 _01829_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08530__B2 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08617_ _03426_ _03561_ _03567_ vssd1 vssd1 vccd1 vccd1 _03568_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_55_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout824_A net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09597_ net484 _04442_ _04515_ _04056_ vssd1 vssd1 vccd1 vccd1 _04516_ sky130_fd_sc_hd__a211o_1
XANTENNA__12209__A3 net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout445_X net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13621__CLK clknet_leaf_58_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08548_ net718 _03498_ vssd1 vssd1 vccd1 vccd1 _03499_ sky130_fd_sc_hd__or2_1
XANTENNA__11324__C _06016_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1917 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12090__A1 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout612_X net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08479_ final_design.cpu.reg_window\[387\] final_design.cpu.reg_window\[419\] net835
+ vssd1 vssd1 vccd1 vccd1 _03430_ sky130_fd_sc_hd__mux2_1
XANTENNA__11621__A net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10510_ net958 _05255_ _05258_ net955 vssd1 vssd1 vccd1 vccd1 _05259_ sky130_fd_sc_hd__o22a_1
XFILLER_0_11_1641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11490_ net183 net640 vssd1 vssd1 vccd1 vccd1 _06113_ sky130_fd_sc_hd__and2_1
XFILLER_0_52_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13771__CLK clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10441_ net1393 net1033 _05204_ net248 vssd1 vssd1 vccd1 vccd1 _00161_ sky130_fd_sc_hd__a22o_1
XANTENNA__10928__B1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10372_ net15 net1025 net1008 final_design.data_from_mem\[21\] vssd1 vssd1 vccd1
+ vccd1 _00125_ sky130_fd_sc_hd__a22o_1
X_13160_ clknet_leaf_35_clk _00391_ net1237 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[148\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout981_X net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12111_ net2059 net222 net391 vssd1 vssd1 vccd1 vccd1 _00835_ sky130_fd_sc_hd__mux2_1
XANTENNA__11767__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13091_ clknet_leaf_0_clk _00322_ net1069 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[79\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14127__CLK clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12042_ net1679 net205 net396 vssd1 vssd1 vccd1 vccd1 _00770_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold290 final_design.cpu.reg_window\[914\] vssd1 vssd1 vccd1 vccd1 net1632 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08141__S net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09010__A2 net1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11353__B1 _06042_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout770 net771 vssd1 vssd1 vccd1 vccd1 net770 sky130_fd_sc_hd__buf_4
XANTENNA__13151__CLK clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout781 net782 vssd1 vssd1 vccd1 vccd1 net781 sky130_fd_sc_hd__buf_2
Xfanout792 net795 vssd1 vssd1 vccd1 vccd1 net792 sky130_fd_sc_hd__clkbuf_4
X_13993_ clknet_leaf_37_clk _01224_ net1231 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[981\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11355__X _06045_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12944_ clknet_leaf_29_clk _00182_ net1193 vssd1 vssd1 vccd1 vccd1 net132 sky130_fd_sc_hd__dfrtp_1
XANTENNA__10459__A2 net1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11656__A1 net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09313__A3 _02091_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12895__Q final_design.data_from_mem\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06758__S1 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12875_ clknet_leaf_17_clk _00113_ net1108 vssd1 vssd1 vccd1 vccd1 final_design.data_from_mem\[9\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__12787__18_A clknet_leaf_27_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11826_ net206 net1989 net264 vssd1 vssd1 vccd1 vccd1 _00578_ sky130_fd_sc_hd__mux2_1
XANTENNA__12869__CLK clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09700__S net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11959__A2 net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11757_ net196 net2105 net418 vssd1 vssd1 vccd1 vccd1 _00520_ sky130_fd_sc_hd__mux2_1
X_10708_ net71 net1043 _05445_ _05446_ vssd1 vssd1 vccd1 vccd1 _05447_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__08316__S net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11688_ net425 net559 _06202_ net294 net2228 vssd1 vssd1 vccd1 vccd1 _00475_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_42_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13427_ clknet_leaf_39_clk _00658_ net1211 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[415\]
+ sky130_fd_sc_hd__dfrtp_1
X_10639_ net801 _05378_ _05381_ _05367_ vssd1 vssd1 vccd1 vccd1 _05382_ sky130_fd_sc_hd__o211a_1
XFILLER_0_24_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13358_ clknet_leaf_42_clk _00589_ net1223 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[346\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10395__A1 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10395__B2 net169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12309_ net1729 net213 net364 vssd1 vssd1 vccd1 vccd1 _01023_ sky130_fd_sc_hd__mux2_1
XANTENNA__07260__B2 net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13289_ clknet_leaf_37_clk _00520_ net1229 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[277\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09147__S _03484_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_18_Right_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_36_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11344__B1 net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07850_ net616 _02797_ _02798_ net550 vssd1 vssd1 vccd1 vccd1 _02801_ sky130_fd_sc_hd__a211oi_2
XANTENNA__09552__A3 _04157_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07890__S net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09671__A net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06801_ final_design.data_from_mem\[22\] net969 _01751_ vssd1 vssd1 vccd1 vccd1 _01752_
+ sky130_fd_sc_hd__o21a_4
X_07781_ _01690_ net604 vssd1 vssd1 vccd1 vccd1 _02732_ sky130_fd_sc_hd__and2_1
Xinput3 DAT_I[10] vssd1 vssd1 vccd1 vccd1 net3 sky130_fd_sc_hd__clkbuf_1
XANTENNA__06771__B1 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09520_ net486 _04435_ _04438_ vssd1 vssd1 vccd1 vccd1 _04439_ sky130_fd_sc_hd__a21o_1
XANTENNA__13644__CLK clknet_leaf_45_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06732_ final_design.cpu.reg_window\[664\] final_design.cpu.reg_window\[696\] net942
+ vssd1 vssd1 vccd1 vccd1 _01683_ sky130_fd_sc_hd__mux2_1
XANTENNA__12301__S net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08287__A net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06663_ final_design.cpu.reg_window\[858\] final_design.cpu.reg_window\[890\] net945
+ vssd1 vssd1 vccd1 vccd1 _01614_ sky130_fd_sc_hd__mux2_1
X_09451_ _04085_ _04093_ vssd1 vssd1 vccd1 vccd1 _04370_ sky130_fd_sc_hd__nand2_1
XFILLER_0_56_1376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07720__C1 _01596_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11537__C_N net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08402_ _02240_ net610 vssd1 vssd1 vccd1 vccd1 _03353_ sky130_fd_sc_hd__nor2_1
X_09382_ _04299_ _04300_ net479 vssd1 vssd1 vccd1 vccd1 _04301_ sky130_fd_sc_hd__mux2_1
X_06594_ final_design.cpu.reg_window\[28\] final_design.cpu.reg_window\[60\] net946
+ vssd1 vssd1 vccd1 vccd1 _01545_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_27_Right_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09699__S0 net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13794__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08333_ final_design.cpu.reg_window\[520\] final_design.cpu.reg_window\[552\] net812
+ vssd1 vssd1 vccd1 vccd1 _03284_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08264_ final_design.cpu.reg_window\[970\] final_design.cpu.reg_window\[1002\] net817
+ vssd1 vssd1 vccd1 vccd1 _03215_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_1737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08226__S net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07215_ final_design.cpu.reg_window\[136\] final_design.cpu.reg_window\[168\] net893
+ vssd1 vssd1 vccd1 vccd1 _02166_ sky130_fd_sc_hd__mux2_1
X_08195_ _03142_ _03143_ _03144_ _03145_ net675 net697 vssd1 vssd1 vccd1 vccd1 _03146_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout405_A _06255_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07146_ net665 _02092_ _02093_ _02096_ vssd1 vssd1 vccd1 vccd1 _02097_ sky130_fd_sc_hd__a211o_2
XFILLER_0_42_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11583__B1 net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07077_ final_design.data_from_mem\[13\] net970 _02027_ vssd1 vssd1 vccd1 vccd1 _02028_
+ sky130_fd_sc_hd__o21a_2
XPHY_EDGE_ROW_36_Right_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13174__CLK clknet_leaf_60_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1009 _05166_ vssd1 vssd1 vccd1 vccd1 net1009 sky130_fd_sc_hd__buf_2
XANTENNA__08426__S1 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout774_A net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout395_X net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07003__A1 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout941_A net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout562_X net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07979_ net603 _02929_ vssd1 vssd1 vccd1 vccd1 _02930_ sky130_fd_sc_hd__nor2_1
X_09718_ _04635_ _04636_ _04599_ _04616_ vssd1 vssd1 vccd1 vccd1 _04637_ sky130_fd_sc_hd__a211o_1
XANTENNA__11638__A1 net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10990_ _05679_ _05700_ _05699_ vssd1 vssd1 vccd1 vccd1 _05716_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_2_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09649_ _03026_ _04427_ _02996_ vssd1 vssd1 vccd1 vccd1 _04568_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_6_1804 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_45_Right_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12660_ _06317_ net1455 net979 vssd1 vssd1 vccd1 vccd1 _01332_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11611_ net226 net630 vssd1 vssd1 vccd1 vccd1 _06163_ sky130_fd_sc_hd__and2_1
XFILLER_0_26_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12591_ net1387 net997 net983 final_design.data_from_mem\[9\] vssd1 vssd1 vccd1 vccd1
+ _01284_ sky130_fd_sc_hd__a22o_1
XANTENNA__08644__B _02772_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11542_ net241 net635 vssd1 vssd1 vccd1 vccd1 _06127_ sky130_fd_sc_hd__and2_1
XANTENNA__08136__S net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11473_ net223 net2344 net309 vssd1 vssd1 vccd1 vccd1 _00355_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input70_A memory_size[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13212_ clknet_leaf_3_clk _00443_ net1066 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[200\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09767__B1 net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10424_ net1584 net1027 _05195_ net245 vssd1 vssd1 vccd1 vccd1 _00153_ sky130_fd_sc_hd__a22o_1
X_14192_ net1251 vssd1 vssd1 vccd1 vccd1 gpio_oeb[4] sky130_fd_sc_hd__buf_2
XANTENNA__13517__CLK clknet_leaf_44_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10377__B2 final_design.data_from_mem\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_54_Right_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13143_ clknet_leaf_5_clk _00374_ net1081 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[131\]
+ sky130_fd_sc_hd__dfrtp_1
X_10355_ net28 net1023 net1006 final_design.data_from_mem\[4\] vssd1 vssd1 vccd1 vccd1
+ _00108_ sky130_fd_sc_hd__o22a_1
X_13074_ clknet_leaf_39_clk _00305_ net1209 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[62\]
+ sky130_fd_sc_hd__dfrtp_1
X_10286_ net741 net731 _01495_ vssd1 vssd1 vccd1 vccd1 _05142_ sky130_fd_sc_hd__and3_2
XFILLER_0_44_1280 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11326__B1 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output157_A net157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12025_ net804 _05841_ vssd1 vssd1 vccd1 vccd1 _06260_ sky130_fd_sc_hd__nand2_4
XANTENNA__13667__CLK clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08659__X _03610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1917 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08742__A1 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07563__X _02514_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06753__B1 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12121__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13976_ clknet_leaf_65_clk _01207_ net1076 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[964\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_63_Right_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_17_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12927_ clknet_leaf_47_clk _00165_ net1198 vssd1 vssd1 vccd1 vccd1 net150 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_17_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12858_ clknet_leaf_18_clk _00096_ net1106 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.ready_data\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_44_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11809_ net2462 net414 net288 _06090_ vssd1 vssd1 vccd1 vccd1 _00562_ sky130_fd_sc_hd__a22o_1
XANTENNA__13047__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11262__C1 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09207__C1 _03610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_72_Right_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07000_ final_design.cpu.reg_window\[143\] final_design.cpu.reg_window\[175\] net888
+ vssd1 vssd1 vccd1 vccd1 _01951_ sky130_fd_sc_hd__mux2_1
XANTENNA__12357__A2 net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13197__CLK clknet_leaf_48_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10368__B2 final_design.data_from_mem\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11565__B1 net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07233__A1 net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10164__X _05058_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06667__S0 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11200__S net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08951_ _02461_ _03889_ _03890_ net621 net258 vssd1 vssd1 vccd1 vccd1 _03891_ sky130_fd_sc_hd__a221o_1
X_07902_ final_design.cpu.reg_window\[919\] final_design.cpu.reg_window\[951\] net852
+ vssd1 vssd1 vccd1 vccd1 _02853_ sky130_fd_sc_hd__mux2_1
XANTENNA__11868__A1 net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08882_ _03655_ _03829_ net1038 vssd1 vssd1 vccd1 vccd1 _03830_ sky130_fd_sc_hd__o21a_1
XANTENNA__07914__A _01722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07092__S0 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07833_ net712 _02783_ vssd1 vssd1 vccd1 vccd1 _02784_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_81_Right_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout188_A _06045_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12031__S net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07764_ final_design.cpu.reg_window\[216\] final_design.cpu.reg_window\[248\] net862
+ vssd1 vssd1 vccd1 vccd1 _02715_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07125__S net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09503_ net88 _04194_ vssd1 vssd1 vccd1 vccd1 _04422_ sky130_fd_sc_hd__nand2_1
XFILLER_0_71_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06715_ final_design.cpu.reg_window\[152\] final_design.cpu.reg_window\[184\] net942
+ vssd1 vssd1 vccd1 vccd1 _01666_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07695_ final_design.cpu.reg_window\[475\] final_design.cpu.reg_window\[507\] net863
+ vssd1 vssd1 vccd1 vccd1 _02646_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout355_A net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09434_ _02838_ _04352_ _03036_ _03035_ vssd1 vssd1 vccd1 vccd1 _04353_ sky130_fd_sc_hd__a211o_1
X_06646_ net884 _01589_ _01595_ _01582_ _01583_ vssd1 vssd1 vccd1 vccd1 _01597_ sky130_fd_sc_hd__a32o_2
XFILLER_0_52_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_1059 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09365_ _02672_ _02702_ _04282_ net448 vssd1 vssd1 vccd1 vccd1 _04284_ sky130_fd_sc_hd__a31o_1
XFILLER_0_47_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout522_A net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06577_ net753 _01527_ vssd1 vssd1 vccd1 vccd1 _01528_ sky130_fd_sc_hd__or2_1
XFILLER_0_75_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12596__A2 net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08316_ final_design.cpu.reg_window\[392\] final_design.cpu.reg_window\[424\] net829
+ vssd1 vssd1 vccd1 vccd1 _03267_ sky130_fd_sc_hd__mux2_1
XANTENNA__09997__B1 _04914_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_2270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09296_ _04211_ _04214_ net473 vssd1 vssd1 vccd1 vccd1 _04215_ sky130_fd_sc_hd__mux2_1
XANTENNA_30 _06257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_1780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout310_X net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08247_ _03195_ _03196_ vssd1 vssd1 vccd1 vccd1 _03198_ sky130_fd_sc_hd__or2_2
XFILLER_0_65_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout408_X net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1052_X net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12348__A2 net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09749__B1 net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10359__A1 net32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08178_ _03116_ _03117_ _03128_ net874 vssd1 vssd1 vccd1 vccd1 _03129_ sky130_fd_sc_hd__a22oi_2
XANTENNA__06552__X _01503_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10359__B2 final_design.data_from_mem\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout891_A net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout989_A _05167_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08421__B1 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07129_ final_design.cpu.reg_window\[843\] final_design.cpu.reg_window\[875\] net909
+ vssd1 vssd1 vccd1 vccd1 _02080_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_1789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_54_2041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10140_ final_design.VGA_data_control.h_count\[5\] _05014_ _05010_ final_design.vga.h_current_state\[1\]
+ final_design.vga.h_current_state\[0\] vssd1 vssd1 vccd1 vccd1 final_design.h_out
+ sky130_fd_sc_hd__a2111o_1
XANTENNA__08972__A1 net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_2052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_2063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput170 net170 vssd1 vssd1 vccd1 vccd1 STB_O sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_73_2697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout777_X net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10071_ net973 _04038_ vssd1 vssd1 vccd1 vccd1 _04989_ sky130_fd_sc_hd__nor2_1
XANTENNA__11859__B2 net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12520__A2 net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout944_X net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13830_ clknet_leaf_51_clk _01061_ net1171 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[818\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13567__RESET_B net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07035__S net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_2479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13761_ clknet_leaf_47_clk _00992_ net1199 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[749\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12284__A1 net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10973_ net84 net1046 net85 vssd1 vssd1 vccd1 vccd1 _05700_ sky130_fd_sc_hd__or3b_1
XANTENNA__09685__C1 _04072_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12712_ final_design.VGA_data_control.v_count\[3\] _06351_ vssd1 vssd1 vccd1 vccd1
+ _06353_ sky130_fd_sc_hd__nand2_1
XANTENNA__07386__S1 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08583__S0 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13692_ clknet_leaf_2_clk _00923_ net1064 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[680\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08655__A _01566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12643_ final_design.VGA_data_control.ready_data\[9\] net1019 net974 final_design.data_from_mem\[9\]
+ vssd1 vssd1 vccd1 vccd1 _06309_ sky130_fd_sc_hd__a22o_1
XFILLER_0_66_852 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12587__A2 net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07138__S1 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12574_ net1052 final_design.uart.working_data\[7\] vssd1 vssd1 vccd1 vccd1 _06292_
+ sky130_fd_sc_hd__and2_1
XANTENNA__09452__A2 net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11525_ net2459 _06120_ _06122_ net434 vssd1 vssd1 vccd1 vccd1 _00392_ sky130_fd_sc_hd__a22o_1
XANTENNA__06897__S0 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12464__X _06283_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12907__CLK clknet_leaf_61_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12339__A2 net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14244_ net1298 vssd1 vssd1 vccd1 vccd1 gpio_out[22] sky130_fd_sc_hd__buf_2
X_11456_ net238 net638 vssd1 vssd1 vccd1 vccd1 _06101_ sky130_fd_sc_hd__and2_1
XFILLER_0_68_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10407_ net1436 net1030 _05186_ net246 vssd1 vssd1 vccd1 vccd1 _00145_ sky130_fd_sc_hd__a22o_1
X_14175_ clknet_leaf_21_clk _01349_ net1161 vssd1 vssd1 vccd1 vccd1 final_design.VGA_adr\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12116__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10425__A _03096_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11387_ net652 _06070_ _06072_ _05843_ vssd1 vssd1 vccd1 vccd1 _06073_ sky130_fd_sc_hd__a31o_1
XFILLER_0_0_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13126_ clknet_leaf_50_clk _00357_ net1168 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[114\]
+ sky130_fd_sc_hd__dfrtp_1
X_10338_ net1503 net1009 net986 final_design.data_from_mem\[23\] vssd1 vssd1 vccd1
+ vccd1 _00095_ sky130_fd_sc_hd__a22o_1
XFILLER_0_24_1662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13057_ clknet_leaf_49_clk _00288_ net1198 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[45\]
+ sky130_fd_sc_hd__dfrtp_1
X_10269_ net1812 _05129_ _05131_ vssd1 vssd1 vccd1 vccd1 _00023_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07518__A2 _01690_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07734__A net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12511__A2 net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12008_ _06210_ net287 net402 net2272 vssd1 vssd1 vccd1 vccd1 _00739_ sky130_fd_sc_hd__a22o_1
XANTENNA__09912__B1 net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12275__A1 net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13959_ clknet_leaf_61_clk _01190_ net1124 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[947\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09140__A1 _04058_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06500_ net762 _01450_ vssd1 vssd1 vccd1 vccd1 _01451_ sky130_fd_sc_hd__or2_1
X_07480_ _02364_ _02429_ _02362_ vssd1 vssd1 vccd1 vccd1 _02431_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_53_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06431_ net51 vssd1 vssd1 vccd1 vccd1 _01386_ sky130_fd_sc_hd__inv_2
XANTENNA__11703__B net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11235__C1 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09150_ _03628_ _04053_ vssd1 vssd1 vccd1 vccd1 _04069_ sky130_fd_sc_hd__nor2_4
XFILLER_0_51_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08101_ net716 _03051_ vssd1 vssd1 vccd1 vccd1 _03052_ sky130_fd_sc_hd__or2_1
X_09081_ _03705_ _03721_ vssd1 vssd1 vccd1 vccd1 _04006_ sky130_fd_sc_hd__xor2_1
XFILLER_0_32_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13832__CLK clknet_leaf_41_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08032_ _02979_ _02980_ _02981_ _02982_ net679 net699 vssd1 vssd1 vccd1 vccd1 _02983_
+ sky130_fd_sc_hd__mux4_1
Xinput50 mem_adr_start[22] vssd1 vssd1 vccd1 vccd1 net50 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput61 mem_adr_start[3] vssd1 vssd1 vccd1 vccd1 net61 sky130_fd_sc_hd__clkbuf_1
Xinput72 memory_size[13] vssd1 vssd1 vccd1 vccd1 net72 sky130_fd_sc_hd__buf_1
Xhold801 final_design.cpu.reg_window\[142\] vssd1 vssd1 vccd1 vccd1 net2143 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkload42_A clknet_leaf_34_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold812 final_design.cpu.reg_window\[273\] vssd1 vssd1 vccd1 vccd1 net2154 sky130_fd_sc_hd__dlygate4sd3_1
Xinput83 memory_size[23] vssd1 vssd1 vccd1 vccd1 net83 sky130_fd_sc_hd__clkbuf_2
Xhold823 final_design.cpu.reg_window\[865\] vssd1 vssd1 vccd1 vccd1 net2165 sky130_fd_sc_hd__dlygate4sd3_1
Xinput94 memory_size[4] vssd1 vssd1 vccd1 vccd1 net94 sky130_fd_sc_hd__buf_1
Xhold834 final_design.cpu.reg_window\[257\] vssd1 vssd1 vccd1 vccd1 net2176 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09600__C1 _04109_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold845 final_design.cpu.reg_window\[206\] vssd1 vssd1 vccd1 vccd1 net2187 sky130_fd_sc_hd__dlygate4sd3_1
Xhold856 final_design.cpu.reg_window\[1008\] vssd1 vssd1 vccd1 vccd1 net2198 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08954__A1 _03655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold867 final_design.cpu.reg_window\[326\] vssd1 vssd1 vccd1 vccd1 net2209 sky130_fd_sc_hd__dlygate4sd3_1
Xhold878 final_design.cpu.reg_window\[551\] vssd1 vssd1 vccd1 vccd1 net2220 sky130_fd_sc_hd__dlygate4sd3_1
Xhold889 final_design.cpu.reg_window\[995\] vssd1 vssd1 vccd1 vccd1 net2231 sky130_fd_sc_hd__dlygate4sd3_1
X_09983_ _04898_ _04901_ vssd1 vssd1 vccd1 vccd1 _04902_ sky130_fd_sc_hd__nand2_1
XANTENNA__13982__CLK clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08934_ _02464_ net625 _03872_ _03875_ vssd1 vssd1 vccd1 vccd1 _03876_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout1012_A _05166_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07644__A net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12502__A2 net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08865_ final_design.CPU_instr_adr\[29\] _01538_ vssd1 vssd1 vccd1 vccd1 _03814_
+ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_4_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout472_A net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11710__B1 net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13212__CLK clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08182__A2 net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07816_ net615 _02763_ _02764_ _01657_ vssd1 vssd1 vccd1 vccd1 _02767_ sky130_fd_sc_hd__a211oi_2
X_08796_ _03679_ _03740_ _03743_ _03744_ _03746_ vssd1 vssd1 vccd1 vccd1 _03747_ sky130_fd_sc_hd__o41a_1
XFILLER_0_58_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07747_ _02685_ _02686_ _02697_ net877 vssd1 vssd1 vccd1 vccd1 _02698_ sky130_fd_sc_hd__a22oi_4
XANTENNA_fanout737_A net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout358_X net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_2310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07678_ final_design.cpu.reg_window\[734\] final_design.cpu.reg_window\[766\] net853
+ vssd1 vssd1 vccd1 vccd1 _02629_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_62_2321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06547__X _01498_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_2955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_2332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_2966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_0_Right_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13362__CLK clknet_leaf_39_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_2977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09417_ _01535_ _01566_ _01596_ _01626_ net453 net462 vssd1 vssd1 vccd1 vccd1 _04336_
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_66_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11613__B net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06629_ final_design.cpu.reg_window\[155\] final_design.cpu.reg_window\[187\] net947
+ vssd1 vssd1 vccd1 vccd1 _01580_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_1829 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout904_A net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08317__S0 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09348_ net481 net470 net527 vssd1 vssd1 vccd1 vccd1 _04267_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11777__B1 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06879__S0 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09279_ _04177_ _04197_ vssd1 vssd1 vccd1 vccd1 _04198_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_30_1187 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11310_ net663 _03890_ net738 vssd1 vssd1 vccd1 vccd1 _06005_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_79_2895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12290_ net581 _06220_ net514 net370 net2094 vssd1 vssd1 vccd1 vccd1 _01005_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_56_2114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_2125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_2759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_2136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11241_ net662 _03955_ net736 vssd1 vssd1 vccd1 vccd1 _05944_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_26_Left_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12741__A2 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11172_ net646 net565 net226 vssd1 vssd1 vccd1 vccd1 _05884_ sky130_fd_sc_hd__and3_1
X_10123_ final_design.VGA_data_control.v_count\[0\] net1051 final_design.VGA_data_control.v_count\[2\]
+ final_design.VGA_data_control.v_count\[3\] vssd1 vssd1 vccd1 vccd1 _05031_ sky130_fd_sc_hd__and4_1
XFILLER_0_41_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13748__RESET_B net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input33_A DAT_I[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10054_ net68 _04940_ _04679_ vssd1 vssd1 vccd1 vccd1 _04973_ sky130_fd_sc_hd__a21bo_1
XANTENNA__07554__A net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07056__S0 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_1879 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13813_ clknet_leaf_57_clk _01044_ net1145 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[801\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13705__CLK clknet_leaf_36_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_35_Left_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11363__X _06052_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07359__S1 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13744_ clknet_leaf_36_clk _00975_ net1236 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[732\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06457__X _01410_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10956_ _01361_ _03859_ net1059 vssd1 vssd1 vccd1 vccd1 _05684_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_1043 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13675_ clknet_leaf_53_clk _00906_ net1187 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[663\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07684__B2 net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10887_ net962 _05617_ vssd1 vssd1 vccd1 vccd1 _05618_ sky130_fd_sc_hd__or2_1
XFILLER_0_39_863 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13855__CLK clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12626_ _06300_ net1394 net980 vssd1 vssd1 vccd1 vccd1 _01315_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_14_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12557_ _06220_ net355 net325 net2216 vssd1 vssd1 vccd1 vccd1 _01261_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07288__X _02239_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11508_ net1674 net237 net522 vssd1 vssd1 vccd1 vccd1 _00377_ sky130_fd_sc_hd__mux2_1
XANTENNA__07531__S1 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12488_ _06148_ net352 net333 net2051 vssd1 vssd1 vccd1 vccd1 _01194_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_44_Left_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold108 final_design.VGA_data_control.data_to_VGA\[16\] vssd1 vssd1 vccd1 vccd1 net1450
+ sky130_fd_sc_hd__dlygate4sd3_1
X_14227_ net1281 vssd1 vssd1 vccd1 vccd1 gpio_out[5] sky130_fd_sc_hd__buf_2
Xhold119 net142 vssd1 vssd1 vccd1 vccd1 net1461 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11439_ net2032 net180 net312 vssd1 vssd1 vccd1 vccd1 _00336_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_1773 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14158_ clknet_leaf_14_clk _01332_ net1110 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.data_to_VGA\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11940__B1 net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13235__CLK clknet_leaf_39_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13109_ clknet_leaf_7_clk _00340_ net1145 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[97\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11538__X _06125_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06980_ final_design.cpu.reg_window\[720\] final_design.cpu.reg_window\[752\] net923
+ vssd1 vssd1 vccd1 vccd1 _01931_ sky130_fd_sc_hd__mux2_1
X_14089_ clknet_leaf_25_clk _01286_ net1155 vssd1 vssd1 vccd1 vccd1 final_design.reqhand.instruction\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08149__C1 net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12496__A1 _06156_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11299__A2 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1170 net1176 vssd1 vssd1 vccd1 vccd1 net1170 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09361__A1 _04046_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1181 net1182 vssd1 vssd1 vccd1 vccd1 net1181 sky130_fd_sc_hd__clkbuf_4
X_08650_ net605 _02668_ _02643_ _01597_ vssd1 vssd1 vccd1 vccd1 _03601_ sky130_fd_sc_hd__o211a_1
Xfanout1192 net1197 vssd1 vssd1 vccd1 vccd1 net1192 sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_53_Left_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13385__CLK clknet_leaf_36_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07601_ final_design.cpu.reg_window\[93\] final_design.cpu.reg_window\[125\] net870
+ vssd1 vssd1 vccd1 vccd1 _02552_ sky130_fd_sc_hd__mux2_1
XANTENNA__12248__A1 net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08581_ final_design.cpu.reg_window\[192\] final_design.cpu.reg_window\[224\] net814
+ vssd1 vssd1 vccd1 vccd1 _03532_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_1733 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09113__A1 _02419_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08547__S0 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13000__RESET_B net1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07532_ final_design.cpu.reg_window\[95\] final_design.cpu.reg_window\[127\] net937
+ vssd1 vssd1 vccd1 vccd1 _02483_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1777 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09664__A2 _04309_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07463_ final_design.cpu.reg_window\[640\] final_design.cpu.reg_window\[672\] net908
+ vssd1 vssd1 vccd1 vccd1 _02414_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09202_ net496 net492 _04099_ _04120_ vssd1 vssd1 vccd1 vccd1 _04121_ sky130_fd_sc_hd__or4_1
X_06414_ final_design.VGA_data_control.v_count\[8\] vssd1 vssd1 vccd1 vccd1 _01369_
+ sky130_fd_sc_hd__inv_2
XANTENNA_wire695_X net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07394_ final_design.cpu.reg_window\[962\] final_design.cpu.reg_window\[994\] net913
+ vssd1 vssd1 vccd1 vccd1 _02345_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09133_ _03607_ _04051_ _02641_ vssd1 vssd1 vccd1 vccd1 _04052_ sky130_fd_sc_hd__o21a_1
XFILLER_0_60_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout220_A net221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_62_Left_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout318_A _04117_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09064_ _02215_ _02437_ vssd1 vssd1 vccd1 vccd1 _03991_ sky130_fd_sc_hd__or2_1
XANTENNA__14010__CLK clknet_leaf_63_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08015_ _01853_ net603 vssd1 vssd1 vccd1 vccd1 _02966_ sky130_fd_sc_hd__nand2_1
Xhold620 final_design.cpu.reg_window\[402\] vssd1 vssd1 vccd1 vccd1 net1962 sky130_fd_sc_hd__dlygate4sd3_1
Xhold631 final_design.cpu.reg_window\[136\] vssd1 vssd1 vccd1 vccd1 net1973 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1227_A net1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold642 final_design.cpu.reg_window\[141\] vssd1 vssd1 vccd1 vccd1 net1984 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_2601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold653 final_design.cpu.reg_window\[600\] vssd1 vssd1 vccd1 vccd1 net1995 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_70_2612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07286__S0 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold664 final_design.cpu.reg_window\[179\] vssd1 vssd1 vccd1 vccd1 net2006 sky130_fd_sc_hd__dlygate4sd3_1
Xhold675 final_design.cpu.reg_window\[947\] vssd1 vssd1 vccd1 vccd1 net2017 sky130_fd_sc_hd__dlygate4sd3_1
Xhold686 final_design.cpu.reg_window\[384\] vssd1 vssd1 vccd1 vccd1 net2028 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout687_A net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold697 final_design.cpu.reg_window\[531\] vssd1 vssd1 vccd1 vccd1 net2039 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14160__CLK clknet_leaf_19_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09966_ _04725_ _04750_ _04768_ _04884_ vssd1 vssd1 vccd1 vccd1 _04885_ sky130_fd_sc_hd__and4_1
XANTENNA__06689__S net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08917_ final_design.CPU_instr_adr\[24\] net1014 _03858_ _03860_ vssd1 vssd1 vccd1
+ vccd1 _00235_ sky130_fd_sc_hd__a22o_1
XANTENNA__13728__CLK clknet_leaf_11_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_71_Left_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09897_ net470 _04815_ net482 vssd1 vssd1 vccd1 vccd1 _04816_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout854_A net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08848_ final_design.CPU_instr_adr\[26\] _03798_ vssd1 vssd1 vccd1 vccd1 _03799_
+ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_68_2530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_3_1_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_2541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10823__A1_N net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_2405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08779_ _03692_ _03694_ _03729_ vssd1 vssd1 vccd1 vccd1 _03730_ sky130_fd_sc_hd__and3_1
XFILLER_0_36_1330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10810_ net1005 _05544_ vssd1 vssd1 vccd1 vccd1 _05545_ sky130_fd_sc_hd__nor2_1
XANTENNA__13878__CLK clknet_leaf_58_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11790_ net2240 net412 net276 _05973_ vssd1 vssd1 vccd1 vccd1 _00546_ sky130_fd_sc_hd__a22o_1
XANTENNA__11998__B1 net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10741_ net40 _05456_ _05460_ vssd1 vssd1 vccd1 vccd1 _05479_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08863__B1 net1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07761__S1 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13460_ clknet_leaf_10_clk _00691_ net1102 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[448\]
+ sky130_fd_sc_hd__dfrtp_1
X_10672_ final_design.CPU_instr_adr\[11\] net1042 net802 vssd1 vssd1 vccd1 vccd1 _05413_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_48_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13108__CLK clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_80_Left_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_11_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12411_ net207 net553 net499 net338 net1693 vssd1 vssd1 vccd1 vccd1 _01121_ sky130_fd_sc_hd__a32o_1
XFILLER_0_63_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10674__S net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13391_ clknet_leaf_42_clk _00622_ net1225 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[379\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12411__A1 net207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09812__C1 net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_20_clk clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_20_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_69_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12342_ _06232_ net500 net361 net2491 vssd1 vssd1 vccd1 vccd1 _01054_ sky130_fd_sc_hd__a22o_1
XANTENNA__08144__S net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13258__CLK clknet_leaf_60_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12273_ net556 _06203_ net502 net368 net1885 vssd1 vssd1 vccd1 vccd1 _00988_ sky130_fd_sc_hd__a32o_1
XFILLER_0_62_1913 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14012_ clknet_leaf_3_clk _01243_ net1079 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[1000\]
+ sky130_fd_sc_hd__dfrtp_1
X_11224_ net426 net556 _05929_ net314 net2038 vssd1 vssd1 vccd1 vccd1 _00284_ sky130_fd_sc_hd__a32o_1
X_11155_ _05839_ _05866_ vssd1 vssd1 vccd1 vccd1 _05869_ sky130_fd_sc_hd__nand2_8
XTAP_TAPCELL_ROW_8_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10106_ final_design.VGA_data_control.v_count\[0\] _05017_ final_design.VGA_data_control.v_count\[1\]
+ vssd1 vssd1 vccd1 vccd1 _05021_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_8_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07029__S0 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11086_ final_design.CPU_instr_adr\[30\] _03811_ net1059 vssd1 vssd1 vccd1 vccd1
+ _05808_ sky130_fd_sc_hd__mux2_1
X_10037_ _04955_ vssd1 vssd1 vccd1 vccd1 _04956_ sky130_fd_sc_hd__inv_2
XANTENNA__11150__A1 _04805_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11988_ _06190_ net285 net407 net1620 vssd1 vssd1 vccd1 vccd1 _00721_ sky130_fd_sc_hd__a22o_1
XANTENNA__11989__B1 net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09646__A2 _04559_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13727_ clknet_leaf_8_clk _00958_ net1131 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[715\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10939_ _05645_ _05662_ _05663_ vssd1 vssd1 vccd1 vccd1 _05667_ sky130_fd_sc_hd__or3_1
XFILLER_0_14_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09498__X _04417_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13658_ clknet_leaf_64_clk _00889_ net1075 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[646\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09939__A net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14033__CLK clknet_leaf_34_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12609_ net1578 net998 net984 final_design.data_from_mem\[27\] vssd1 vssd1 vccd1
+ vccd1 _01302_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_26_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13589_ clknet_leaf_58_clk _00820_ net1133 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[577\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_11_clk clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_11_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_30_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14183__CLK clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10716__A1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11913__A0 net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10716__B2 _04036_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_6_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout407 _06255_ vssd1 vssd1 vccd1 vccd1 net407 sky130_fd_sc_hd__clkbuf_4
X_09820_ _03295_ _03569_ _03575_ net321 vssd1 vssd1 vccd1 vccd1 _04739_ sky130_fd_sc_hd__a211o_1
Xfanout418 net419 vssd1 vssd1 vccd1 vccd1 net418 sky130_fd_sc_hd__clkbuf_8
XANTENNA__12304__S net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout429 net430 vssd1 vssd1 vccd1 vccd1 net429 sky130_fd_sc_hd__buf_4
X_09751_ net491 _04222_ _04261_ _04667_ _04669_ vssd1 vssd1 vccd1 vccd1 _04670_ sky130_fd_sc_hd__o311a_1
X_06963_ final_design.cpu.reg_window\[272\] final_design.cpu.reg_window\[304\] net925
+ vssd1 vssd1 vccd1 vccd1 _01914_ sky130_fd_sc_hd__mux2_1
X_08702_ _03635_ _03645_ _03650_ _03652_ net731 vssd1 vssd1 vccd1 vccd1 _03653_ sky130_fd_sc_hd__o311a_1
X_09682_ _03163_ net443 vssd1 vssd1 vccd1 vccd1 _04601_ sky130_fd_sc_hd__nor2_1
X_06894_ final_design.cpu.reg_window\[659\] final_design.cpu.reg_window\[691\] net902
+ vssd1 vssd1 vccd1 vccd1 _01845_ sky130_fd_sc_hd__mux2_1
X_08633_ _03166_ _03581_ _03583_ vssd1 vssd1 vccd1 vccd1 _03584_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_59_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11692__A2 net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08737__B _02097_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout268_A net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11444__A net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07991__S1 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08564_ _02394_ net608 vssd1 vssd1 vccd1 vccd1 _03515_ sky130_fd_sc_hd__nor2_1
XFILLER_0_76_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11163__B net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07515_ _01723_ _01725_ vssd1 vssd1 vccd1 vccd1 _02466_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_1913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08495_ final_design.cpu.reg_window\[579\] final_design.cpu.reg_window\[611\] net825
+ vssd1 vssd1 vccd1 vccd1 _03446_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12641__B2 final_design.data_from_mem\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout435_A net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07446_ final_design.cpu.reg_window\[256\] final_design.cpu.reg_window\[288\] net909
+ vssd1 vssd1 vccd1 vccd1 _02397_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09201__X _04120_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_21_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout223_X net223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07377_ final_design.reqhand.instruction\[10\] net972 _02327_ vssd1 vssd1 vccd1 vccd1
+ _02328_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout602_A net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06871__A2 _01498_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13400__CLK clknet_leaf_63_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_2810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09116_ net995 net992 net1040 vssd1 vssd1 vccd1 vccd1 _04035_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_60_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10507__B net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1356 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09047_ _03728_ _03975_ vssd1 vssd1 vccd1 vccd1 _03976_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_44_1643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold450 final_design.cpu.reg_window\[69\] vssd1 vssd1 vccd1 vccd1 net1792 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout971_A _01415_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13550__CLK clknet_leaf_44_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold461 final_design.cpu.reg_window\[700\] vssd1 vssd1 vccd1 vccd1 net1803 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout592_X net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold472 final_design.cpu.reg_window\[919\] vssd1 vssd1 vccd1 vccd1 net1814 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09573__A1 net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold483 final_design.cpu.reg_window\[170\] vssd1 vssd1 vccd1 vccd1 net1825 sky130_fd_sc_hd__dlygate4sd3_1
Xhold494 final_design.cpu.reg_window\[187\] vssd1 vssd1 vccd1 vccd1 net1836 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_1717 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout930 net931 vssd1 vssd1 vccd1 vccd1 net930 sky130_fd_sc_hd__clkbuf_4
Xfanout941 net942 vssd1 vssd1 vccd1 vccd1 net941 sky130_fd_sc_hd__clkbuf_4
X_09949_ _04112_ _04867_ _04443_ vssd1 vssd1 vccd1 vccd1 _04868_ sky130_fd_sc_hd__o21ba_1
Xfanout952 net953 vssd1 vssd1 vccd1 vccd1 net952 sky130_fd_sc_hd__buf_2
Xfanout963 _04036_ vssd1 vssd1 vccd1 vccd1 net963 sky130_fd_sc_hd__clkbuf_2
Xfanout974 _06299_ vssd1 vssd1 vccd1 vccd1 net974 sky130_fd_sc_hd__buf_2
XANTENNA__09590__Y _04509_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout985 _06296_ vssd1 vssd1 vccd1 vccd1 net985 sky130_fd_sc_hd__clkbuf_2
X_12960_ clknet_leaf_32_clk _00198_ net1233 vssd1 vssd1 vccd1 vccd1 net118 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_77_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout996 net997 vssd1 vssd1 vccd1 vccd1 net996 sky130_fd_sc_hd__buf_2
Xhold1150 final_design.cpu.reg_window\[555\] vssd1 vssd1 vccd1 vccd1 net2492 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_77_1463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09523__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11911_ net191 net1909 net274 vssd1 vssd1 vccd1 vccd1 _00651_ sky130_fd_sc_hd__mux2_1
Xhold1161 final_design.cpu.reg_window\[116\] vssd1 vssd1 vccd1 vccd1 net2503 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1172 final_design.cpu.reg_window\[125\] vssd1 vssd1 vccd1 vccd1 net2514 sky130_fd_sc_hd__dlygate4sd3_1
X_12891_ clknet_leaf_17_clk _00129_ net1113 vssd1 vssd1 vccd1 vccd1 final_design.data_from_mem\[25\]
+ sky130_fd_sc_hd__dfrtp_4
Xhold1183 final_design.CPU_instr_adr\[4\] vssd1 vssd1 vccd1 vccd1 net2525 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1194 final_design.cpu.reg_window\[308\] vssd1 vssd1 vccd1 vccd1 net2536 sky130_fd_sc_hd__dlygate4sd3_1
X_11842_ net176 net2350 net266 vssd1 vssd1 vccd1 vccd1 _00594_ sky130_fd_sc_hd__mux2_1
XANTENNA__08139__S net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14056__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1160 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_0_191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11773_ net2520 net413 _06229_ net428 vssd1 vssd1 vccd1 vccd1 _00533_ sky130_fd_sc_hd__a22o_1
XFILLER_0_71_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13512_ clknet_leaf_41_clk _00743_ net1224 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[500\]
+ sky130_fd_sc_hd__dfrtp_1
X_10724_ net729 _04613_ net249 vssd1 vssd1 vccd1 vccd1 _05462_ sky130_fd_sc_hd__and3_1
XFILLER_0_49_991 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_22_clk_X clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13443_ clknet_leaf_1_clk _00674_ net1071 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[431\]
+ sky130_fd_sc_hd__dfrtp_1
X_10655_ net965 _05396_ vssd1 vssd1 vccd1 vccd1 _05397_ sky130_fd_sc_hd__nand2_1
XFILLER_0_67_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13080__CLK clknet_leaf_62_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkload17 clknet_leaf_17_clk vssd1 vssd1 vccd1 vccd1 clkload17/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_23_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13374_ clknet_leaf_9_clk _00605_ net1103 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[362\]
+ sky130_fd_sc_hd__dfrtp_1
X_10586_ net97 final_design.VGA_adr\[5\] vssd1 vssd1 vccd1 vccd1 _05331_ sky130_fd_sc_hd__nand2_1
Xclkload28 clknet_leaf_49_clk vssd1 vssd1 vccd1 vccd1 clkload28/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__10417__B _05190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload39 clknet_leaf_30_clk vssd1 vssd1 vccd1 vccd1 clkload39/Y sky130_fd_sc_hd__inv_6
X_12325_ net2285 net183 net366 vssd1 vssd1 vccd1 vccd1 _01039_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_37_clk_X clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12256_ net577 _06185_ _06264_ net374 net2090 vssd1 vssd1 vccd1 vccd1 _00972_ sky130_fd_sc_hd__a32o_1
XANTENNA__06911__A net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_16 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11207_ _03615_ _05913_ vssd1 vssd1 vccd1 vccd1 _05914_ sky130_fd_sc_hd__nor2_2
X_12187_ net2317 net192 net382 vssd1 vssd1 vccd1 vccd1 _00906_ sky130_fd_sc_hd__mux2_1
XANTENNA__12124__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11138_ _01495_ _03614_ vssd1 vssd1 vccd1 vccd1 _05853_ sky130_fd_sc_hd__nor2_1
XANTENNA__07670__S0 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11069_ _01388_ _05790_ vssd1 vssd1 vccd1 vccd1 _05792_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_30_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_0_clk clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_0_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_30_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_3003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_3014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_3025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_3036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07878__A1 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11674__A2 net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_3047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1861 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06550__A1 final_design.data_from_mem\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_28_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07300_ final_design.cpu.reg_window\[453\] final_design.cpu.reg_window\[485\] net919
+ vssd1 vssd1 vccd1 vccd1 _02251_ sky130_fd_sc_hd__mux2_1
XANTENNA__13423__CLK clknet_leaf_38_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08280_ _03195_ _03196_ _03227_ _03228_ vssd1 vssd1 vccd1 vccd1 _03231_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_24_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1299 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07231_ _02178_ _02179_ _02180_ _02181_ net766 net786 vssd1 vssd1 vccd1 vccd1 _02182_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__11711__B net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06805__B _01503_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07162_ net758 _02112_ net745 vssd1 vssd1 vccd1 vccd1 _02113_ sky130_fd_sc_hd__o21a_1
XANTENNA__13573__CLK clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07093_ net757 _02043_ vssd1 vssd1 vccd1 vccd1 _02044_ sky130_fd_sc_hd__or2_1
XFILLER_0_48_1064 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_880 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09555__A1 net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout204 _05989_ vssd1 vssd1 vccd1 vccd1 net204 sky130_fd_sc_hd__clkbuf_2
XANTENNA__12034__S net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout215 _05941_ vssd1 vssd1 vccd1 vccd1 net215 sky130_fd_sc_hd__buf_2
Xfanout226 net227 vssd1 vssd1 vccd1 vccd1 net226 sky130_fd_sc_hd__clkbuf_2
Xfanout237 net238 vssd1 vssd1 vccd1 vccd1 net237 sky130_fd_sc_hd__clkbuf_2
X_09803_ net321 _04721_ vssd1 vssd1 vccd1 vccd1 _04722_ sky130_fd_sc_hd__nor2_1
Xfanout248 net249 vssd1 vssd1 vccd1 vccd1 net248 sky130_fd_sc_hd__buf_4
X_07995_ final_design.cpu.reg_window\[144\] final_design.cpu.reg_window\[176\] net846
+ vssd1 vssd1 vccd1 vccd1 _02946_ sky130_fd_sc_hd__mux2_1
Xfanout259 _03654_ vssd1 vssd1 vccd1 vccd1 net259 sky130_fd_sc_hd__buf_2
XANTENNA_fanout385_A _06266_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09734_ _04124_ _04652_ _04651_ net263 vssd1 vssd1 vccd1 vccd1 _04653_ sky130_fd_sc_hd__o211ai_2
X_06946_ final_design.cpu.reg_window\[849\] final_design.cpu.reg_window\[881\] net925
+ vssd1 vssd1 vccd1 vccd1 _01897_ sky130_fd_sc_hd__mux2_1
XANTENNA__09858__A2 net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14079__CLK clknet_leaf_19_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07652__A _01570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09665_ net319 _04301_ _04305_ net320 vssd1 vssd1 vccd1 vccd1 _04584_ sky130_fd_sc_hd__a22o_1
X_06877_ final_design.cpu.reg_window\[467\] final_design.cpu.reg_window\[499\] net911
+ vssd1 vssd1 vccd1 vccd1 _01828_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout552_A _01686_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06539__Y _01490_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08616_ _03359_ _03564_ _03565_ _03327_ _03566_ vssd1 vssd1 vccd1 vccd1 _03567_ sky130_fd_sc_hd__a221o_1
X_09596_ net471 _04240_ net481 vssd1 vssd1 vccd1 vccd1 _04515_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_38_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08547_ _03494_ _03495_ _03496_ _03497_ net681 net699 vssd1 vssd1 vccd1 vccd1 _03498_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_38_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout340_X net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout817_A net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_1721 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout438_X net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08478_ final_design.cpu.reg_window\[451\] final_design.cpu.reg_window\[483\] net823
+ vssd1 vssd1 vccd1 vccd1 _03429_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13916__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11621__B net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07429_ final_design.cpu.reg_window\[897\] final_design.cpu.reg_window\[929\] net914
+ vssd1 vssd1 vccd1 vccd1 _02380_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10440_ _02830_ net592 vssd1 vssd1 vccd1 vccd1 _05204_ sky130_fd_sc_hd__nor2_1
XFILLER_0_66_1120 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10371_ net14 net1024 net1006 final_design.data_from_mem\[20\] vssd1 vssd1 vccd1
+ vccd1 _00124_ sky130_fd_sc_hd__o22a_1
XANTENNA__12940__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12110_ net1877 net205 net388 vssd1 vssd1 vccd1 vccd1 _00834_ sky130_fd_sc_hd__mux2_1
XANTENNA__08422__S net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13090_ clknet_leaf_3_clk _00321_ net1068 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[78\]
+ sky130_fd_sc_hd__dfrtp_1
X_12041_ net1728 net208 net396 vssd1 vssd1 vccd1 vccd1 _00769_ sky130_fd_sc_hd__mux2_1
XFILLER_0_40_1304 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold280 final_design.cpu.reg_window\[163\] vssd1 vssd1 vccd1 vccd1 net1622 sky130_fd_sc_hd__dlygate4sd3_1
Xhold291 final_design.cpu.reg_window\[184\] vssd1 vssd1 vccd1 vccd1 net1633 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11353__A1 _01660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12550__B1 net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11353__B2 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout760 _01426_ vssd1 vssd1 vccd1 vccd1 net760 sky130_fd_sc_hd__buf_4
Xfanout771 _01422_ vssd1 vssd1 vccd1 vccd1 net771 sky130_fd_sc_hd__buf_4
Xfanout782 _01419_ vssd1 vssd1 vccd1 vccd1 net782 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11105__A1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13992_ clknet_leaf_42_clk _01223_ net1224 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[980\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout793 net795 vssd1 vssd1 vccd1 vccd1 net793 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11105__B2 net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08506__C1 _02326_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12943_ clknet_leaf_29_clk _00181_ net1193 vssd1 vssd1 vccd1 vccd1 net131 sky130_fd_sc_hd__dfrtp_1
XANTENNA__11656__A2 net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08010__X _02961_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13446__CLK clknet_leaf_51_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_64_clk_A clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12874_ clknet_leaf_15_clk _00112_ net1094 vssd1 vssd1 vccd1 vccd1 final_design.data_from_mem\[8\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_62_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09157__S0 net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11825_ net207 net2071 net264 vssd1 vssd1 vccd1 vccd1 _00577_ sky130_fd_sc_hd__mux2_1
XANTENNA__12605__B2 final_design.data_from_mem\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10616__B1 net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09482__A0 net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11756_ net197 net2160 net418 vssd1 vssd1 vccd1 vccd1 _00519_ sky130_fd_sc_hd__mux2_1
XANTENNA__12081__A2 net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13596__CLK clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10707_ net72 net1043 vssd1 vssd1 vccd1 vccd1 _05446_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_42_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12119__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11687_ net220 net626 vssd1 vssd1 vccd1 vccd1 _06202_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_42_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13426_ clknet_leaf_38_clk _00657_ net1190 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[414\]
+ sky130_fd_sc_hd__dfrtp_1
X_10638_ net961 _05380_ vssd1 vssd1 vccd1 vccd1 _05381_ sky130_fd_sc_hd__or2_1
XFILLER_0_29_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10147__B net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10919__B2 net1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10654__A1_N net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13357_ clknet_leaf_44_clk _00588_ net1209 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[345\]
+ sky130_fd_sc_hd__dfrtp_1
X_10569_ _05288_ _05313_ vssd1 vssd1 vccd1 vccd1 _05315_ sky130_fd_sc_hd__or2_1
XFILLER_0_23_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10395__A2 net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12308_ net1811 net214 net364 vssd1 vssd1 vccd1 vccd1 _01022_ sky130_fd_sc_hd__mux2_1
X_13288_ clknet_leaf_41_clk _00519_ net1224 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[276\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10434__Y _05201_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12239_ net557 _06169_ net502 net372 net1502 vssd1 vssd1 vccd1 vccd1 _00956_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_36_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11344__A1 final_design.data_from_mem\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_17_clk_A clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12541__B1 net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07643__S0 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06800_ final_design.reqhand.instruction\[22\] net971 vssd1 vssd1 vccd1 vccd1 _01751_
+ sky130_fd_sc_hd__or2_1
X_07780_ _02718_ _02719_ _02730_ net877 vssd1 vssd1 vccd1 vccd1 _02731_ sky130_fd_sc_hd__a22oi_4
XFILLER_0_36_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput4 DAT_I[11] vssd1 vssd1 vccd1 vccd1 net4 sky130_fd_sc_hd__clkbuf_1
X_06731_ final_design.cpu.reg_window\[728\] final_design.cpu.reg_window\[760\] net942
+ vssd1 vssd1 vccd1 vccd1 _01682_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_1322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1907 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09450_ _02767_ net445 net443 vssd1 vssd1 vccd1 vccd1 _04369_ sky130_fd_sc_hd__o21a_1
X_06662_ net753 _01606_ net748 vssd1 vssd1 vccd1 vccd1 _01613_ sky130_fd_sc_hd__o21a_1
XFILLER_0_8_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08401_ net875 _03351_ _03340_ _03339_ vssd1 vssd1 vccd1 vccd1 _03352_ sky130_fd_sc_hd__o2bb2a_2
XANTENNA__13939__CLK clknet_leaf_41_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09381_ net545 net544 net542 net541 net459 net469 vssd1 vssd1 vccd1 vccd1 _04300_
+ sky130_fd_sc_hd__mux4_2
X_06593_ final_design.cpu.reg_window\[92\] final_design.cpu.reg_window\[124\] net940
+ vssd1 vssd1 vccd1 vccd1 _01544_ sky130_fd_sc_hd__mux2_1
XANTENNA__09699__S1 net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08332_ final_design.cpu.reg_window\[584\] final_design.cpu.reg_window\[616\] net807
+ vssd1 vssd1 vccd1 vccd1 _03283_ sky130_fd_sc_hd__mux2_1
XANTENNA__07079__A2 _02029_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1705 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08263_ final_design.cpu.reg_window\[778\] final_design.cpu.reg_window\[810\] net817
+ vssd1 vssd1 vccd1 vccd1 _03214_ sky130_fd_sc_hd__mux2_1
XANTENNA__11280__B1 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12029__S net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1749 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07214_ final_design.cpu.reg_window\[200\] final_design.cpu.reg_window\[232\] net893
+ vssd1 vssd1 vccd1 vccd1 _02165_ sky130_fd_sc_hd__mux2_1
X_12784__15 clknet_leaf_28_clk vssd1 vssd1 vccd1 vccd1 net1325 sky130_fd_sc_hd__inv_2
X_08194_ final_design.cpu.reg_window\[142\] final_design.cpu.reg_window\[174\] net812
+ vssd1 vssd1 vccd1 vccd1 _03145_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_1905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07145_ _01463_ net740 _02095_ vssd1 vssd1 vccd1 vccd1 _02096_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout300_A net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1042_A _01371_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11583__A1 net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13319__CLK clknet_leaf_59_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07076_ net1041 net993 net990 final_design.reqhand.instruction\[13\] vssd1 vssd1
+ vccd1 vccd1 _02027_ sky130_fd_sc_hd__a31o_1
XFILLER_0_77_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12532__B1 net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1072 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout290_X net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout767_A net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout388_X net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13469__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07978_ net879 _02928_ _02917_ _02911_ vssd1 vssd1 vccd1 vccd1 _02929_ sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_57_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09717_ net727 _04626_ _04630_ _04634_ vssd1 vssd1 vccd1 vccd1 _04636_ sky130_fd_sc_hd__or4b_1
XANTENNA__11175__Y _05886_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06929_ net886 _01879_ _01868_ _01862_ vssd1 vssd1 vccd1 vccd1 _01880_ sky130_fd_sc_hd__o2bb2a_2
XANTENNA__11638__A2 net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout934_A net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout555_X net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09700__A1 _04618_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08503__A2 _03450_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09648_ _02996_ _03026_ _04427_ vssd1 vssd1 vccd1 vccd1 _04567_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_2_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_1816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_1851 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout722_X net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09579_ _03071_ _03102_ _04496_ _03581_ vssd1 vssd1 vccd1 vccd1 _04498_ sky130_fd_sc_hd__a31oi_1
XANTENNA__11191__X _05900_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11610_ net428 net566 _06162_ net299 net1475 vssd1 vssd1 vccd1 vccd1 _00437_ sky130_fd_sc_hd__a32o_1
XFILLER_0_38_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12063__A2 net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12590_ net1444 net997 net983 final_design.data_from_mem\[8\] vssd1 vssd1 vccd1 vccd1
+ _01283_ sky130_fd_sc_hd__a22o_1
XANTENNA__09464__B1 net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11271__B1 _05970_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11541_ net428 net566 _06126_ net303 net1687 vssd1 vssd1 vccd1 vccd1 _00404_ sky130_fd_sc_hd__a32o_1
XFILLER_0_9_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11472_ net205 net2252 net306 vssd1 vssd1 vccd1 vccd1 _00354_ sky130_fd_sc_hd__mux2_1
X_13211_ clknet_leaf_66_clk _00442_ net1063 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[199\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09767__A1 net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10423_ _03065_ _05190_ vssd1 vssd1 vccd1 vccd1 _05195_ sky130_fd_sc_hd__nor2_1
X_14191_ net1250 vssd1 vssd1 vccd1 vccd1 gpio_oeb[3] sky130_fd_sc_hd__buf_2
XFILLER_0_81_1415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10377__A2 net1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08660__B _03610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13142_ clknet_leaf_60_clk _00373_ net1140 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[130\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input63_A mem_adr_start[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10354_ net27 net1025 net1008 final_design.data_from_mem\[3\] vssd1 vssd1 vccd1 vccd1
+ _00107_ sky130_fd_sc_hd__a22o_1
X_13073_ clknet_leaf_34_clk _00304_ net1242 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[61\]
+ sky130_fd_sc_hd__dfrtp_1
X_10285_ net2549 _05139_ _05141_ net798 vssd1 vssd1 vccd1 vccd1 _00030_ sky130_fd_sc_hd__o211a_1
XANTENNA__11326__A1 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12523__B1 net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09772__A net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12024_ net804 _05841_ vssd1 vssd1 vccd1 vccd1 _06259_ sky130_fd_sc_hd__and2_1
XFILLER_0_79_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_1877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11877__A2 net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08742__A2 _01537_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08388__A net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06753__A1 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout590 net591 vssd1 vssd1 vccd1 vccd1 net590 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12836__CLK clknet_leaf_19_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13975_ clknet_leaf_6_clk _01206_ net1129 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[963\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkload9_A clknet_leaf_56_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12926_ clknet_leaf_49_clk _00164_ net1181 vssd1 vssd1 vccd1 vccd1 net149 sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_17_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12857_ clknet_leaf_17_clk _00095_ net1109 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.ready_data\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_48_1860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_44_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11808_ net2461 net414 net286 _06082_ vssd1 vssd1 vccd1 vccd1 _00561_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_44_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07075__A1_N net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11739_ net227 net2335 net417 vssd1 vssd1 vccd1 vccd1 _00502_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11801__A2 net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09207__B1 _04125_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09758__A1 net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13409_ clknet_leaf_48_clk _00640_ net1200 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[397\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11565__A1 net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06667__S1 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10605__B final_design.VGA_adr\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08950_ _03669_ _03752_ vssd1 vssd1 vccd1 vccd1 _03890_ sky130_fd_sc_hd__xnor2_1
XANTENNA__13611__CLK clknet_leaf_52_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12514__B1 net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11317__B2 net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07901_ final_design.cpu.reg_window\[983\] final_design.cpu.reg_window\[1015\] net849
+ vssd1 vssd1 vccd1 vccd1 _02852_ sky130_fd_sc_hd__mux2_1
X_08881_ _03800_ _03828_ vssd1 vssd1 vccd1 vccd1 _03829_ sky130_fd_sc_hd__nor2_1
XFILLER_0_47_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07832_ _02779_ _02780_ _02781_ _02782_ net685 net706 vssd1 vssd1 vccd1 vccd1 _02783_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__12312__S net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07092__S1 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13761__CLK clknet_leaf_47_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07763_ final_design.cpu.reg_window\[24\] final_design.cpu.reg_window\[56\] net862
+ vssd1 vssd1 vccd1 vccd1 _02714_ sky130_fd_sc_hd__mux2_1
X_09502_ net451 _04392_ _04419_ net727 vssd1 vssd1 vccd1 vccd1 _04421_ sky130_fd_sc_hd__a211o_2
X_06714_ final_design.cpu.reg_window\[216\] final_design.cpu.reg_window\[248\] net942
+ vssd1 vssd1 vccd1 vccd1 _01665_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07694_ final_design.cpu.reg_window\[283\] final_design.cpu.reg_window\[315\] net869
+ vssd1 vssd1 vccd1 vccd1 _02645_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07930__A net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09433_ net260 _03592_ _03033_ vssd1 vssd1 vccd1 vccd1 _04352_ sky130_fd_sc_hd__o21bai_2
X_06645_ net884 _01589_ _01595_ _01582_ _01583_ vssd1 vssd1 vccd1 vccd1 _01596_ sky130_fd_sc_hd__a32oi_4
XANTENNA_fanout250_A net251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout348_A net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14117__CLK clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09364_ _02702_ _04282_ _02672_ vssd1 vssd1 vccd1 vccd1 _04283_ sky130_fd_sc_hd__a21oi_1
X_06576_ _01523_ _01524_ _01525_ _01526_ net777 net794 vssd1 vssd1 vccd1 vccd1 _01527_
+ sky130_fd_sc_hd__mux4_1
X_08315_ final_design.cpu.reg_window\[456\] final_design.cpu.reg_window\[488\] net810
+ vssd1 vssd1 vccd1 vccd1 _03266_ sky130_fd_sc_hd__mux2_1
XANTENNA__09997__A1 _04124_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_2260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_20 final_design.reqhand.data_from_UART\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09295_ net462 _04208_ _04213_ vssd1 vssd1 vccd1 vccd1 _04214_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_60_2271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout515_A net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08246_ net538 _03194_ vssd1 vssd1 vccd1 vccd1 _03197_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_62_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13141__CLK clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08177_ _03122_ _03127_ net707 vssd1 vssd1 vccd1 vccd1 _03128_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout303_X net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10359__A2 net1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07128_ net752 _02072_ net746 vssd1 vssd1 vccd1 vccd1 _02079_ sky130_fd_sc_hd__o21a_1
XANTENNA__08421__A1 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout884_A net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_2042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07059_ final_design.cpu.reg_window\[13\] final_design.cpu.reg_window\[45\] net930
+ vssd1 vssd1 vccd1 vccd1 _02010_ sky130_fd_sc_hd__mux2_1
XANTENNA__13291__CLK clknet_leaf_38_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_2053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput160 net160 vssd1 vssd1 vccd1 vccd1 DAT_O[4] sky130_fd_sc_hd__buf_2
XANTENNA_fanout1212_X net1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_2064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput171 net171 vssd1 vssd1 vccd1 vccd1 WE_O sky130_fd_sc_hd__buf_2
XANTENNA__12505__B1 net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12859__CLK clknet_leaf_17_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10070_ wb_manage.curr_state\[0\] net801 _04988_ _01372_ wb_manage.curr_state\[1\]
+ vssd1 vssd1 vccd1 vccd1 _00004_ sky130_fd_sc_hd__a32o_1
XANTENNA__11859__A2 net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout672_X net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11627__A net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06735__B2 net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout937_X net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13760_ clknet_leaf_11_clk _00991_ net1087 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[748\]
+ sky130_fd_sc_hd__dfrtp_1
X_10972_ _05697_ _05698_ _05678_ vssd1 vssd1 vccd1 vccd1 _05699_ sky130_fd_sc_hd__o21ai_1
XANTENNA__08032__S0 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12711_ final_design.VGA_data_control.v_count\[3\] _06351_ vssd1 vssd1 vccd1 vccd1
+ _06352_ sky130_fd_sc_hd__or2_1
X_13691_ clknet_leaf_65_clk _00922_ net1070 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[679\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08583__S1 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11362__A net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12642_ _06308_ net1580 net978 vssd1 vssd1 vccd1 vccd1 _01323_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12573_ net1806 _06291_ _06286_ vssd1 vssd1 vccd1 vccd1 _01271_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11795__B2 net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11524_ net580 net196 _06116_ vssd1 vssd1 vccd1 vccd1 _06122_ sky130_fd_sc_hd__and3_1
XFILLER_0_81_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06897__S1 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14243_ net1297 vssd1 vssd1 vccd1 vccd1 gpio_out[21] sky130_fd_sc_hd__buf_2
XFILLER_0_0_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11455_ net225 net2458 net307 vssd1 vssd1 vccd1 vccd1 _00344_ sky130_fd_sc_hd__mux2_1
XANTENNA__13634__CLK clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11547__B2 net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09204__A3 _04117_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10406_ _03415_ _05181_ vssd1 vssd1 vccd1 vccd1 _05186_ sky130_fd_sc_hd__nor2_1
XFILLER_0_61_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14174_ clknet_leaf_21_clk _01348_ net1160 vssd1 vssd1 vccd1 vccd1 final_design.VGA_adr\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11386_ net643 _06071_ _05947_ _01538_ vssd1 vssd1 vccd1 vccd1 _06072_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__10425__B _05190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14181__Q final_design.VGA_adr\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13125_ clknet_leaf_49_clk _00356_ net1184 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[113\]
+ sky130_fd_sc_hd__dfrtp_1
X_10337_ net1494 net1009 net986 final_design.data_from_mem\[22\] vssd1 vssd1 vccd1
+ vccd1 _00094_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13056_ clknet_leaf_11_clk _00287_ net1086 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[44\]
+ sky130_fd_sc_hd__dfrtp_1
X_10268_ final_design.uart.BAUD_counter\[25\] _05129_ net797 vssd1 vssd1 vccd1 vccd1
+ _05131_ sky130_fd_sc_hd__o21ai_1
XANTENNA__13784__CLK clknet_leaf_65_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12007_ _06209_ net276 net400 net1990 vssd1 vssd1 vccd1 vccd1 _00738_ sky130_fd_sc_hd__a22o_1
XANTENNA__12132__S net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10199_ _05072_ _05081_ _05084_ _05087_ vssd1 vssd1 vccd1 vccd1 _05088_ sky130_fd_sc_hd__or4_1
XANTENNA__08271__S0 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13014__CLK clknet_leaf_60_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13958_ clknet_leaf_51_clk _01189_ net1174 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[946\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12909_ clknet_leaf_61_clk _00147_ net1140 vssd1 vssd1 vccd1 vccd1 net162 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_75_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13889_ clknet_leaf_47_clk _01120_ net1202 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[877\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_820 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06430_ net44 vssd1 vssd1 vccd1 vccd1 _01385_ sky130_fd_sc_hd__inv_2
XFILLER_0_75_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13164__CLK clknet_leaf_47_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08100_ _03047_ _03048_ _03049_ _03050_ net675 net697 vssd1 vssd1 vccd1 vccd1 _03051_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__11786__B2 _05952_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09080_ _02270_ _02434_ vssd1 vssd1 vccd1 vccd1 _04005_ sky130_fd_sc_hd__or2_1
XANTENNA__11250__A3 _05952_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08031_ final_design.cpu.reg_window\[915\] final_design.cpu.reg_window\[947\] net830
+ vssd1 vssd1 vccd1 vccd1 _02982_ sky130_fd_sc_hd__mux2_1
Xinput40 mem_adr_start[13] vssd1 vssd1 vccd1 vccd1 net40 sky130_fd_sc_hd__buf_1
XFILLER_0_82_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06662__B1 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07468__Y _02419_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12307__S net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput51 mem_adr_start[23] vssd1 vssd1 vccd1 vccd1 net51 sky130_fd_sc_hd__clkbuf_1
Xinput62 mem_adr_start[4] vssd1 vssd1 vccd1 vccd1 net62 sky130_fd_sc_hd__clkbuf_1
Xhold802 final_design.cpu.reg_window\[929\] vssd1 vssd1 vccd1 vccd1 net2144 sky130_fd_sc_hd__dlygate4sd3_1
Xinput73 memory_size[14] vssd1 vssd1 vccd1 vccd1 net73 sky130_fd_sc_hd__buf_1
XANTENNA__07197__A net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput84 memory_size[24] vssd1 vssd1 vccd1 vccd1 net84 sky130_fd_sc_hd__buf_1
Xhold813 final_design.cpu.reg_window\[866\] vssd1 vssd1 vccd1 vccd1 net2155 sky130_fd_sc_hd__dlygate4sd3_1
Xinput95 memory_size[5] vssd1 vssd1 vccd1 vccd1 net95 sky130_fd_sc_hd__buf_1
Xhold824 final_design.cpu.reg_window\[954\] vssd1 vssd1 vccd1 vccd1 net2166 sky130_fd_sc_hd__dlygate4sd3_1
Xhold835 final_design.cpu.reg_window\[286\] vssd1 vssd1 vccd1 vccd1 net2177 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_978 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkload35_A clknet_leaf_46_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold846 final_design.cpu.reg_window\[53\] vssd1 vssd1 vccd1 vccd1 net2188 sky130_fd_sc_hd__dlygate4sd3_1
Xhold857 final_design.cpu.reg_window\[392\] vssd1 vssd1 vccd1 vccd1 net2199 sky130_fd_sc_hd__dlygate4sd3_1
Xhold868 final_design.cpu.reg_window\[769\] vssd1 vssd1 vccd1 vccd1 net2210 sky130_fd_sc_hd__dlygate4sd3_1
X_09982_ _03327_ _04899_ _04900_ net447 vssd1 vssd1 vccd1 vccd1 _04901_ sky130_fd_sc_hd__a211o_1
Xhold879 final_design.cpu.reg_window\[415\] vssd1 vssd1 vccd1 vccd1 net2221 sky130_fd_sc_hd__dlygate4sd3_1
X_08933_ net625 _03874_ _03655_ vssd1 vssd1 vccd1 vccd1 _03875_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_58_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout298_A net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12042__S net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08864_ net2543 net1014 _03809_ _03813_ vssd1 vssd1 vccd1 vccd1 _00241_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout1005_A _05172_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11710__A1 net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07815_ net604 _02763_ _02739_ _01657_ vssd1 vssd1 vccd1 vccd1 _02766_ sky130_fd_sc_hd__o211a_1
XFILLER_0_58_1225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08795_ final_design.CPU_instr_adr\[16\] _01939_ vssd1 vssd1 vccd1 vccd1 _03746_
+ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout465_A net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07746_ _02691_ _02696_ net711 vssd1 vssd1 vccd1 vccd1 _02697_ sky130_fd_sc_hd__mux2_1
XANTENNA__12266__A2 net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13507__CLK clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07660__A _01507_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07677_ _02624_ _02625_ _02626_ _02627_ net684 net703 vssd1 vssd1 vccd1 vccd1 _02628_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_62_2311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout253_X net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout632_A net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_2322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06576__S0 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_2333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_2956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09416_ _04084_ _04202_ _04234_ _04073_ vssd1 vssd1 vccd1 vccd1 _04335_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_81_2967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06628_ final_design.cpu.reg_window\[219\] final_design.cpu.reg_window\[251\] net945
+ vssd1 vssd1 vccd1 vccd1 _01579_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_81_2978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12018__A2 net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1870 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10029__A1 net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08317__S1 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09347_ net527 net482 vssd1 vssd1 vccd1 vccd1 _04266_ sky130_fd_sc_hd__nor2_1
XANTENNA__11226__B1 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06559_ _01508_ _01509_ vssd1 vssd1 vccd1 vccd1 _01510_ sky130_fd_sc_hd__nand2b_1
XANTENNA_fanout420_X net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1162_X net1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13657__CLK clknet_leaf_52_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout518_X net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09278_ net92 _04196_ vssd1 vssd1 vccd1 vccd1 _04197_ sky130_fd_sc_hd__xor2_2
XFILLER_0_7_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1917 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06879__S1 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08229_ net710 _03173_ net724 vssd1 vssd1 vccd1 vccd1 _03180_ sky130_fd_sc_hd__o21a_1
XANTENNA__07850__C1 net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_2896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_2104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11529__A1 net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_2115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_2126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11240_ final_design.data_from_mem\[12\] _05914_ _05917_ vssd1 vssd1 vccd1 vccd1
+ _05943_ sky130_fd_sc_hd__a21o_1
XANTENNA__09874__X _04793_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_2137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_1696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11171_ _04825_ net653 _05843_ _05882_ vssd1 vssd1 vccd1 vccd1 _05883_ sky130_fd_sc_hd__a211oi_1
X_10122_ _01368_ _01370_ _05027_ _05030_ _04999_ vssd1 vssd1 vccd1 vccd1 final_design.vga.v_next_count\[7\]
+ sky130_fd_sc_hd__o311a_1
XANTENNA__13037__CLK clknet_leaf_44_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10053_ _04954_ _04956_ _04971_ net730 vssd1 vssd1 vccd1 vccd1 _04972_ sky130_fd_sc_hd__a22o_1
XANTENNA__07554__B _02504_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07056__S1 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06708__A1 final_design.data_from_mem\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input26_A DAT_I[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13812_ clknet_leaf_8_clk _01043_ net1153 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[800\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13187__CLK clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07570__A net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10955_ _05681_ _05682_ vssd1 vssd1 vccd1 vccd1 _05683_ sky130_fd_sc_hd__or2_1
X_13743_ clknet_leaf_43_clk _00974_ net1218 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[731\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12009__A2 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10886_ net960 _05615_ _05616_ net956 vssd1 vssd1 vccd1 vccd1 _05617_ sky130_fd_sc_hd__o2bb2a_1
X_13674_ clknet_leaf_60_clk _00905_ net1141 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[662\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12625_ final_design.VGA_data_control.ready_data\[0\] net1022 net977 final_design.data_from_mem\[0\]
+ vssd1 vssd1 vccd1 vccd1 _06300_ sky130_fd_sc_hd__a22o_1
XFILLER_0_39_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_14_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12556_ _06219_ net352 net324 net1855 vssd1 vssd1 vccd1 vccd1 _01260_ sky130_fd_sc_hd__a22o_1
XFILLER_0_81_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_16 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11507_ net2283 net224 net522 vssd1 vssd1 vccd1 vccd1 _00376_ sky130_fd_sc_hd__mux2_1
X_12487_ _06147_ net348 net331 net2233 vssd1 vssd1 vccd1 vccd1 _01193_ sky130_fd_sc_hd__a22o_1
XANTENNA__10436__A _03022_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold109 net152 vssd1 vssd1 vccd1 vccd1 net1451 sky130_fd_sc_hd__dlygate4sd3_1
X_14226_ net1280 vssd1 vssd1 vccd1 vccd1 gpio_out[4] sky130_fd_sc_hd__buf_2
X_11438_ net2131 net182 net312 vssd1 vssd1 vccd1 vccd1 _00335_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_1725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14157_ clknet_leaf_18_clk _01331_ net1112 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.data_to_VGA\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_46_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11369_ _01599_ _05947_ _06056_ net644 vssd1 vssd1 vccd1 vccd1 _06057_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_10_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08492__S0 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13108_ clknet_leaf_13_clk _00339_ net1088 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[96\]
+ sky130_fd_sc_hd__dfrtp_1
X_14088_ clknet_leaf_9_clk _01285_ net1152 vssd1 vssd1 vccd1 vccd1 final_design.reqhand.instruction\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10442__Y _05205_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13039_ clknet_leaf_42_clk _00270_ net1219 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_28_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12496__A2 net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09897__B1 net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1160 net1161 vssd1 vssd1 vccd1 vccd1 net1160 sky130_fd_sc_hd__clkbuf_4
Xfanout1171 net1176 vssd1 vssd1 vccd1 vccd1 net1171 sky130_fd_sc_hd__clkbuf_2
Xfanout1182 net1192 vssd1 vssd1 vccd1 vccd1 net1182 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_28_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1193 net1197 vssd1 vssd1 vccd1 vccd1 net1193 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_59_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07600_ _02547_ _02548_ _02549_ _02550_ net687 net694 vssd1 vssd1 vccd1 vccd1 _02551_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_72_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08580_ final_design.cpu.reg_window\[0\] final_design.cpu.reg_window\[32\] net814
+ vssd1 vssd1 vccd1 vccd1 _03531_ sky130_fd_sc_hd__mux2_1
XANTENNA__06795__S net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07531_ _02478_ _02479_ _02480_ _02481_ net776 net793 vssd1 vssd1 vccd1 vccd1 _02482_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_72_1745 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09744__S0 net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08547__S1 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1789 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07462_ final_design.cpu.reg_window\[704\] final_design.cpu.reg_window\[736\] net908
+ vssd1 vssd1 vccd1 vccd1 _02413_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_1188 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09201_ net594 _04112_ vssd1 vssd1 vccd1 vccd1 _04120_ sky130_fd_sc_hd__or2_1
X_06413_ final_design.VGA_data_control.v_count\[7\] vssd1 vssd1 vccd1 vccd1 _01368_
+ sky130_fd_sc_hd__inv_2
XANTENNA__11208__B1 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07393_ net752 _02337_ net746 vssd1 vssd1 vccd1 vccd1 _02344_ sky130_fd_sc_hd__o21a_1
XFILLER_0_56_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09132_ _02610_ _04050_ vssd1 vssd1 vccd1 vccd1 _04051_ sky130_fd_sc_hd__and2_1
XANTENNA__12420__A2 net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09200__A net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09063_ final_design.CPU_instr_adr\[8\] _03990_ net1037 vssd1 vssd1 vccd1 vccd1 _00219_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12037__S net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout213_A _05951_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09694__X _04613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08014_ _01908_ _02904_ _02930_ _02964_ vssd1 vssd1 vccd1 vccd1 _02965_ sky130_fd_sc_hd__o31a_1
Xhold610 final_design.cpu.reg_window\[399\] vssd1 vssd1 vccd1 vccd1 net1952 sky130_fd_sc_hd__dlygate4sd3_1
Xhold621 final_design.cpu.reg_window\[435\] vssd1 vssd1 vccd1 vccd1 net1963 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12184__A1 net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold632 final_design.cpu.reg_window\[579\] vssd1 vssd1 vccd1 vccd1 net1974 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold643 final_design.cpu.reg_window\[739\] vssd1 vssd1 vccd1 vccd1 net1985 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_2602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold654 final_design.cpu.reg_window\[332\] vssd1 vssd1 vccd1 vccd1 net1996 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_70_2613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07286__S1 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold665 final_design.cpu.reg_window\[88\] vssd1 vssd1 vccd1 vccd1 net2007 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1122_A net1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold676 final_design.cpu.reg_window\[367\] vssd1 vssd1 vccd1 vccd1 net2018 sky130_fd_sc_hd__dlygate4sd3_1
Xhold687 final_design.cpu.reg_window\[278\] vssd1 vssd1 vccd1 vccd1 net2029 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11931__B2 net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07655__A _01567_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10290__S0 net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold698 final_design.cpu.reg_window\[881\] vssd1 vssd1 vccd1 vccd1 net2040 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08250__S net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09965_ _04788_ _04828_ _04882_ _04883_ vssd1 vssd1 vccd1 vccd1 _04884_ sky130_fd_sc_hd__and4_1
XANTENNA_fanout582_A net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08916_ net257 _03859_ net1014 vssd1 vssd1 vccd1 vccd1 _03860_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12487__A2 net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09896_ net537 net535 net534 net533 net455 net461 vssd1 vssd1 vccd1 vccd1 _04815_
+ sky130_fd_sc_hd__mux4_2
XANTENNA_fanout1008_X net1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09352__A2 net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08847_ final_design.CPU_instr_adr\[25\] final_design.CPU_instr_adr\[24\] _03797_
+ vssd1 vssd1 vccd1 vccd1 _03798_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_68_2520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout370_X net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_2531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_2542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06797__S0 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout847_A net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08778_ _03725_ _03727_ _03695_ _03696_ vssd1 vssd1 vccd1 vccd1 _03729_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_64_2406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08486__A net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07729_ final_design.cpu.reg_window\[90\] final_design.cpu.reg_window\[122\] net865
+ vssd1 vssd1 vccd1 vccd1 _02680_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout635_X net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_1741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10740_ net41 _05476_ vssd1 vssd1 vccd1 vccd1 _05478_ sky130_fd_sc_hd__xor2_1
XFILLER_0_67_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08863__A1 _03655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10671_ _05410_ _05411_ vssd1 vssd1 vccd1 vccd1 _05412_ sky130_fd_sc_hd__xor2_1
XANTENNA_fanout802_X net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12410_ _06106_ net353 net341 net2097 vssd1 vssd1 vccd1 vccd1 _01120_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_11_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13390_ clknet_leaf_42_clk _00621_ net1223 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[378\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12411__A2 net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12341_ net2383 net360 net344 _05935_ vssd1 vssd1 vccd1 vccd1 _01053_ sky130_fd_sc_hd__a22o_1
XFILLER_0_63_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10422__B2 net246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12272_ net557 _06202_ net503 net368 net1864 vssd1 vssd1 vccd1 vccd1 _00987_ sky130_fd_sc_hd__a32o_1
X_14011_ clknet_leaf_66_clk _01242_ net1070 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[999\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_62_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11223_ net646 net218 vssd1 vssd1 vccd1 vccd1 _05929_ sky130_fd_sc_hd__and2_1
X_11154_ _05839_ _05866_ vssd1 vssd1 vccd1 vccd1 _05868_ sky130_fd_sc_hd__and2_4
XFILLER_0_43_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10105_ _05019_ vssd1 vssd1 vccd1 vccd1 _05020_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_8_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11085_ _05801_ _05806_ vssd1 vssd1 vccd1 vccd1 _05807_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_8_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07029__S1 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12478__A2 net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11518__C _06116_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10036_ net80 _04189_ vssd1 vssd1 vccd1 vccd1 _04955_ sky130_fd_sc_hd__xor2_2
XANTENNA_input29_X net29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11686__B1 net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13822__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09726__S0 net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11987_ _06189_ net293 net406 net2191 vssd1 vssd1 vccd1 vccd1 _00720_ sky130_fd_sc_hd__a22o_1
XFILLER_0_58_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13726_ clknet_leaf_11_clk _00957_ net1097 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[714\]
+ sky130_fd_sc_hd__dfrtp_1
X_10938_ net1003 _05665_ _05666_ net1033 net1345 vssd1 vssd1 vccd1 vccd1 _00196_ sky130_fd_sc_hd__a32o_1
XFILLER_0_14_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13972__CLK clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10869_ net48 _05599_ vssd1 vssd1 vccd1 vccd1 _05601_ sky130_fd_sc_hd__nor2_1
XFILLER_0_73_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13657_ clknet_leaf_52_clk _00888_ net1170 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[645\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12608_ net1424 net998 net984 final_design.data_from_mem\[26\] vssd1 vssd1 vccd1
+ vccd1 _01301_ sky130_fd_sc_hd__a22o_1
XFILLER_0_27_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08335__S net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12402__A2 net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06644__A net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13588_ clknet_leaf_10_clk _00819_ net1102 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[576\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11610__B1 net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10413__B2 net246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1224 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12539_ _06202_ net343 net322 net2254 vssd1 vssd1 vccd1 vccd1 _01243_ sky130_fd_sc_hd__a22o_1
XFILLER_0_30_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13202__CLK clknet_leaf_39_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14209_ net1267 vssd1 vssd1 vccd1 vccd1 gpio_oeb[21] sky130_fd_sc_hd__buf_2
XFILLER_0_2_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07475__A _02419_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08070__S net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11709__B net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13352__CLK clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout408 net409 vssd1 vssd1 vccd1 vccd1 net408 sky130_fd_sc_hd__buf_4
Xfanout419 _06226_ vssd1 vssd1 vccd1 vccd1 net419 sky130_fd_sc_hd__clkbuf_8
X_06962_ final_design.cpu.reg_window\[336\] final_design.cpu.reg_window\[368\] net927
+ vssd1 vssd1 vccd1 vccd1 _01913_ sky130_fd_sc_hd__mux2_1
X_09750_ _03198_ net446 _04222_ _04268_ _04668_ vssd1 vssd1 vccd1 vccd1 _04669_ sky130_fd_sc_hd__o221a_1
XANTENNA__12469__A2 net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09690__A net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08701_ _03645_ _03651_ vssd1 vssd1 vccd1 vccd1 _03652_ sky130_fd_sc_hd__nand2_2
XFILLER_0_39_1905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09681_ _03165_ _04505_ vssd1 vssd1 vccd1 vccd1 _04600_ sky130_fd_sc_hd__xnor2_1
X_06893_ final_design.cpu.reg_window\[723\] final_design.cpu.reg_window\[755\] net911
+ vssd1 vssd1 vccd1 vccd1 _01844_ sky130_fd_sc_hd__mux2_1
XANTENNA__06779__S0 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08632_ net543 _03104_ _03130_ _03134_ _03582_ vssd1 vssd1 vccd1 vccd1 _03583_ sky130_fd_sc_hd__o32a_1
XANTENNA__12320__S net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07414__S net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08563_ net876 _03506_ _03512_ _03499_ _03500_ vssd1 vssd1 vccd1 vccd1 _03514_ sky130_fd_sc_hd__a32o_1
XFILLER_0_77_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07514_ _01759_ _01789_ _02463_ _01757_ vssd1 vssd1 vccd1 vccd1 _02465_ sky130_fd_sc_hd__o31a_1
XFILLER_0_76_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11163__C net242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08494_ final_design.cpu.reg_window\[643\] final_design.cpu.reg_window\[675\] net826
+ vssd1 vssd1 vccd1 vccd1 _03445_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07445_ final_design.cpu.reg_window\[320\] final_design.cpu.reg_window\[352\] net909
+ vssd1 vssd1 vccd1 vccd1 _02396_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout330_A net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1072_A net1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout428_A net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11460__A net221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07376_ final_design.data_from_mem\[10\] net970 vssd1 vssd1 vccd1 vccd1 _02327_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_21_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_2800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09115_ _04034_ final_design.CPU_instr_adr\[0\] _03812_ vssd1 vssd1 vccd1 vccd1 _00209_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_76_2811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11601__B1 net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08073__A2 _03022_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10507__C net1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09046_ _03693_ _03695_ vssd1 vssd1 vccd1 vccd1 _03975_ sky130_fd_sc_hd__nor2_1
XANTENNA__14080__RESET_B net1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold440 final_design.cpu.reg_window\[753\] vssd1 vssd1 vccd1 vccd1 net1782 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold451 final_design.cpu.reg_window\[648\] vssd1 vssd1 vccd1 vccd1 net1793 sky130_fd_sc_hd__dlygate4sd3_1
Xhold462 final_design.cpu.reg_window\[517\] vssd1 vssd1 vccd1 vccd1 net1804 sky130_fd_sc_hd__dlygate4sd3_1
Xhold473 final_design.cpu.reg_window\[903\] vssd1 vssd1 vccd1 vccd1 net1815 sky130_fd_sc_hd__dlygate4sd3_1
Xhold484 final_design.cpu.reg_window\[534\] vssd1 vssd1 vccd1 vccd1 net1826 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11619__B net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold495 final_design.cpu.reg_window\[574\] vssd1 vssd1 vccd1 vccd1 net1837 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout964_A net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout585_X net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout920 net922 vssd1 vssd1 vccd1 vccd1 net920 sky130_fd_sc_hd__clkbuf_4
Xfanout931 net932 vssd1 vssd1 vccd1 vccd1 net931 sky130_fd_sc_hd__buf_4
XANTENNA__11380__A2 _06065_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout942 net945 vssd1 vssd1 vccd1 vccd1 net942 sky130_fd_sc_hd__clkbuf_4
X_09948_ _04755_ _04866_ net481 vssd1 vssd1 vccd1 vccd1 _04867_ sky130_fd_sc_hd__mux2_1
XANTENNA__13845__CLK clknet_leaf_57_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout953 _01420_ vssd1 vssd1 vccd1 vccd1 net953 sky130_fd_sc_hd__clkbuf_8
Xfanout964 net967 vssd1 vssd1 vccd1 vccd1 net964 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08646__A_N _01686_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout975 _06299_ vssd1 vssd1 vccd1 vccd1 net975 sky130_fd_sc_hd__clkbuf_2
Xfanout986 _05167_ vssd1 vssd1 vccd1 vccd1 net986 sky130_fd_sc_hd__buf_2
XANTENNA__11668__B1 net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout997 net999 vssd1 vssd1 vccd1 vccd1 net997 sky130_fd_sc_hd__clkbuf_4
X_09879_ net528 net456 _04061_ net465 vssd1 vssd1 vccd1 vccd1 _04798_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout752_X net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1140 final_design.cpu.reg_window\[620\] vssd1 vssd1 vccd1 vccd1 net2482 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1151 final_design.cpu.reg_window\[185\] vssd1 vssd1 vccd1 vccd1 net2493 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11635__A net206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11910_ net193 _06248_ _06249_ net274 net2266 vssd1 vssd1 vccd1 vccd1 _00650_ sky130_fd_sc_hd__a32o_1
Xhold1162 final_design.cpu.reg_window\[117\] vssd1 vssd1 vccd1 vccd1 net2504 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12230__S net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1173 final_design.cpu.reg_window\[956\] vssd1 vssd1 vccd1 vccd1 net2515 sky130_fd_sc_hd__dlygate4sd3_1
X_12890_ clknet_leaf_18_clk _00128_ net1112 vssd1 vssd1 vccd1 vccd1 final_design.data_from_mem\[24\]
+ sky130_fd_sc_hd__dfrtp_4
Xhold1184 final_design.cpu.reg_window\[829\] vssd1 vssd1 vccd1 vccd1 net2526 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1195 final_design.uart.bits_received\[3\] vssd1 vssd1 vccd1 vccd1 net2537 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13995__CLK clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11841_ net178 net1994 net266 vssd1 vssd1 vccd1 vccd1 _00593_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11772_ _05849_ net555 net241 vssd1 vssd1 vccd1 vccd1 _06229_ sky130_fd_sc_hd__and3_1
XANTENNA__12093__B1 net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10723_ _05458_ _05459_ _05461_ net1032 net1371 vssd1 vssd1 vccd1 vccd1 _00186_ sky130_fd_sc_hd__a32o_1
X_13511_ clknet_leaf_63_clk _00742_ net1122 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[499\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06735__Y _01686_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13225__CLK clknet_leaf_36_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input93_A memory_size[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10654_ net957 _05395_ _05394_ net960 vssd1 vssd1 vccd1 vccd1 _05396_ sky130_fd_sc_hd__a2bb2o_1
X_13442_ clknet_leaf_11_clk _00673_ net1097 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[430\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13373_ clknet_leaf_5_clk _00604_ net1081 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[361\]
+ sky130_fd_sc_hd__dfrtp_1
X_10585_ net728 _04903_ net247 net668 vssd1 vssd1 vccd1 vccd1 _05330_ sky130_fd_sc_hd__a31o_1
Xclkload18 clknet_leaf_18_clk vssd1 vssd1 vccd1 vccd1 clkload18/X sky130_fd_sc_hd__clkbuf_4
Xclkload29 clknet_leaf_51_clk vssd1 vssd1 vccd1 vccd1 clkload29/X sky130_fd_sc_hd__clkbuf_8
X_12324_ net1746 net185 net367 vssd1 vssd1 vccd1 vccd1 _01038_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_1408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09775__A net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13375__CLK clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11369__X _06057_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14245__1299 vssd1 vssd1 vccd1 vccd1 _14245__1299/HI net1299 sky130_fd_sc_hd__conb_1
X_12255_ net582 _06184_ net514 net375 net1515 vssd1 vssd1 vccd1 vccd1 _00971_ sky130_fd_sc_hd__a32o_1
XANTENNA__09494__B _04087_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1875 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11206_ net245 _05854_ vssd1 vssd1 vccd1 vccd1 _05913_ sky130_fd_sc_hd__nand2_1
X_12186_ net1605 net195 net381 vssd1 vssd1 vccd1 vccd1 _00905_ sky130_fd_sc_hd__mux2_1
X_11137_ final_design.CPU_instr_adr\[0\] net734 net662 _04032_ net654 vssd1 vssd1
+ vccd1 vccd1 _05852_ sky130_fd_sc_hd__a221o_1
XANTENNA__07670__S1 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11068_ net57 _05790_ vssd1 vssd1 vccd1 vccd1 _05791_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_34_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_3004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10019_ _03642_ net447 vssd1 vssd1 vccd1 vccd1 _04938_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_82_3015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12140__S net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_3026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10331__B1 net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_3037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_3048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14000__CLK clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1873 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12084__B1 net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11831__A0 net197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13709_ clknet_leaf_48_clk _00940_ net1200 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[697\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_28_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1879 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_28_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09669__B net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06645__Y _01596_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14150__CLK clknet_leaf_15_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07230_ final_design.cpu.reg_window\[904\] final_design.cpu.reg_window\[936\] net897
+ vssd1 vssd1 vccd1 vccd1 _02181_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13718__CLK clknet_leaf_59_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07161_ _02108_ _02109_ _02110_ _02111_ net765 net786 vssd1 vssd1 vccd1 vccd1 _02112_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_48_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07092_ _02039_ _02040_ _02041_ _02042_ net765 net786 vssd1 vssd1 vccd1 vccd1 _02043_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_48_1076 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_1833 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12315__S net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13868__CLK clknet_leaf_46_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11347__C1 net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11898__A0 net209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_1877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08212__C1 net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout205 net206 vssd1 vssd1 vccd1 vccd1 net205 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_10_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout216 net217 vssd1 vssd1 vccd1 vccd1 net216 sky130_fd_sc_hd__buf_2
Xfanout227 _05883_ vssd1 vssd1 vccd1 vccd1 net227 sky130_fd_sc_hd__buf_2
X_09802_ _03358_ _04720_ vssd1 vssd1 vccd1 vccd1 _04721_ sky130_fd_sc_hd__xnor2_1
Xfanout238 _05904_ vssd1 vssd1 vccd1 vccd1 net238 sky130_fd_sc_hd__clkbuf_2
Xfanout249 _04986_ vssd1 vssd1 vccd1 vccd1 net249 sky130_fd_sc_hd__buf_4
X_07994_ final_design.cpu.reg_window\[208\] final_design.cpu.reg_window\[240\] net846
+ vssd1 vssd1 vccd1 vccd1 _02945_ sky130_fd_sc_hd__mux2_1
XANTENNA__12892__CLK clknet_leaf_15_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06945_ net756 _01889_ net747 vssd1 vssd1 vccd1 vccd1 _01896_ sky130_fd_sc_hd__o21ai_1
X_09733_ _03071_ _04496_ vssd1 vssd1 vccd1 vccd1 _04652_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout280_A net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12311__A1 net207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout378_A net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12050__S net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06876_ final_design.cpu.reg_window\[275\] final_design.cpu.reg_window\[307\] net911
+ vssd1 vssd1 vccd1 vccd1 _01827_ sky130_fd_sc_hd__mux2_1
X_09664_ _04108_ _04309_ _04117_ vssd1 vssd1 vccd1 vccd1 _04583_ sky130_fd_sc_hd__o21a_1
XANTENNA__10322__B1 net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10873__A1 _05508_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08615_ _02211_ _03297_ _03322_ vssd1 vssd1 vccd1 vccd1 _03566_ sky130_fd_sc_hd__and3b_1
X_09595_ _02704_ _04049_ net321 vssd1 vssd1 vccd1 vccd1 _04514_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout545_A _01908_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13248__CLK clknet_leaf_11_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12075__B1 net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08546_ final_design.cpu.reg_window\[129\] final_design.cpu.reg_window\[161\] net836
+ vssd1 vssd1 vccd1 vccd1 _03497_ sky130_fd_sc_hd__mux2_1
XANTENNA__08764__A final_design.CPU_instr_adr\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11822__A0 net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1733 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08477_ final_design.cpu.reg_window\[259\] final_design.cpu.reg_window\[291\] net831
+ vssd1 vssd1 vccd1 vccd1 _03428_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout333_X net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout712_A net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12090__A3 net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1777 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07428_ final_design.cpu.reg_window\[961\] final_design.cpu.reg_window\[993\] net913
+ vssd1 vssd1 vccd1 vccd1 _02379_ sky130_fd_sc_hd__mux2_1
XANTENNA__13398__CLK clknet_leaf_59_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12378__A1 net207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07359_ _02306_ _02307_ _02308_ _02309_ net767 net787 vssd1 vssd1 vccd1 vccd1 _02310_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout500_X net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10389__B1 net1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10928__A2 net1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10370_ net12 net1026 net1008 final_design.data_from_mem\[19\] vssd1 vssd1 vccd1
+ vccd1 _00123_ sky130_fd_sc_hd__a22o_1
XFILLER_0_61_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09029_ _02445_ _03959_ vssd1 vssd1 vccd1 vccd1 _03960_ sky130_fd_sc_hd__xor2_1
XANTENNA__12800__31_A clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12040_ net1863 net210 net398 vssd1 vssd1 vccd1 vccd1 _00768_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_1452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold270 final_design.cpu.reg_window\[203\] vssd1 vssd1 vccd1 vccd1 net1612 sky130_fd_sc_hd__dlygate4sd3_1
Xhold281 final_design.cpu.reg_window\[59\] vssd1 vssd1 vccd1 vccd1 net1623 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout967_X net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold292 final_design.cpu.reg_window\[239\] vssd1 vssd1 vccd1 vccd1 net1634 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11353__A2 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout750 net751 vssd1 vssd1 vccd1 vccd1 net750 sky130_fd_sc_hd__buf_2
XANTENNA__14023__CLK clknet_leaf_63_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout761 net762 vssd1 vssd1 vccd1 vccd1 net761 sky130_fd_sc_hd__buf_2
Xfanout772 net779 vssd1 vssd1 vccd1 vccd1 net772 sky130_fd_sc_hd__buf_4
X_13991_ clknet_leaf_63_clk _01222_ net1123 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[979\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout783 net784 vssd1 vssd1 vccd1 vccd1 net783 sky130_fd_sc_hd__buf_4
XANTENNA__12302__A1 net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout794 net795 vssd1 vssd1 vccd1 vccd1 net794 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_38_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09703__C1 _04341_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07562__B net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12942_ clknet_leaf_23_clk _00180_ net1165 vssd1 vssd1 vccd1 vccd1 net130 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_77_1272 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06459__A net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07054__S net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10864__A1 net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10864__B2 net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12873_ clknet_leaf_14_clk _00111_ net1111 vssd1 vssd1 vccd1 vccd1 final_design.data_from_mem\[7\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__14173__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11824_ net209 net2036 net266 vssd1 vssd1 vccd1 vccd1 _00576_ sky130_fd_sc_hd__mux2_1
XANTENNA__12066__B1 net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09157__S1 net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11813__A0 net242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11755_ net200 net2379 net417 vssd1 vssd1 vccd1 vccd1 _00518_ sky130_fd_sc_hd__mux2_1
XANTENNA__09482__A1 net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10706_ net72 net1043 vssd1 vssd1 vccd1 vccd1 _05445_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_42_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11686_ net558 net420 _06201_ net294 net1741 vssd1 vssd1 vccd1 vccd1 _00474_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_42_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13425_ clknet_leaf_35_clk _00656_ net1241 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[413\]
+ sky130_fd_sc_hd__dfrtp_1
X_10637_ net958 _05377_ _05379_ net957 vssd1 vssd1 vccd1 vccd1 _05380_ sky130_fd_sc_hd__o22a_1
XFILLER_0_23_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10568_ _05288_ _05313_ vssd1 vssd1 vccd1 vccd1 _05314_ sky130_fd_sc_hd__nand2_1
X_13356_ clknet_leaf_45_clk _00587_ net1216 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[344\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12307_ net1765 net217 net364 vssd1 vssd1 vccd1 vccd1 _01021_ sky130_fd_sc_hd__mux2_1
XANTENNA__12135__S net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10499_ net1002 _05247_ _05248_ net1029 net123 vssd1 vssd1 vccd1 vccd1 _00175_ sky130_fd_sc_hd__a32o_1
X_13287_ clknet_leaf_63_clk _00518_ net1121 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[275\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10444__A _02894_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12238_ net557 _06168_ net503 net372 net1541 vssd1 vssd1 vccd1 vccd1 _00955_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_36_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11344__A2 net235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12169_ net1955 net225 net382 vssd1 vssd1 vccd1 vccd1 _00888_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_32_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07643__S1 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06771__A2 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput5 DAT_I[12] vssd1 vssd1 vccd1 vccd1 net5 sky130_fd_sc_hd__clkbuf_1
X_06730_ final_design.cpu.reg_window\[536\] final_design.cpu.reg_window\[568\] net935
+ vssd1 vssd1 vccd1 vccd1 _01681_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06661_ net761 _01611_ vssd1 vssd1 vccd1 vccd1 _01612_ sky130_fd_sc_hd__or2_1
XFILLER_0_36_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08400_ _03345_ _03350_ net709 vssd1 vssd1 vccd1 vccd1 _03351_ sky130_fd_sc_hd__mux2_1
X_09380_ net550 net549 net548 net546 net458 net469 vssd1 vssd1 vccd1 vccd1 _04299_
+ sky130_fd_sc_hd__mux4_1
X_06592_ final_design.cpu.reg_window\[156\] final_design.cpu.reg_window\[188\] net940
+ vssd1 vssd1 vccd1 vccd1 _01543_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08584__A net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13540__CLK clknet_leaf_54_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08331_ final_design.cpu.reg_window\[648\] final_design.cpu.reg_window\[680\] net808
+ vssd1 vssd1 vccd1 vccd1 _03282_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11804__B1 net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08276__A2 _03224_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12072__A3 net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1717 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1917 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08262_ final_design.cpu.reg_window\[842\] final_design.cpu.reg_window\[874\] net828
+ vssd1 vssd1 vccd1 vccd1 _03213_ sky130_fd_sc_hd__mux2_1
XANTENNA__08681__C1 _02542_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07213_ _02160_ _02161_ _02162_ _02163_ net766 net785 vssd1 vssd1 vccd1 vccd1 _02164_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_55_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08193_ final_design.cpu.reg_window\[206\] final_design.cpu.reg_window\[238\] net812
+ vssd1 vssd1 vccd1 vccd1 _03144_ sky130_fd_sc_hd__mux2_1
XANTENNA__13690__CLK clknet_leaf_63_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07144_ final_design.reqhand.instruction\[7\] final_design.data_from_mem\[7\] net971
+ vssd1 vssd1 vccd1 vccd1 _02095_ sky130_fd_sc_hd__mux2_2
XFILLER_0_82_1917 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06832__A net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11583__A2 net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07075_ net885 _02025_ _02014_ _02008_ vssd1 vssd1 vccd1 vccd1 _02026_ sky130_fd_sc_hd__o2bb2a_2
XANTENNA__12045__S net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1035_A net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07139__S net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14046__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10073__B net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout495_A _03419_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1202_A net1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07977_ _02922_ _02927_ net714 vssd1 vssd1 vccd1 vccd1 _02928_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout283_X net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout662_A net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_21_clk_X clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12780__11_A clknet_leaf_28_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13070__CLK clknet_leaf_45_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09716_ net727 _04626_ _04630_ _04633_ _04185_ vssd1 vssd1 vccd1 vccd1 _04635_ sky130_fd_sc_hd__o311ai_1
X_06928_ _01873_ _01878_ net756 vssd1 vssd1 vccd1 vccd1 _01879_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_1543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07398__S0 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout450_X net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09647_ _04046_ _04553_ _04554_ _04564_ vssd1 vssd1 vccd1 vccd1 _04566_ sky130_fd_sc_hd__a31o_1
X_06859_ final_design.cpu.reg_window\[660\] final_design.cpu.reg_window\[692\] net947
+ vssd1 vssd1 vccd1 vccd1 _01810_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1192_X net1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout548_X net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout927_A net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14244__1298 vssd1 vssd1 vccd1 vccd1 _14244__1298/HI net1298 sky130_fd_sc_hd__conb_1
XANTENNA_clkbuf_leaf_36_clk_X clknet_leaf_36_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09578_ _03071_ _04496_ _03580_ vssd1 vssd1 vccd1 vccd1 _04497_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_17_1863 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07602__S net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12599__B2 final_design.data_from_mem\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08529_ _03474_ _03479_ net710 vssd1 vssd1 vccd1 vccd1 _03480_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout715_X net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10529__A net1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12063__A3 net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11271__A1 net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11540_ net228 net635 vssd1 vssd1 vccd1 vccd1 _06126_ sky130_fd_sc_hd__and2_1
XFILLER_0_68_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11471_ net206 net638 vssd1 vssd1 vccd1 vccd1 _06107_ sky130_fd_sc_hd__and2_1
XFILLER_0_0_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10422_ net1611 net1030 _05194_ net246 vssd1 vssd1 vccd1 vccd1 _00152_ sky130_fd_sc_hd__a22o_1
X_13210_ clknet_leaf_1_clk _00441_ net1082 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[198\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12220__B1 net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14190_ net1249 vssd1 vssd1 vccd1 vccd1 gpio_oeb[2] sky130_fd_sc_hd__buf_2
X_13141_ clknet_leaf_6_clk _00372_ net1134 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[129\]
+ sky130_fd_sc_hd__dfrtp_1
X_10353_ net24 net1025 _05170_ final_design.data_from_mem\[2\] vssd1 vssd1 vccd1 vccd1
+ _00106_ sky130_fd_sc_hd__a22o_1
XFILLER_0_63_1861 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13072_ clknet_leaf_33_clk _00303_ net1238 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[60\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input56_A mem_adr_start[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10284_ final_design.uart.BAUD_counter\[31\] _05139_ vssd1 vssd1 vccd1 vccd1 _05141_
+ sky130_fd_sc_hd__nand2_1
X_12023_ _06225_ net289 net403 net2296 vssd1 vssd1 vccd1 vccd1 _00754_ sky130_fd_sc_hd__a22o_1
XANTENNA__13413__CLK clknet_leaf_48_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06888__S net913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1889 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08669__A _01999_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09117__X _04036_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout580 net587 vssd1 vssd1 vccd1 vccd1 net580 sky130_fd_sc_hd__clkbuf_2
Xfanout591 _05844_ vssd1 vssd1 vccd1 vccd1 net591 sky130_fd_sc_hd__buf_2
XANTENNA__12287__B1 net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13974_ clknet_leaf_59_clk _01205_ net1138 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[962\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09152__B1 net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14179__Q final_design.VGA_adr\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13563__CLK clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12925_ clknet_leaf_61_clk _00163_ net1137 vssd1 vssd1 vccd1 vccd1 net148 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12856_ clknet_leaf_17_clk _00094_ net1109 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.ready_data\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_1821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_48_1850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11542__B net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11807_ net2481 net414 net292 _06075_ vssd1 vssd1 vccd1 vccd1 _00560_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_44_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11738_ net242 net1910 net417 vssd1 vssd1 vccd1 vccd1 _00501_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09207__A1 _02545_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11669_ net805 _02358_ net803 vssd1 vssd1 vccd1 vccd1 _06192_ sky130_fd_sc_hd__and3_2
XFILLER_0_71_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07748__A _01630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13408_ clknet_leaf_10_clk _00639_ net1101 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[396\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12211__B1 net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14069__CLK clknet_leaf_15_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07313__S0 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11565__A2 net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13339_ clknet_leaf_64_clk _00570_ net1074 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[327\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_38_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1901 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11317__A2 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13093__CLK clknet_leaf_49_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07900_ net714 _02844_ net723 vssd1 vssd1 vccd1 vccd1 _02851_ sky130_fd_sc_hd__o21a_1
XANTENNA__09682__B net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08880_ final_design.CPU_instr_adr\[27\] _03799_ final_design.CPU_instr_adr\[28\]
+ vssd1 vssd1 vccd1 vccd1 _03828_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11868__A3 net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07831_ final_design.cpu.reg_window\[405\] final_design.cpu.reg_window\[437\] net858
+ vssd1 vssd1 vccd1 vccd1 _02782_ sky130_fd_sc_hd__mux2_1
XANTENNA__11717__B net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13906__CLK clknet_leaf_44_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12278__B1 net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07762_ final_design.cpu.reg_window\[88\] final_design.cpu.reg_window\[120\] net862
+ vssd1 vssd1 vccd1 vccd1 _02713_ sky130_fd_sc_hd__mux2_1
X_09501_ net451 _04392_ _04419_ vssd1 vssd1 vccd1 vccd1 _04420_ sky130_fd_sc_hd__a21o_1
X_06713_ final_design.cpu.reg_window\[24\] final_design.cpu.reg_window\[56\] net942
+ vssd1 vssd1 vccd1 vccd1 _01664_ sky130_fd_sc_hd__mux2_1
X_07693_ final_design.cpu.reg_window\[347\] final_design.cpu.reg_window\[379\] net869
+ vssd1 vssd1 vccd1 vccd1 _02644_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09694__A1 net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12293__A3 net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11733__A net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12930__CLK clknet_leaf_47_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06644_ net761 _01594_ vssd1 vssd1 vccd1 vccd1 _01595_ sky130_fd_sc_hd__or2_1
X_09432_ _02935_ net260 _03589_ vssd1 vssd1 vccd1 vccd1 _04351_ sky130_fd_sc_hd__or3_1
XANTENNA__11452__B net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09363_ _02735_ _02768_ _04281_ _02766_ _02705_ vssd1 vssd1 vccd1 vccd1 _04282_ sky130_fd_sc_hd__a311o_1
X_06575_ final_design.cpu.reg_window\[925\] final_design.cpu.reg_window\[957\] net949
+ vssd1 vssd1 vccd1 vccd1 _01526_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout243_A net244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1861 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08314_ final_design.cpu.reg_window\[264\] final_design.cpu.reg_window\[296\] net820
+ vssd1 vssd1 vccd1 vccd1 _03265_ sky130_fd_sc_hd__mux2_1
X_09294_ net467 _04203_ _04207_ vssd1 vssd1 vccd1 vccd1 _04213_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_60_2250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_10 _06285_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_2261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_21 net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_2272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08245_ net611 _03192_ _03193_ net538 vssd1 vssd1 vccd1 vccd1 _03196_ sky130_fd_sc_hd__a211oi_1
XANTENNA__12564__A net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout410_A net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06833__Y _01784_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1152_A net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout508_A net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08176_ _03123_ _03124_ _03125_ _03126_ net674 net691 vssd1 vssd1 vccd1 vccd1 _03127_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__12202__B1 net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08406__C1 _02239_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09749__A2 net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08253__S net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07127_ net760 _02077_ vssd1 vssd1 vccd1 vccd1 _02078_ sky130_fd_sc_hd__or2_1
XFILLER_0_63_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_1867 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_63_clk_A clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13436__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10764__B1 net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1038_X net1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_2190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07058_ final_design.cpu.reg_window\[77\] final_design.cpu.reg_window\[109\] net930
+ vssd1 vssd1 vccd1 vccd1 _02009_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_54_2043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput150 net150 vssd1 vssd1 vccd1 vccd1 DAT_O[24] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_54_2054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput161 net161 vssd1 vssd1 vccd1 vccd1 DAT_O[5] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_54_2065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout877_A net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput172 net172 vssd1 vssd1 vccd1 vccd1 gpio_out[0] sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_73_2699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout498_X net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13586__CLK clknet_leaf_38_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11627__B net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout665_X net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12269__B1 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_6_Left_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10971_ net85 net1045 vssd1 vssd1 vccd1 vccd1 _05698_ sky130_fd_sc_hd__nor2_1
XANTENNA__09685__A1 net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12739__A _05058_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08032__S1 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12284__A3 net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12710_ _06349_ _06350_ vssd1 vssd1 vccd1 vccd1 _06351_ sky130_fd_sc_hd__nor2_2
XANTENNA__07696__A0 final_design.cpu.reg_window\[411\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13690_ clknet_leaf_63_clk _00921_ net1121 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[678\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06737__A net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12641_ final_design.VGA_data_control.ready_data\[8\] net1019 net974 final_design.data_from_mem\[8\]
+ vssd1 vssd1 vccd1 vccd1 _06308_ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_16_clk_A clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_567 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12572_ final_design.uart.receiving final_design.uart.working_data\[6\] vssd1 vssd1
+ vccd1 vccd1 _06291_ sky130_fd_sc_hd__and2_1
XFILLER_0_80_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07543__S0 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11795__A2 net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11523_ net1847 net197 net523 vssd1 vssd1 vccd1 vccd1 _00391_ sky130_fd_sc_hd__mux2_1
Xwire211 _05958_ vssd1 vssd1 vccd1 vccd1 net211 sky130_fd_sc_hd__buf_2
XFILLER_0_68_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08671__B _01598_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14242_ net1296 vssd1 vssd1 vccd1 vccd1 gpio_out[20] sky130_fd_sc_hd__buf_2
X_11454_ net225 net639 vssd1 vssd1 vccd1 vccd1 _06100_ sky130_fd_sc_hd__and2_1
XFILLER_0_46_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11547__A2 net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10405_ net1454 net1027 _05185_ net246 vssd1 vssd1 vccd1 vccd1 _00144_ sky130_fd_sc_hd__a22o_1
X_14173_ clknet_leaf_21_clk _01347_ net1160 vssd1 vssd1 vccd1 vccd1 final_design.VGA_adr\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_11385_ final_design.data_from_mem\[29\] net236 net234 vssd1 vssd1 vccd1 vccd1 _06071_
+ sky130_fd_sc_hd__a21o_1
XANTENNA__09070__C1 net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13124_ clknet_leaf_53_clk _00355_ net1187 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[112\]
+ sky130_fd_sc_hd__dfrtp_1
X_10336_ net1507 net1009 net986 final_design.data_from_mem\[21\] vssd1 vssd1 vccd1
+ vccd1 _00093_ sky130_fd_sc_hd__a22o_1
XANTENNA__13929__CLK clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11377__X _06064_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10267_ _05129_ _05130_ vssd1 vssd1 vccd1 vccd1 _00022_ sky130_fd_sc_hd__nor2_1
X_13055_ clknet_leaf_8_clk _00286_ net1154 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[43\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10722__A net1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12006_ _06208_ net278 net400 net2250 vssd1 vssd1 vccd1 vccd1 _00737_ sky130_fd_sc_hd__a22o_1
X_10198_ _05076_ _05085_ _05086_ vssd1 vssd1 vccd1 vccd1 _05087_ sky130_fd_sc_hd__or3_1
XFILLER_0_20_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08271__S1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12953__CLK clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09007__B net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09125__B1 net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13957_ clknet_leaf_50_clk _01188_ net1181 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[945\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12275__A3 net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12908_ clknet_leaf_61_clk _00146_ net1140 vssd1 vssd1 vccd1 vccd1 net161 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_48_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13888_ clknet_leaf_10_clk _01119_ net1101 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[876\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13309__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12839_ clknet_leaf_19_clk _00077_ net1156 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.ready_data\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09428__A1 _04334_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11235__A1 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08862__A net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11786__A2 net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13459__CLK clknet_leaf_40_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08030_ final_design.cpu.reg_window\[979\] final_design.cpu.reg_window\[1011\] net830
+ vssd1 vssd1 vccd1 vccd1 _02981_ sky130_fd_sc_hd__mux2_1
XANTENNA__06662__A1 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput30 DAT_I[6] vssd1 vssd1 vccd1 vccd1 net30 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput41 mem_adr_start[14] vssd1 vssd1 vccd1 vccd1 net41 sky130_fd_sc_hd__buf_1
XFILLER_0_71_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput52 mem_adr_start[24] vssd1 vssd1 vccd1 vccd1 net52 sky130_fd_sc_hd__clkbuf_1
Xinput63 mem_adr_start[5] vssd1 vssd1 vccd1 vccd1 net63 sky130_fd_sc_hd__buf_1
Xhold803 final_design.cpu.reg_window\[347\] vssd1 vssd1 vccd1 vccd1 net2145 sky130_fd_sc_hd__dlygate4sd3_1
Xinput74 memory_size[15] vssd1 vssd1 vccd1 vccd1 net74 sky130_fd_sc_hd__buf_1
Xhold814 final_design.cpu.reg_window\[253\] vssd1 vssd1 vccd1 vccd1 net2156 sky130_fd_sc_hd__dlygate4sd3_1
Xinput85 memory_size[25] vssd1 vssd1 vccd1 vccd1 net85 sky130_fd_sc_hd__buf_1
XANTENNA__09061__C1 _03655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold825 final_design.cpu.reg_window\[540\] vssd1 vssd1 vccd1 vccd1 net2167 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08403__A2 _03352_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput96 memory_size[6] vssd1 vssd1 vccd1 vccd1 net96 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__10746__B1 _04990_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold836 final_design.cpu.reg_window\[68\] vssd1 vssd1 vccd1 vccd1 net2178 sky130_fd_sc_hd__dlygate4sd3_1
Xhold847 final_design.cpu.reg_window\[618\] vssd1 vssd1 vccd1 vccd1 net2189 sky130_fd_sc_hd__dlygate4sd3_1
Xhold858 final_design.cpu.reg_window\[819\] vssd1 vssd1 vccd1 vccd1 net2200 sky130_fd_sc_hd__dlygate4sd3_1
X_09981_ _03327_ _03356_ _04706_ vssd1 vssd1 vccd1 vccd1 _04900_ sky130_fd_sc_hd__and3b_1
Xhold869 final_design.cpu.reg_window\[861\] vssd1 vssd1 vccd1 vccd1 net2211 sky130_fd_sc_hd__dlygate4sd3_1
X_14243__1297 vssd1 vssd1 vccd1 vccd1 _14243__1297/HI net1297 sky130_fd_sc_hd__conb_1
XANTENNA_clkload28_A clknet_leaf_49_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08932_ _03862_ _03873_ vssd1 vssd1 vccd1 vccd1 _03874_ sky130_fd_sc_hd__or2_1
XANTENNA__12323__S net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12499__B1 net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07417__S net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09903__A2 _04559_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1805 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08863_ _03655_ _03811_ net1038 vssd1 vssd1 vccd1 vccd1 _03813_ sky130_fd_sc_hd__o21a_1
XANTENNA__11171__B1 _05843_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout193_A _06031_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11710__A2 net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07814_ net604 _02763_ _02739_ vssd1 vssd1 vccd1 vccd1 _02765_ sky130_fd_sc_hd__o21a_1
XFILLER_0_77_1849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08794_ _03679_ _03740_ _03743_ _03744_ vssd1 vssd1 vccd1 vccd1 _03745_ sky130_fd_sc_hd__or4_1
XFILLER_0_58_1237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07745_ _02692_ _02693_ _02694_ _02695_ net686 net694 vssd1 vssd1 vccd1 vccd1 _02696_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_79_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout360_A net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout458_A net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_66_2470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07676_ final_design.cpu.reg_window\[926\] final_design.cpu.reg_window\[958\] net855
+ vssd1 vssd1 vccd1 vccd1 _02627_ sky130_fd_sc_hd__mux2_1
XANTENNA__06557__A _01453_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_2312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07773__S0 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07152__S net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06576__S1 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_2323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_2957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09415_ _04107_ _04241_ _04116_ vssd1 vssd1 vccd1 vccd1 _04334_ sky130_fd_sc_hd__a21oi_2
XTAP_TAPCELL_ROW_62_2334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_2968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06627_ final_design.cpu.reg_window\[27\] final_design.cpu.reg_window\[59\] net941
+ vssd1 vssd1 vccd1 vccd1 _01578_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_2979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout246_X net246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1882 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout625_A _02506_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11226__A1 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12423__B1 net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09346_ net473 _04075_ _04086_ vssd1 vssd1 vccd1 vccd1 _04265_ sky130_fd_sc_hd__or3_1
XANTENNA__09868__A net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06558_ _01453_ _01507_ vssd1 vssd1 vccd1 vccd1 _01509_ sky130_fd_sc_hd__or2_1
XFILLER_0_14_1877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11777__A2 net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09277_ net89 net91 _04195_ vssd1 vssd1 vccd1 vccd1 _04196_ sky130_fd_sc_hd__or3_1
X_06489_ final_design.cpu.reg_window\[862\] final_design.cpu.reg_window\[894\] net936
+ vssd1 vssd1 vccd1 vccd1 _01440_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout413_X net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08228_ net718 _03178_ vssd1 vssd1 vccd1 vccd1 _03179_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_79_2886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_2105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_2897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_2116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_2127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08159_ _03106_ _03107_ _03108_ _03109_ net676 net696 vssd1 vssd1 vccd1 vccd1 _03110_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__10737__B1 net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11170_ net651 _05879_ _05881_ vssd1 vssd1 vccd1 vccd1 _05882_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout782_X net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10121_ final_design.VGA_data_control.v_count\[6\] _05026_ final_design.VGA_data_control.v_count\[7\]
+ vssd1 vssd1 vccd1 vccd1 _05030_ sky130_fd_sc_hd__a21o_1
XANTENNA__12976__CLK clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07327__S net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10052_ _04659_ _04676_ vssd1 vssd1 vccd1 vccd1 _04971_ sky130_fd_sc_hd__nor2_1
XFILLER_0_41_1274 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11162__B1 net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13811_ clknet_leaf_40_clk _01042_ net1211 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[799\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07851__A net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input19_A DAT_I[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12257__A3 net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11373__A net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13742_ clknet_leaf_43_clk _00973_ net1218 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[730\]
+ sky130_fd_sc_hd__dfrtp_1
X_10954_ _05676_ _05680_ vssd1 vssd1 vccd1 vccd1 _05682_ sky130_fd_sc_hd__and2b_1
XFILLER_0_39_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13673_ clknet_leaf_37_clk _00904_ net1228 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[661\]
+ sky130_fd_sc_hd__dfrtp_1
X_10885_ final_design.CPU_instr_adr\[21\] _03887_ net1059 vssd1 vssd1 vccd1 vccd1
+ _05616_ sky130_fd_sc_hd__mux2_1
XANTENNA__11217__A1 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13601__CLK clknet_leaf_47_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12624_ _05165_ net1022 vssd1 vssd1 vccd1 vccd1 _06299_ sky130_fd_sc_hd__nor2_2
XFILLER_0_54_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09778__A net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12414__B1 net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_14_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12555_ _06218_ net355 net324 net2063 vssd1 vssd1 vccd1 vccd1 _01259_ sky130_fd_sc_hd__a22o_1
X_11506_ net1619 net239 net521 vssd1 vssd1 vccd1 vccd1 _00375_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_28 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12486_ _06146_ net354 net332 net2086 vssd1 vssd1 vccd1 vccd1 _01192_ sky130_fd_sc_hd__a22o_1
XANTENNA__10436__B net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13751__CLK clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14225_ final_design.cpu.Error vssd1 vssd1 vccd1 vccd1 net175 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_80_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11437_ net1701 net185 net312 vssd1 vssd1 vccd1 vccd1 _00334_ sky130_fd_sc_hd__mux2_1
XANTENNA__09594__B1 net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14156_ clknet_leaf_18_clk _01330_ net1113 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.data_to_VGA\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11368_ final_design.data_from_mem\[27\] net236 net234 vssd1 vssd1 vccd1 vccd1 _06056_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_22_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08492__S1 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11548__A net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11940__A2 net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13107_ clknet_leaf_36_clk _00338_ net1210 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[95\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14107__CLK clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10319_ net1526 net1011 net988 final_design.data_from_mem\[4\] vssd1 vssd1 vccd1
+ vccd1 _00076_ sky130_fd_sc_hd__a22o_1
XANTENNA__12143__S net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10452__A _02698_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14087_ clknet_leaf_8_clk _01284_ net1152 vssd1 vssd1 vccd1 vccd1 final_design.reqhand.instruction\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_11299_ _04451_ net652 net590 _05995_ vssd1 vssd1 vccd1 vccd1 _05996_ sky130_fd_sc_hd__o211a_2
X_13038_ clknet_leaf_45_clk _00269_ net1213 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09897__A1 net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1150 net1167 vssd1 vssd1 vccd1 vccd1 net1150 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_28_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1161 net1162 vssd1 vssd1 vccd1 vccd1 net1161 sky130_fd_sc_hd__clkbuf_4
Xfanout1172 net1175 vssd1 vssd1 vccd1 vccd1 net1172 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06929__X _01880_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1183 net1192 vssd1 vssd1 vccd1 vccd1 net1183 sky130_fd_sc_hd__clkbuf_2
Xfanout1194 net1197 vssd1 vssd1 vccd1 vccd1 net1194 sky130_fd_sc_hd__clkbuf_4
XANTENNA__13131__CLK clknet_leaf_38_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06648__Y _01599_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07530_ final_design.cpu.reg_window\[415\] final_design.cpu.reg_window\[447\] net939
+ vssd1 vssd1 vccd1 vccd1 _02481_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09744__S1 net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07461_ _02408_ _02409_ _02410_ _02411_ net768 net788 vssd1 vssd1 vccd1 vccd1 _02412_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_9_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13281__CLK clknet_leaf_48_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09200_ net482 _04116_ vssd1 vssd1 vccd1 vccd1 _04119_ sky130_fd_sc_hd__nand2_2
X_06412_ net1018 vssd1 vssd1 vccd1 vccd1 _01367_ sky130_fd_sc_hd__inv_2
XANTENNA__11208__A1 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07392_ net760 _02342_ vssd1 vssd1 vccd1 vccd1 _02343_ sky130_fd_sc_hd__or2_1
XANTENNA__12405__B1 net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12849__CLK clknet_leaf_17_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09131_ _02706_ _02771_ _03594_ _03603_ vssd1 vssd1 vccd1 vccd1 _04050_ sky130_fd_sc_hd__a31o_1
XANTENNA__12318__S net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10967__B1 net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12420__A3 net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09062_ net254 _03987_ _03989_ vssd1 vssd1 vccd1 vccd1 _03990_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09200__B _04116_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08013_ _02932_ _02933_ _02963_ vssd1 vssd1 vccd1 vccd1 _02964_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_8_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold600 final_design.cpu.reg_window\[850\] vssd1 vssd1 vccd1 vccd1 net1942 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout206_A _05972_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold611 final_design.cpu.reg_window\[606\] vssd1 vssd1 vccd1 vccd1 net1953 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold622 final_design.cpu.reg_window\[674\] vssd1 vssd1 vccd1 vccd1 net1964 sky130_fd_sc_hd__dlygate4sd3_1
Xhold633 final_design.cpu.reg_window\[802\] vssd1 vssd1 vccd1 vccd1 net1975 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07936__A net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold644 final_design.cpu.reg_window\[456\] vssd1 vssd1 vccd1 vccd1 net1986 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_70_2603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold655 final_design.cpu.reg_window\[393\] vssd1 vssd1 vccd1 vccd1 net1997 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold666 final_design.cpu.reg_window\[489\] vssd1 vssd1 vccd1 vccd1 net2008 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11931__A2 net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold677 final_design.cpu.reg_window\[283\] vssd1 vssd1 vccd1 vccd1 net2019 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11458__A net244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold688 final_design.cpu.reg_window\[654\] vssd1 vssd1 vccd1 vccd1 net2030 sky130_fd_sc_hd__dlygate4sd3_1
X_09964_ _04848_ _04849_ _04881_ vssd1 vssd1 vccd1 vccd1 _04883_ sky130_fd_sc_hd__and3_1
Xhold699 final_design.cpu.reg_window\[327\] vssd1 vssd1 vccd1 vccd1 net2041 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12053__S net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10290__S1 net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1115_A net1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08915_ final_design.CPU_instr_adr\[24\] _03797_ vssd1 vssd1 vccd1 vccd1 _03859_
+ sky130_fd_sc_hd__xnor2_1
XANTENNA__11144__A0 net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09895_ _04794_ _04796_ net460 vssd1 vssd1 vccd1 vccd1 _04814_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_1613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11892__S net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout575_A net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout196_X net196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08846_ final_design.CPU_instr_adr\[23\] _03796_ vssd1 vssd1 vccd1 vccd1 _03797_
+ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_68_2521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_2532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07671__A net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_2543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06797__S1 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08777_ _03725_ _03727_ _03696_ vssd1 vssd1 vccd1 vccd1 _03728_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout742_A net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_2407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12239__A3 net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06571__B1 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout363_X net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13624__CLK clknet_leaf_65_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07728_ _02675_ _02676_ _02677_ _02678_ net686 net704 vssd1 vssd1 vccd1 vccd1 _02679_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__11998__A2 net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07659_ _02573_ _02575_ _02605_ _02607_ vssd1 vssd1 vccd1 vccd1 _02610_ sky130_fd_sc_hd__o22a_1
XFILLER_0_36_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout628_X net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09598__A _04097_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10670_ _05389_ _05393_ _05391_ vssd1 vssd1 vccd1 vccd1 _05411_ sky130_fd_sc_hd__o21a_1
XFILLER_0_36_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13774__CLK clknet_leaf_43_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09329_ net450 _04199_ _04245_ _04247_ vssd1 vssd1 vccd1 vccd1 _04248_ sky130_fd_sc_hd__a22o_1
XFILLER_0_63_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12411__A3 net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08171__S0 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10422__A2 net1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12340_ net2373 net360 net342 _05929_ vssd1 vssd1 vccd1 vccd1 _01052_ sky130_fd_sc_hd__a22o_1
XFILLER_0_35_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout997_X net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12271_ net562 _06201_ net502 net368 net1982 vssd1 vssd1 vccd1 vccd1 _00986_ sky130_fd_sc_hd__a32o_1
XFILLER_0_47_1461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14010_ clknet_leaf_63_clk _01241_ net1121 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[998\]
+ sky130_fd_sc_hd__dfrtp_1
X_11222_ net588 _05926_ _05927_ vssd1 vssd1 vccd1 vccd1 _05928_ sky130_fd_sc_hd__and3_1
XANTENNA__11383__B1 _01491_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11153_ net673 _02358_ _05838_ vssd1 vssd1 vccd1 vccd1 _05867_ sky130_fd_sc_hd__or3_1
X_10104_ final_design.VGA_data_control.v_count\[0\] final_design.VGA_data_control.v_count\[1\]
+ _05017_ vssd1 vssd1 vccd1 vccd1 _05019_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_8_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13154__CLK clknet_leaf_11_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11084_ _05804_ _05805_ vssd1 vssd1 vccd1 vccd1 _05806_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_8_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10035_ net727 _04950_ _04952_ vssd1 vssd1 vccd1 vccd1 _04954_ sky130_fd_sc_hd__or3_4
XFILLER_0_76_1123 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06468__Y _01419_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09726__S1 net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11986_ _06188_ net288 net406 net2067 vssd1 vssd1 vccd1 vccd1 _00719_ sky130_fd_sc_hd__a22o_1
XFILLER_0_59_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11989__A2 net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09500__B1 _04417_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13725_ clknet_leaf_2_clk _00956_ net1065 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[713\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10937_ _05643_ _05647_ _05664_ vssd1 vssd1 vccd1 vccd1 _05666_ sky130_fd_sc_hd__o21ai_1
XPHY_EDGE_ROW_9_Left_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14242__1296 vssd1 vssd1 vccd1 vccd1 _14242__1296/HI net1296 sky130_fd_sc_hd__conb_1
XFILLER_0_67_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13656_ clknet_leaf_65_clk _00887_ net1073 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[644\]
+ sky130_fd_sc_hd__dfrtp_1
X_10868_ net48 _05599_ vssd1 vssd1 vccd1 vccd1 _05600_ sky130_fd_sc_hd__and2_1
XFILLER_0_6_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12607_ net1458 net998 net984 final_design.data_from_mem\[25\] vssd1 vssd1 vccd1
+ vccd1 _01300_ sky130_fd_sc_hd__a22o_1
XANTENNA__11550__B net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09301__A net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12138__S net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13587_ clknet_leaf_40_clk _00818_ net1207 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[575\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10799_ _05532_ _05533_ vssd1 vssd1 vccd1 vccd1 _05534_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_26_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06617__A1 final_design.data_from_mem\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11610__A1 net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12538_ _06201_ net342 net322 net2273 vssd1 vssd1 vccd1 vccd1 _01242_ sky130_fd_sc_hd__a22o_1
XANTENNA__10166__B _05058_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1236 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12469_ _06253_ net498 net330 net2000 vssd1 vssd1 vccd1 vccd1 _01175_ sky130_fd_sc_hd__a22o_1
XFILLER_0_1_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09567__A0 net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14208_ net1266 vssd1 vssd1 vccd1 vccd1 gpio_oeb[20] sky130_fd_sc_hd__buf_2
XANTENNA__07756__A _01690_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11374__B1 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14139_ clknet_leaf_20_clk final_design.vga.h_next_count\[8\] net1115 vssd1 vssd1
+ vccd1 vccd1 final_design.VGA_data_control.h_count\[8\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout409 net411 vssd1 vssd1 vccd1 vccd1 net409 sky130_fd_sc_hd__buf_4
XFILLER_0_61_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09971__A net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07593__A2 _02540_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06961_ _01908_ _01910_ vssd1 vssd1 vccd1 vccd1 _01912_ sky130_fd_sc_hd__or2_1
XANTENNA__11126__B1 net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08700_ _03629_ _03650_ vssd1 vssd1 vccd1 vccd1 _03651_ sky130_fd_sc_hd__nor2_1
XANTENNA__13647__CLK clknet_leaf_44_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09680_ _04577_ _04598_ vssd1 vssd1 vccd1 vccd1 _04599_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10910__A net1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06892_ net751 _01842_ vssd1 vssd1 vccd1 vccd1 _01843_ sky130_fd_sc_hd__nor2_1
XFILLER_0_39_1917 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06779__S1 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07976__S0 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08631_ net599 _03160_ _03135_ _01996_ vssd1 vssd1 vccd1 vccd1 _03582_ sky130_fd_sc_hd__o211ai_2
XANTENNA__11284__Y _05982_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11725__B net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07750__C1 _01626_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08562_ net876 _03506_ _03512_ _03499_ _03500_ vssd1 vssd1 vccd1 vccd1 _03513_ sky130_fd_sc_hd__a32oi_4
XANTENNA__07728__S0 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13797__CLK clknet_leaf_52_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07513_ _01759_ _01789_ _02463_ vssd1 vssd1 vccd1 vccd1 _02464_ sky130_fd_sc_hd__or3_1
X_08493_ final_design.cpu.reg_window\[707\] final_design.cpu.reg_window\[739\] net826
+ vssd1 vssd1 vccd1 vccd1 _03444_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07444_ _02390_ _02394_ vssd1 vssd1 vccd1 vccd1 _02395_ sky130_fd_sc_hd__nand2_1
XFILLER_0_71_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10437__A1_N net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11460__B net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_21_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13027__CLK clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07375_ net882 _02318_ _02324_ _02311_ _02312_ vssd1 vssd1 vccd1 vccd1 _02326_ sky130_fd_sc_hd__a32o_2
XANTENNA__12048__S net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout323_A _06285_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1065_A net1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09114_ net619 _04032_ _04033_ _02426_ vssd1 vssd1 vccd1 vccd1 _04034_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_76_2801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_2812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11887__S net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09045_ final_design.CPU_instr_adr\[10\] _03974_ net1037 vssd1 vssd1 vccd1 vccd1
+ _00221_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1232_A net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout209_X net209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13177__CLK clknet_leaf_59_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold430 final_design.cpu.reg_window\[166\] vssd1 vssd1 vccd1 vccd1 net1772 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06570__A net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold441 final_design.cpu.reg_window\[247\] vssd1 vssd1 vccd1 vccd1 net1783 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11365__B1 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold452 final_design.cpu.reg_window\[457\] vssd1 vssd1 vccd1 vccd1 net1794 sky130_fd_sc_hd__dlygate4sd3_1
Xhold463 final_design.cpu.reg_window\[89\] vssd1 vssd1 vccd1 vccd1 net1805 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11188__A net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold474 final_design.cpu.reg_window\[346\] vssd1 vssd1 vccd1 vccd1 net1816 sky130_fd_sc_hd__dlygate4sd3_1
Xhold485 final_design.cpu.reg_window\[453\] vssd1 vssd1 vccd1 vccd1 net1827 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11089__A2_N net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1118_X net1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold496 final_design.cpu.reg_window\[74\] vssd1 vssd1 vccd1 vccd1 net1838 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout910 net953 vssd1 vssd1 vccd1 vccd1 net910 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_5_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout921 net922 vssd1 vssd1 vccd1 vccd1 net921 sky130_fd_sc_hd__clkbuf_4
Xfanout932 net953 vssd1 vssd1 vccd1 vccd1 net932 sky130_fd_sc_hd__buf_2
X_09947_ _04710_ _04865_ net471 vssd1 vssd1 vccd1 vccd1 _04866_ sky130_fd_sc_hd__mux2_1
Xfanout943 net944 vssd1 vssd1 vccd1 vccd1 net943 sky130_fd_sc_hd__clkbuf_4
Xfanout954 _05039_ vssd1 vssd1 vccd1 vccd1 net954 sky130_fd_sc_hd__buf_2
XANTENNA_fanout578_X net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout965 net967 vssd1 vssd1 vccd1 vccd1 net965 sky130_fd_sc_hd__clkbuf_2
Xfanout976 _06299_ vssd1 vssd1 vccd1 vccd1 net976 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11668__A1 net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout987 _05167_ vssd1 vssd1 vccd1 vccd1 net987 sky130_fd_sc_hd__clkbuf_2
X_09878_ net529 net456 _04063_ net460 vssd1 vssd1 vccd1 vccd1 _04797_ sky130_fd_sc_hd__a211o_1
Xfanout998 net999 vssd1 vssd1 vccd1 vccd1 net998 sky130_fd_sc_hd__clkbuf_4
Xhold1130 final_design.cpu.reg_window\[893\] vssd1 vssd1 vccd1 vccd1 net2472 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1141 final_design.cpu.reg_window\[921\] vssd1 vssd1 vccd1 vccd1 net2483 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11635__B net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1152 final_design.cpu.reg_window\[416\] vssd1 vssd1 vccd1 vccd1 net2494 sky130_fd_sc_hd__dlygate4sd3_1
X_08829_ final_design.CPU_instr_adr\[31\] _02504_ vssd1 vssd1 vccd1 vccd1 _03780_
+ sky130_fd_sc_hd__xnor2_1
Xhold1163 final_design.cpu.reg_window\[704\] vssd1 vssd1 vccd1 vccd1 net2505 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_77_1487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout745_X net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1174 final_design.cpu.reg_window\[313\] vssd1 vssd1 vccd1 vccd1 net2516 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10340__B2 final_design.data_from_mem\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1185 final_design.cpu.reg_window\[377\] vssd1 vssd1 vccd1 vccd1 net2527 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1196 final_design.CPU_instr_adr\[6\] vssd1 vssd1 vccd1 vccd1 net2538 sky130_fd_sc_hd__dlygate4sd3_1
X_11840_ net181 net2316 net266 vssd1 vssd1 vccd1 vccd1 _00592_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12093__A1 net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11771_ net2510 net413 net282 _05865_ vssd1 vssd1 vccd1 vccd1 _00532_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout912_X net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12747__A final_design.VGA_adr\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13510_ clknet_leaf_51_clk _00741_ net1169 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[498\]
+ sky130_fd_sc_hd__dfrtp_1
X_10722_ net1005 _05460_ vssd1 vssd1 vccd1 vccd1 _05461_ sky130_fd_sc_hd__nor2_1
XFILLER_0_3_1414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13441_ clknet_leaf_48_clk _00672_ net1200 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[429\]
+ sky130_fd_sc_hd__dfrtp_1
X_10653_ final_design.CPU_instr_adr\[10\] _03968_ net1058 vssd1 vssd1 vccd1 vccd1
+ _05395_ sky130_fd_sc_hd__mux2_1
XANTENNA_input86_A memory_size[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13372_ clknet_leaf_4_clk _00603_ net1083 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[360\]
+ sky130_fd_sc_hd__dfrtp_1
X_10584_ _05309_ _05327_ _05325_ vssd1 vssd1 vccd1 vccd1 _05329_ sky130_fd_sc_hd__a21oi_2
XANTENNA__08960__A net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload19 clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 clkload19/X sky130_fd_sc_hd__clkbuf_8
XANTENNA__12984__RESET_B net1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12323_ net2057 net186 net367 vssd1 vssd1 vccd1 vccd1 _01037_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_40_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09775__B _04693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07576__A net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12254_ net574 _06183_ net509 net375 net1785 vssd1 vssd1 vccd1 vccd1 _00970_ sky130_fd_sc_hd__a32o_1
XFILLER_0_62_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11205_ net245 _05854_ vssd1 vssd1 vccd1 vccd1 _05912_ sky130_fd_sc_hd__and2_1
XFILLER_0_27_1887 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12185_ _06122_ net501 _06270_ net2229 vssd1 vssd1 vccd1 vccd1 _00904_ sky130_fd_sc_hd__a22o_1
XFILLER_0_43_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11136_ net671 _05848_ _05850_ vssd1 vssd1 vccd1 vccd1 _05851_ sky130_fd_sc_hd__or3_4
XANTENNA__11385__X _06071_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09316__A3 _02325_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11067_ net966 _05789_ _05787_ _05778_ vssd1 vssd1 vccd1 vccd1 _05790_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_34_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_3005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10018_ _03612_ _03635_ _04053_ _04935_ vssd1 vssd1 vccd1 vccd1 _04937_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_82_3016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_3027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10331__B2 final_design.data_from_mem\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_3038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_3049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12608__B1 net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06630__S0 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_1825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_1885 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11969_ _06171_ net281 net405 net1821 vssd1 vssd1 vccd1 vccd1 _00702_ sky130_fd_sc_hd__a22o_1
XANTENNA__08827__A2 _01538_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13708_ clknet_leaf_45_clk _00939_ net1215 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[696\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_28_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07250__S net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13639_ clknet_leaf_62_clk _00870_ net1119 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[627\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_32_1582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11044__C1 net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07160_ final_design.cpu.reg_window\[138\] final_design.cpu.reg_window\[170\] net896
+ vssd1 vssd1 vccd1 vccd1 _02111_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11595__B1 net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07091_ final_design.cpu.reg_window\[140\] final_design.cpu.reg_window\[172\] net895
+ vssd1 vssd1 vccd1 vccd1 _02042_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_1801 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1845 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07015__B2 net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1889 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout206 _05972_ vssd1 vssd1 vccd1 vccd1 net206 sky130_fd_sc_hd__clkbuf_2
X_09801_ _03391_ _04718_ _03564_ vssd1 vssd1 vccd1 vccd1 _04720_ sky130_fd_sc_hd__a21o_1
Xfanout217 _05934_ vssd1 vssd1 vccd1 vccd1 net217 sky130_fd_sc_hd__buf_2
Xfanout228 _05864_ vssd1 vssd1 vccd1 vccd1 net228 sky130_fd_sc_hd__buf_2
Xfanout239 net240 vssd1 vssd1 vccd1 vccd1 net239 sky130_fd_sc_hd__buf_2
XANTENNA_clkload10_A clknet_leaf_57_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07993_ final_design.cpu.reg_window\[16\] final_design.cpu.reg_window\[48\] net846
+ vssd1 vssd1 vccd1 vccd1 _02944_ sky130_fd_sc_hd__mux2_1
X_09732_ net318 _04399_ _04647_ _04341_ _04650_ vssd1 vssd1 vccd1 vccd1 _04651_ sky130_fd_sc_hd__o221a_1
X_06944_ net763 _01894_ vssd1 vssd1 vccd1 vccd1 _01895_ sky130_fd_sc_hd__nor2_1
XFILLER_0_78_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09206__A _04124_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09663_ net494 _04581_ _04231_ vssd1 vssd1 vccd1 vccd1 _04582_ sky130_fd_sc_hd__a21o_1
X_06875_ final_design.cpu.reg_window\[339\] final_design.cpu.reg_window\[371\] net911
+ vssd1 vssd1 vccd1 vccd1 _01826_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout273_A net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06549__B net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08614_ net532 _03354_ vssd1 vssd1 vccd1 vccd1 _03565_ sky130_fd_sc_hd__nor2_1
X_09594_ _04282_ _04512_ net449 vssd1 vssd1 vccd1 vccd1 _04513_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_82_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_1903 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12075__A1 net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08545_ final_design.cpu.reg_window\[193\] final_design.cpu.reg_window\[225\] net836
+ vssd1 vssd1 vccd1 vccd1 _03496_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout440_A _04094_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1182_A net1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_59_Left_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11471__A net206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout538_A _02091_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08476_ final_design.cpu.reg_window\[323\] final_design.cpu.reg_window\[355\] net831
+ vssd1 vssd1 vccd1 vccd1 _03427_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08256__S net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1745 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_1611 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07427_ final_design.cpu.reg_window\[769\] final_design.cpu.reg_window\[801\] net914
+ vssd1 vssd1 vccd1 vccd1 _02378_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout705_A net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1789 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout326_X net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08126__S0 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1068_X net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07358_ final_design.cpu.reg_window\[131\] final_design.cpu.reg_window\[163\] net901
+ vssd1 vssd1 vccd1 vccd1 _02309_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10389__A1 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07289_ net741 _01628_ net666 vssd1 vssd1 vccd1 vccd1 _02240_ sky130_fd_sc_hd__mux2_2
XANTENNA_fanout1235_X net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11410__S net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09087__S net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13812__CLK clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09028_ _02100_ _02101_ vssd1 vssd1 vccd1 vccd1 _03959_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_68_Left_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11338__B1 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold260 final_design.VGA_data_control.data_to_VGA\[20\] vssd1 vssd1 vccd1 vccd1 net1602
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold271 final_design.cpu.reg_window\[58\] vssd1 vssd1 vccd1 vccd1 net1613 sky130_fd_sc_hd__dlygate4sd3_1
Xhold282 final_design.cpu.reg_window\[578\] vssd1 vssd1 vccd1 vccd1 net1624 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12550__A2 net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09951__B1 net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold293 final_design.cpu.reg_window\[906\] vssd1 vssd1 vccd1 vccd1 net1635 sky130_fd_sc_hd__dlygate4sd3_1
X_14241__1295 vssd1 vssd1 vccd1 vccd1 _14241__1295/HI net1295 sky130_fd_sc_hd__conb_1
XANTENNA_fanout862_X net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13962__CLK clknet_leaf_60_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout751 net752 vssd1 vssd1 vccd1 vccd1 net751 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_1773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout762 net763 vssd1 vssd1 vccd1 vccd1 net762 sky130_fd_sc_hd__clkbuf_4
X_13990_ clknet_leaf_51_clk _01221_ net1172 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[978\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout773 net779 vssd1 vssd1 vccd1 vccd1 net773 sky130_fd_sc_hd__buf_4
Xfanout784 _01419_ vssd1 vssd1 vccd1 vccd1 net784 sky130_fd_sc_hd__clkbuf_8
Xfanout795 _01418_ vssd1 vssd1 vccd1 vccd1 net795 sky130_fd_sc_hd__buf_4
X_12941_ clknet_leaf_22_clk _00179_ net1165 vssd1 vssd1 vccd1 vccd1 net129 sky130_fd_sc_hd__dfrtp_1
XANTENNA__10959__A1_N net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07562__C net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06459__B net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12872_ clknet_leaf_25_clk _00110_ net1157 vssd1 vssd1 vccd1 vccd1 final_design.data_from_mem\[6\]
+ sky130_fd_sc_hd__dfrtp_4
XPHY_EDGE_ROW_77_Left_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13183__RESET_B net1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12066__A1 net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11823_ net213 net1996 net264 vssd1 vssd1 vccd1 vccd1 _00575_ sky130_fd_sc_hd__mux2_1
XANTENNA__11381__A net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09122__Y _04041_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11754_ net201 net1853 net417 vssd1 vssd1 vccd1 vccd1 _00517_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07070__S net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09482__A2 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13342__CLK clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10705_ _04632_ net253 vssd1 vssd1 vccd1 vccd1 _05444_ sky130_fd_sc_hd__nor2_1
X_11685_ net243 net626 vssd1 vssd1 vccd1 vccd1 _06201_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_42_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13424_ clknet_leaf_37_clk _00655_ net1232 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[412\]
+ sky130_fd_sc_hd__dfrtp_1
X_10636_ final_design.CPU_instr_adr\[9\] _03981_ net1058 vssd1 vssd1 vccd1 vccd1 _05379_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08690__A _02419_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11577__B1 net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13355_ clknet_leaf_38_clk _00586_ net1189 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[343\]
+ sky130_fd_sc_hd__dfrtp_1
X_10567_ _05311_ _05312_ vssd1 vssd1 vccd1 vccd1 _05313_ sky130_fd_sc_hd__nand2_1
XFILLER_0_12_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13492__CLK clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08993__A1 net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12306_ net1880 net219 net364 vssd1 vssd1 vccd1 vccd1 _01020_ sky130_fd_sc_hd__mux2_1
X_13286_ clknet_leaf_51_clk _00517_ net1170 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[274\]
+ sky130_fd_sc_hd__dfrtp_1
X_10498_ _05233_ _05246_ vssd1 vssd1 vccd1 vccd1 _05248_ sky130_fd_sc_hd__nand2_1
XANTENNA__10444__B net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11329__B1 _06021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12237_ net558 _06167_ net502 net372 net1417 vssd1 vssd1 vccd1 vccd1 _00954_ sky130_fd_sc_hd__a32o_1
XFILLER_0_23_1515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12541__A2 net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12168_ net1753 net240 net380 vssd1 vssd1 vccd1 vccd1 _00887_ sky130_fd_sc_hd__mux2_1
X_11119_ _05064_ _05834_ vssd1 vssd1 vccd1 vccd1 _05836_ sky130_fd_sc_hd__or2_1
XANTENNA__10460__A _02635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12151__S net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12099_ net1705 net240 net388 vssd1 vssd1 vccd1 vccd1 _00823_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07245__S net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput6 DAT_I[13] vssd1 vssd1 vccd1 vccd1 net6 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11843__X _06238_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06660_ _01607_ _01608_ _01609_ _01610_ net775 net783 vssd1 vssd1 vccd1 vccd1 _01611_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__07720__A2 _02668_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06591_ final_design.cpu.reg_window\[220\] final_design.cpu.reg_window\[252\] net938
+ vssd1 vssd1 vccd1 vccd1 _01542_ sky130_fd_sc_hd__mux2_1
XANTENNA__08584__B _03534_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08356__S0 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08330_ final_design.cpu.reg_window\[712\] final_design.cpu.reg_window\[744\] net808
+ vssd1 vssd1 vccd1 vccd1 _03281_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11804__B2 _06053_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08261_ net716 _03211_ net722 vssd1 vssd1 vccd1 vccd1 _03212_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_69_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13835__CLK clknet_leaf_52_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07212_ final_design.cpu.reg_window\[392\] final_design.cpu.reg_window\[424\] net899
+ vssd1 vssd1 vccd1 vccd1 _02163_ sky130_fd_sc_hd__mux2_1
X_08192_ final_design.cpu.reg_window\[14\] final_design.cpu.reg_window\[46\] net812
+ vssd1 vssd1 vccd1 vccd1 _03143_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07143_ _01463_ net740 vssd1 vssd1 vccd1 vccd1 _02094_ sky130_fd_sc_hd__nand2_4
XANTENNA__12326__S net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09630__C1 net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07074_ _02019_ _02024_ net762 vssd1 vssd1 vccd1 vccd1 _02025_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_1620 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13985__CLK clknet_leaf_47_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10791__B2 net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08599__X _03550_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10073__C net251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1028_A net1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12532__A2 net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11740__A0 net240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout390_A net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13215__CLK clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07976_ _02923_ _02924_ _02925_ _02926_ net683 net693 vssd1 vssd1 vccd1 vccd1 _02927_
+ sky130_fd_sc_hd__mux4_1
X_09715_ _04185_ _04633_ vssd1 vssd1 vccd1 vccd1 _04634_ sky130_fd_sc_hd__nand2_1
X_06927_ _01874_ _01875_ _01876_ _01877_ net773 net784 vssd1 vssd1 vccd1 vccd1 _01878_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_74_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout655_A _05142_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout276_X net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07398__S1 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09646_ net485 _04559_ _04560_ _04224_ _04113_ vssd1 vssd1 vccd1 vccd1 _04565_ sky130_fd_sc_hd__a221o_1
X_06858_ final_design.cpu.reg_window\[724\] final_design.cpu.reg_window\[756\] net947
+ vssd1 vssd1 vccd1 vccd1 _01809_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_2_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13365__CLK clknet_leaf_55_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12048__A1 net196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09577_ _03231_ _04495_ _03572_ vssd1 vssd1 vccd1 vccd1 _04496_ sky130_fd_sc_hd__a21bo_1
XANTENNA_fanout822_A net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06789_ final_design.cpu.reg_window\[726\] final_design.cpu.reg_window\[758\] net920
+ vssd1 vssd1 vccd1 vccd1 _01740_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout443_X net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10059__B1 _04632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08528_ _03475_ _03476_ _03477_ _03478_ net679 net692 vssd1 vssd1 vccd1 vccd1 _03479_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_17_1875 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08459_ final_design.cpu.reg_window\[644\] final_design.cpu.reg_window\[676\] net819
+ vssd1 vssd1 vccd1 vccd1 _03410_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_14_Right_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11470_ net208 net2429 net306 vssd1 vssd1 vccd1 vccd1 _00353_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_1463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11559__B1 net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10421_ _03192_ _05190_ vssd1 vssd1 vccd1 vccd1 _05194_ sky130_fd_sc_hd__nor2_1
XFILLER_0_6_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13140_ clknet_leaf_12_clk _00371_ net1090 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[128\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_60_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10352_ net13 net1025 _05170_ final_design.data_from_mem\[1\] vssd1 vssd1 vccd1 vccd1
+ _00105_ sky130_fd_sc_hd__a22o_1
XANTENNA__10782__A1 net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10782__B2 net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13071_ clknet_leaf_42_clk _00302_ net1222 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[59\]
+ sky130_fd_sc_hd__dfrtp_1
X_10283_ _05139_ _05140_ vssd1 vssd1 vccd1 vccd1 _00029_ sky130_fd_sc_hd__nor2_1
XFILLER_0_63_1873 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12523__A2 net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12022_ _06224_ net290 net402 net2366 vssd1 vssd1 vccd1 vccd1 _00753_ sky130_fd_sc_hd__a22o_1
XANTENNA_input49_A mem_adr_start[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10534__A1 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_23_Right_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_50_1900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08669__B _02029_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_50_1911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14140__CLK clknet_leaf_17_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07065__S net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout570 net571 vssd1 vssd1 vccd1 vccd1 net570 sky130_fd_sc_hd__clkbuf_2
Xfanout581 net582 vssd1 vssd1 vccd1 vccd1 net581 sky130_fd_sc_hd__buf_2
Xfanout592 net593 vssd1 vssd1 vccd1 vccd1 net592 sky130_fd_sc_hd__clkbuf_8
XANTENNA__13708__CLK clknet_leaf_45_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13973_ clknet_leaf_57_clk _01204_ net1144 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[961\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12287__A1 net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12924_ clknet_leaf_49_clk _00162_ net1198 vssd1 vssd1 vccd1 vccd1 net147 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_17_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12039__A1 net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12855_ clknet_leaf_16_clk _00093_ net1109 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.ready_data\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_48_1840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06476__Y _01427_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1833 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_1328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13858__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11806_ net2487 net414 net288 _06068_ vssd1 vssd1 vccd1 vccd1 _00559_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_32_Right_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_44_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11798__B1 net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11737_ net229 net2176 net417 vssd1 vssd1 vccd1 vccd1 _00500_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11262__A2 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08663__B1 _02029_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11668_ net437 net579 _06191_ net300 net1559 vssd1 vssd1 vccd1 vccd1 _00466_ sky130_fd_sc_hd__a32o_1
XANTENNA__12882__CLK clknet_leaf_17_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13407_ clknet_leaf_7_clk _00638_ net1149 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[395\]
+ sky130_fd_sc_hd__dfrtp_1
X_10619_ net66 _05361_ vssd1 vssd1 vccd1 vccd1 _05363_ sky130_fd_sc_hd__nor2_1
XFILLER_0_25_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12146__S net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11599_ net437 net579 _06155_ net304 net1895 vssd1 vssd1 vccd1 vccd1 _00433_ sky130_fd_sc_hd__a32o_1
XFILLER_0_3_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07313__S1 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13338_ clknet_leaf_58_clk _00569_ net1132 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[326\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_38_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_38_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11970__B1 net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13238__CLK clknet_leaf_60_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13269_ clknet_leaf_56_clk _00500_ net1144 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[257\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_1913 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_41_Right_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12514__A2 net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11722__B1 net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07830_ final_design.cpu.reg_window\[469\] final_design.cpu.reg_window\[501\] net859
+ vssd1 vssd1 vccd1 vccd1 _02781_ sky130_fd_sc_hd__mux2_1
XANTENNA__13388__CLK clknet_leaf_45_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07761_ _02708_ _02709_ _02710_ _02711_ net686 net704 vssd1 vssd1 vccd1 vccd1 _02712_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__12278__A1 net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09500_ _04124_ _04418_ _04417_ net262 vssd1 vssd1 vccd1 vccd1 _04419_ sky130_fd_sc_hd__o211a_1
X_06712_ final_design.cpu.reg_window\[88\] final_design.cpu.reg_window\[120\] net942
+ vssd1 vssd1 vccd1 vccd1 _01663_ sky130_fd_sc_hd__mux2_1
X_07692_ _01599_ net615 vssd1 vssd1 vccd1 vccd1 _02643_ sky130_fd_sc_hd__or2_1
XFILLER_0_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_1739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09431_ _03585_ _03589_ vssd1 vssd1 vccd1 vccd1 _04350_ sky130_fd_sc_hd__or2_1
X_06643_ _01590_ _01591_ _01592_ _01593_ net775 net783 vssd1 vssd1 vccd1 vccd1 _01594_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__11733__B net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_50_Right_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06901__B1 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08329__S0 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09362_ _04158_ _04164_ _02738_ _04133_ vssd1 vssd1 vccd1 vccd1 _04281_ sky130_fd_sc_hd__a211o_1
X_06574_ final_design.cpu.reg_window\[989\] final_design.cpu.reg_window\[1021\] net949
+ vssd1 vssd1 vccd1 vccd1 _01525_ sky130_fd_sc_hd__mux2_1
X_08313_ final_design.cpu.reg_window\[328\] final_design.cpu.reg_window\[360\] net820
+ vssd1 vssd1 vccd1 vccd1 _03264_ sky130_fd_sc_hd__mux2_1
XANTENNA__06546__C net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07001__S0 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_2240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_1873 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09293_ _02641_ net445 _04206_ _04209_ vssd1 vssd1 vccd1 vccd1 _04212_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_60_2251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14240__1294 vssd1 vssd1 vccd1 vccd1 _14240__1294/HI net1294 sky130_fd_sc_hd__conb_1
XANTENNA_11 net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_2262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout236_A _05982_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_22 net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_2273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10461__B1 _05214_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08244_ net598 _03192_ _03168_ net538 vssd1 vssd1 vccd1 vccd1 _03195_ sky130_fd_sc_hd__o211a_1
XANTENNA__14013__CLK clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12202__A1 net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08175_ final_design.cpu.reg_window\[527\] final_design.cpu.reg_window\[559\] net806
+ vssd1 vssd1 vccd1 vccd1 _03126_ sky130_fd_sc_hd__mux2_1
XANTENNA__12056__S net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout403_A _06257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1145_A net1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07126_ _02073_ _02074_ _02075_ _02076_ net771 net790 vssd1 vssd1 vccd1 vccd1 _02077_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_82_1737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_1879 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_2180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11961__B1 net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11895__S net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_2191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07057_ net755 _02007_ vssd1 vssd1 vccd1 vccd1 _02008_ sky130_fd_sc_hd__nor2_1
XANTENNA__09873__B _04109_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14163__CLK clknet_leaf_17_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput140 net140 vssd1 vssd1 vccd1 vccd1 DAT_O[15] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_54_2044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput151 net151 vssd1 vssd1 vccd1 vccd1 DAT_O[25] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_54_2055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_2066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput162 net162 vssd1 vssd1 vccd1 vccd1 DAT_O[6] sky130_fd_sc_hd__buf_2
XANTENNA__12505__A2 net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput173 net173 vssd1 vssd1 vccd1 vccd1 gpio_out[1] sky130_fd_sc_hd__clkbuf_4
XANTENNA__07068__S0 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10812__B net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout772_A net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout393_X net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11196__A net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09382__A1 _04300_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07393__B1 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12269__A1 net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07959_ _02906_ _02907_ _02908_ _02909_ net683 net702 vssd1 vssd1 vccd1 vccd1 _02910_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout658_X net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10970_ net85 net1045 vssd1 vssd1 vccd1 vccd1 _05697_ sky130_fd_sc_hd__and2_1
XANTENNA__11643__B net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09629_ _02868_ _02898_ _04331_ vssd1 vssd1 vccd1 vccd1 _04548_ sky130_fd_sc_hd__and3b_1
XFILLER_0_74_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout825_X net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12640_ _06307_ net1413 net980 vssd1 vssd1 vccd1 vccd1 _01322_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12441__A1 net219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12571_ net2528 _06290_ _06286_ vssd1 vssd1 vccd1 vccd1 _01270_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_50_clk clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_50_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_38_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11522_ net2012 net199 net522 vssd1 vssd1 vccd1 vccd1 _00390_ sky130_fd_sc_hd__mux2_1
XANTENNA__07543__S1 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08444__S net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14241_ net1295 vssd1 vssd1 vccd1 vccd1 gpio_out[19] sky130_fd_sc_hd__buf_2
X_11453_ net239 net2255 net306 vssd1 vssd1 vccd1 vccd1 _00343_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10404_ _03450_ _05181_ vssd1 vssd1 vccd1 vccd1 _05185_ sky130_fd_sc_hd__nor2_1
X_14172_ clknet_leaf_20_clk _01346_ net1158 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.data_to_VGA\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11384_ net739 _03821_ _06069_ vssd1 vssd1 vccd1 vccd1 _06070_ sky130_fd_sc_hd__a21o_1
XANTENNA__10755__A1 _04040_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10755__B2 _04042_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11952__B1 net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13123_ clknet_leaf_0_clk _00354_ net1061 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[111\]
+ sky130_fd_sc_hd__dfrtp_1
X_10335_ net1542 net1009 net986 final_design.data_from_mem\[20\] vssd1 vssd1 vccd1
+ vccd1 _00092_ sky130_fd_sc_hd__a22o_1
X_13054_ clknet_leaf_13_clk _00285_ net1088 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[42\]
+ sky130_fd_sc_hd__dfrtp_1
X_10266_ final_design.uart.BAUD_counter\[24\] _05128_ net797 vssd1 vssd1 vccd1 vccd1
+ _05130_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_44_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11704__B1 net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12005_ _06207_ net285 net402 net2268 vssd1 vssd1 vccd1 vccd1 _00736_ sky130_fd_sc_hd__a22o_1
X_10197_ final_design.uart.BAUD_counter\[5\] final_design.uart.BAUD_counter\[4\] final_design.uart.BAUD_counter\[8\]
+ final_design.uart.BAUD_counter\[9\] vssd1 vssd1 vccd1 vccd1 _05086_ sky130_fd_sc_hd__or4b_1
XANTENNA__09125__A1 net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11393__X _06078_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13680__CLK clknet_leaf_36_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13956_ clknet_leaf_54_clk _01187_ net1178 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[944\]
+ sky130_fd_sc_hd__dfrtp_1
X_12907_ clknet_leaf_61_clk _00145_ net1140 vssd1 vssd1 vccd1 vccd1 net160 sky130_fd_sc_hd__dfrtp_1
XANTENNA__07231__S0 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13887_ clknet_leaf_7_clk _01118_ net1131 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[875\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11045__S net1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12838_ clknet_leaf_18_clk _00076_ net1111 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.ready_data\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14036__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07439__A1 net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11235__A2 _05936_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12432__A1 net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12769_ final_design.VGA_adr\[9\] net796 vssd1 vssd1 vccd1 vccd1 _01356_ sky130_fd_sc_hd__and2_1
XFILLER_0_51_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_41_clk clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_41_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_51_1084 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08862__B net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10443__B1 _05205_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput20 DAT_I[26] vssd1 vssd1 vccd1 vccd1 net20 sky130_fd_sc_hd__clkbuf_1
XANTENNA_clkbuf_leaf_20_clk_X clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput31 DAT_I[7] vssd1 vssd1 vccd1 vccd1 net31 sky130_fd_sc_hd__clkbuf_2
XANTENNA__13060__CLK clknet_leaf_54_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput42 mem_adr_start[15] vssd1 vssd1 vccd1 vccd1 net42 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput53 mem_adr_start[25] vssd1 vssd1 vccd1 vccd1 net53 sky130_fd_sc_hd__buf_1
XFILLER_0_64_1412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput64 mem_adr_start[6] vssd1 vssd1 vccd1 vccd1 net64 sky130_fd_sc_hd__buf_1
XFILLER_0_68_1592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput75 memory_size[16] vssd1 vssd1 vccd1 vccd1 net75 sky130_fd_sc_hd__buf_1
Xhold804 final_design.cpu.reg_window\[342\] vssd1 vssd1 vccd1 vccd1 net2146 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput86 memory_size[26] vssd1 vssd1 vccd1 vccd1 net86 sky130_fd_sc_hd__buf_2
XANTENNA__10746__A1 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold815 final_design.cpu.reg_window\[65\] vssd1 vssd1 vccd1 vccd1 net2157 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold826 final_design.cpu.reg_window\[860\] vssd1 vssd1 vccd1 vccd1 net2168 sky130_fd_sc_hd__dlygate4sd3_1
Xinput97 memory_size[7] vssd1 vssd1 vccd1 vccd1 net97 sky130_fd_sc_hd__buf_1
XANTENNA__11943__B1 net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold837 final_design.cpu.reg_window\[948\] vssd1 vssd1 vccd1 vccd1 net2179 sky130_fd_sc_hd__dlygate4sd3_1
Xhold848 final_design.cpu.reg_window\[565\] vssd1 vssd1 vccd1 vccd1 net2190 sky130_fd_sc_hd__dlygate4sd3_1
X_09980_ _03356_ _04706_ vssd1 vssd1 vccd1 vccd1 _04899_ sky130_fd_sc_hd__nand2_1
Xhold859 final_design.cpu.reg_window\[822\] vssd1 vssd1 vccd1 vccd1 net2201 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_35_clk_X clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08931_ _03758_ _03861_ vssd1 vssd1 vccd1 vccd1 _03873_ sky130_fd_sc_hd__nor2_1
XFILLER_0_58_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12901__Q net167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08862_ net1013 net254 vssd1 vssd1 vccd1 vccd1 _03812_ sky130_fd_sc_hd__or2_1
XFILLER_0_23_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_1817 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11171__A1 _04825_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07813_ _01660_ net615 vssd1 vssd1 vccd1 vccd1 _02764_ sky130_fd_sc_hd__nor2_1
X_08793_ _03680_ _03681_ vssd1 vssd1 vccd1 vccd1 _03744_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout186_A net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07744_ final_design.cpu.reg_window\[538\] final_design.cpu.reg_window\[570\] net861
+ vssd1 vssd1 vccd1 vccd1 _02695_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08529__S net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06838__A _01785_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08875__B1 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_2460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07675_ final_design.cpu.reg_window\[990\] final_design.cpu.reg_window\[1022\] net853
+ vssd1 vssd1 vccd1 vccd1 _02626_ sky130_fd_sc_hd__mux2_1
XANTENNA__12671__B2 final_design.data_from_mem\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_2471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout353_A net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06557__B _01507_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_2313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1095_A net1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09414_ _04331_ _04332_ net448 vssd1 vssd1 vccd1 vccd1 _04333_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_62_2324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07773__S1 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06626_ final_design.cpu.reg_window\[91\] final_design.cpu.reg_window\[123\] net943
+ vssd1 vssd1 vccd1 vccd1 _01577_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_81_2958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_2335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_2969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09345_ _04057_ _04076_ net474 vssd1 vssd1 vccd1 vccd1 _04264_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_1856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10029__A3 _04838_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06557_ _01453_ _01507_ vssd1 vssd1 vccd1 vccd1 _01508_ sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_32_clk clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_32_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__13403__CLK clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout618_A _02513_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_1889 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09276_ net88 _04194_ vssd1 vssd1 vccd1 vccd1 _04195_ sky130_fd_sc_hd__or2_2
XANTENNA__08264__S net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06488_ net755 _01430_ net747 vssd1 vssd1 vccd1 vccd1 _01439_ sky130_fd_sc_hd__o21a_1
XFILLER_0_74_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08227_ _03174_ _03175_ _03176_ _03177_ net681 net699 vssd1 vssd1 vccd1 vccd1 _03178_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout1050_X net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_2887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout406_X net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_2898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_2106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_2117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08158_ final_design.cpu.reg_window\[399\] final_design.cpu.reg_window\[431\] net810
+ vssd1 vssd1 vccd1 vccd1 _03109_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_56_2128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13553__CLK clknet_leaf_34_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout987_A _05167_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11934__B1 net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07109_ final_design.data_from_mem\[12\] net1039 net994 net991 vssd1 vssd1 vccd1
+ vccd1 _02060_ sky130_fd_sc_hd__or4_2
X_08089_ _02902_ _03033_ _03037_ _03039_ vssd1 vssd1 vccd1 vccd1 _03040_ sky130_fd_sc_hd__a211oi_2
X_10120_ _01370_ _05027_ _05029_ _04999_ vssd1 vssd1 vccd1 vccd1 final_design.vga.v_next_count\[6\]
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_41_1220 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout775_X net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10051_ _04654_ _04656_ _04700_ _04748_ _04749_ vssd1 vssd1 vccd1 vccd1 _04970_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_21_1849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout942_X net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07461__S0 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12771__2 clknet_leaf_25_clk vssd1 vssd1 vccd1 vccd1 net1312 sky130_fd_sc_hd__inv_2
X_13810_ clknet_leaf_44_clk _01041_ net1209 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[798\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14059__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13741_ clknet_leaf_48_clk _00972_ net1201 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[729\]
+ sky130_fd_sc_hd__dfrtp_1
X_10953_ _05680_ _05676_ vssd1 vssd1 vccd1 vccd1 _05681_ sky130_fd_sc_hd__and2b_1
XANTENNA__07213__S0 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13672_ clknet_leaf_40_clk _00903_ net1220 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[660\]
+ sky130_fd_sc_hd__dfrtp_1
X_10884_ _05613_ _05614_ vssd1 vssd1 vccd1 vccd1 _05615_ sky130_fd_sc_hd__nand2_1
X_12623_ final_design.VGA_data_control.state\[0\] final_design.VGA_data_control.state\[1\]
+ vssd1 vssd1 vccd1 vccd1 _06298_ sky130_fd_sc_hd__xor2_2
XFILLER_0_2_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13083__CLK clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_23_clk clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_23_clk sky130_fd_sc_hd__clkbuf_8
X_12554_ _06217_ net352 net325 net2291 vssd1 vssd1 vccd1 vccd1 _01258_ sky130_fd_sc_hd__a22o_1
XANTENNA__09291__A0 _01626_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11505_ net1865 net226 net521 vssd1 vssd1 vccd1 vccd1 _00374_ sky130_fd_sc_hd__mux2_1
X_12485_ _06145_ net357 net332 net2179 vssd1 vssd1 vccd1 vccd1 _01191_ sky130_fd_sc_hd__a22o_1
XFILLER_0_80_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14224_ final_design.pixel_data vssd1 vssd1 vccd1 vccd1 net174 sky130_fd_sc_hd__clkbuf_1
X_11436_ net1840 net186 net312 vssd1 vssd1 vccd1 vccd1 _00333_ sky130_fd_sc_hd__mux2_1
XANTENNA__11925__B1 net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14155_ clknet_leaf_18_clk _01329_ net1113 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.data_to_VGA\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_11367_ net739 _03837_ _06054_ vssd1 vssd1 vccd1 vccd1 _06055_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12920__CLK clknet_leaf_61_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13106_ clknet_leaf_39_clk _00337_ net1210 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[94\]
+ sky130_fd_sc_hd__dfrtp_1
X_10318_ net1512 net1012 net988 final_design.data_from_mem\[3\] vssd1 vssd1 vccd1
+ vccd1 _00075_ sky130_fd_sc_hd__a22o_1
XANTENNA__11548__B net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14086_ clknet_leaf_9_clk _01283_ net1151 vssd1 vssd1 vccd1 vccd1 final_design.reqhand.instruction\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_11298_ net643 _05994_ _05993_ vssd1 vssd1 vccd1 vccd1 _05995_ sky130_fd_sc_hd__a21o_1
XANTENNA__10452__B net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08149__A2 _03096_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13037_ clknet_leaf_44_clk _00268_ net1202 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_10249_ final_design.uart.BAUD_counter\[18\] _05118_ vssd1 vssd1 vccd1 vccd1 _05119_
+ sky130_fd_sc_hd__and2_1
XANTENNA__12350__B1 net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1140 net1141 vssd1 vssd1 vccd1 vccd1 net1140 sky130_fd_sc_hd__clkbuf_4
Xfanout1151 net1153 vssd1 vssd1 vccd1 vccd1 net1151 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_28_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1162 net1167 vssd1 vssd1 vccd1 vccd1 net1162 sky130_fd_sc_hd__clkbuf_4
Xfanout1173 net1175 vssd1 vssd1 vccd1 vccd1 net1173 sky130_fd_sc_hd__clkbuf_2
Xfanout1184 net1186 vssd1 vssd1 vccd1 vccd1 net1184 sky130_fd_sc_hd__clkbuf_4
Xfanout1195 net1197 vssd1 vssd1 vccd1 vccd1 net1195 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11564__A net209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13939_ clknet_leaf_41_clk _01170_ net1219 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[927\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12653__B2 final_design.data_from_mem\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_62_clk_A clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13426__CLK clknet_leaf_38_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10664__B1 net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07460_ final_design.cpu.reg_window\[896\] final_design.cpu.reg_window\[928\] net909
+ vssd1 vssd1 vccd1 vccd1 _02411_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_22_Left_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09321__X _04240_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06411_ final_design.CPU_instr_adr\[4\] vssd1 vssd1 vccd1 vccd1 _01366_ sky130_fd_sc_hd__inv_2
X_07391_ _02338_ _02339_ _02340_ _02341_ net770 net789 vssd1 vssd1 vccd1 vccd1 _02342_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_45_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_1821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11503__S net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_14_clk clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_14_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__10416__B1 _05191_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09130_ _02771_ _03594_ _03599_ vssd1 vssd1 vccd1 vccd1 _04049_ sky130_fd_sc_hd__a21boi_1
XANTENNA__09282__A0 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07489__A _02185_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13576__CLK clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09061_ net622 _03983_ _03985_ _03655_ vssd1 vssd1 vccd1 vccd1 _03989_ sky130_fd_sc_hd__o211a_1
XFILLER_0_60_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08012_ net613 _02961_ _02937_ net544 vssd1 vssd1 vccd1 vccd1 _02963_ sky130_fd_sc_hd__a211o_1
Xhold601 final_design.cpu.reg_window\[550\] vssd1 vssd1 vccd1 vccd1 net1943 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold612 final_design.cpu.reg_window\[146\] vssd1 vssd1 vccd1 vccd1 net1954 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_74_2740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold623 final_design.cpu.reg_window\[767\] vssd1 vssd1 vccd1 vccd1 net1965 sky130_fd_sc_hd__dlygate4sd3_1
Xhold634 final_design.cpu.reg_window\[56\] vssd1 vssd1 vccd1 vccd1 net1976 sky130_fd_sc_hd__dlygate4sd3_1
Xhold645 final_design.cpu.reg_window\[868\] vssd1 vssd1 vccd1 vccd1 net1987 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_31_Left_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_70_2604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold656 final_design.cpu.reg_window\[62\] vssd1 vssd1 vccd1 vccd1 net1998 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11392__A1 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold667 final_design.cpu.reg_window\[434\] vssd1 vssd1 vccd1 vccd1 net2009 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07428__S net913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09963_ _04851_ _04864_ vssd1 vssd1 vccd1 vccd1 _04882_ sky130_fd_sc_hd__xor2_1
XANTENNA__11458__B net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_4_Right_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold678 final_design.cpu.reg_window\[128\] vssd1 vssd1 vccd1 vccd1 net2020 sky130_fd_sc_hd__dlygate4sd3_1
Xhold689 final_design.cpu.reg_window\[412\] vssd1 vssd1 vccd1 vccd1 net2031 sky130_fd_sc_hd__dlygate4sd3_1
X_08914_ _02468_ _03856_ _03857_ net621 net257 vssd1 vssd1 vccd1 vccd1 _03858_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout1010_A _05166_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09894_ _03558_ _03559_ _03638_ vssd1 vssd1 vccd1 vccd1 _04813_ sky130_fd_sc_hd__and3_1
XANTENNA_clkbuf_leaf_15_clk_A clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12341__B1 net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08845_ final_design.CPU_instr_adr\[22\] final_design.CPU_instr_adr\[21\] _03795_
+ vssd1 vssd1 vccd1 vccd1 _03796_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout470_A _03485_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_2522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_2533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout568_A net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_2544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08776_ _03696_ _03726_ vssd1 vssd1 vccd1 vccd1 _03727_ sky130_fd_sc_hd__nor2_1
XANTENNA__06571__A1 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_2408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07727_ final_design.cpu.reg_window\[410\] final_design.cpu.reg_window\[442\] net864
+ vssd1 vssd1 vccd1 vccd1 _02678_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_40_Left_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout735_A net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout356_X net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07658_ _02608_ vssd1 vssd1 vccd1 vccd1 _02609_ sky130_fd_sc_hd__inv_2
XANTENNA__13919__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06609_ final_design.cpu.reg_window\[732\] final_design.cpu.reg_window\[764\] net946
+ vssd1 vssd1 vccd1 vccd1 _01560_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout523_X net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07589_ net878 _02521_ _02527_ _02533_ _02539_ vssd1 vssd1 vccd1 vccd1 _02540_ sky130_fd_sc_hd__o32a_4
XFILLER_0_14_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11413__S net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09328_ net321 _04052_ _04246_ vssd1 vssd1 vccd1 vccd1 _04247_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_11_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09812__A2 _04368_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09259_ net90 net93 net94 vssd1 vssd1 vccd1 vccd1 _04178_ sky130_fd_sc_hd__and3_1
XANTENNA__08171__S1 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12943__CLK clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12270_ net563 _06200_ net505 net368 net1664 vssd1 vssd1 vccd1 vccd1 _00985_ sky130_fd_sc_hd__a32o_1
XFILLER_0_62_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11907__A0 net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout892_X net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11221_ _04744_ net653 vssd1 vssd1 vccd1 vccd1 _05927_ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_1473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11383__A1 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09119__A net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11152_ _02358_ _05838_ net672 vssd1 vssd1 vccd1 vccd1 _05866_ sky130_fd_sc_hd__o21ai_4
XANTENNA__07682__S0 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10103_ final_design.VGA_data_control.v_count\[0\] _05017_ _05018_ vssd1 vssd1 vccd1
+ vccd1 final_design.vga.v_next_count\[0\] sky130_fd_sc_hd__o21a_1
X_11083_ net91 _05780_ vssd1 vssd1 vccd1 vccd1 _05805_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_8_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_8_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12332__B1 net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08536__C1 _02356_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input31_A DAT_I[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10034_ _04950_ _04952_ vssd1 vssd1 vccd1 vccd1 _04953_ sky130_fd_sc_hd__nor2_1
XFILLER_0_76_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11686__A2 net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08677__B _03617_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13449__CLK clknet_leaf_36_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_906 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11985_ _06187_ net291 net406 net1918 vssd1 vssd1 vccd1 vccd1 _00718_ sky130_fd_sc_hd__a22o_1
XANTENNA__11671__X _06194_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09500__A1 _04124_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10936_ _05643_ _05647_ _05664_ vssd1 vssd1 vccd1 vccd1 _05665_ sky130_fd_sc_hd__or3_1
X_13724_ clknet_leaf_2_clk _00955_ net1065 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[712\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13599__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10867_ net669 _05584_ _05598_ net966 _05597_ vssd1 vssd1 vccd1 vccd1 _05599_ sky130_fd_sc_hd__o221a_1
X_13655_ clknet_leaf_4_clk _00886_ net1084 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[643\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10287__X _05143_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12399__B1 net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12606_ net1477 net996 net982 final_design.data_from_mem\[24\] vssd1 vssd1 vccd1
+ vccd1 _01299_ sky130_fd_sc_hd__a22o_1
X_13586_ clknet_leaf_38_clk _00817_ net1205 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[574\]
+ sky130_fd_sc_hd__dfrtp_1
X_10798_ _05512_ _05514_ _05531_ vssd1 vssd1 vccd1 vccd1 _05533_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_67_1805 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12537_ _06200_ net346 net322 net1931 vssd1 vssd1 vccd1 vccd1 _01241_ sky130_fd_sc_hd__a22o_1
XANTENNA__11610__A2 net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12468_ _06128_ net346 net331 net2385 vssd1 vssd1 vccd1 vccd1 _01174_ sky130_fd_sc_hd__a22o_1
XFILLER_0_48_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09567__A1 net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14207_ net1265 vssd1 vssd1 vccd1 vccd1 gpio_oeb[19] sky130_fd_sc_hd__buf_2
X_11419_ net1744 net218 net310 vssd1 vssd1 vccd1 vccd1 _00316_ sky130_fd_sc_hd__mux2_1
XANTENNA__12154__S net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12399_ _06097_ net349 net339 net2155 vssd1 vssd1 vccd1 vccd1 _01109_ sky130_fd_sc_hd__a22o_1
XANTENNA__11374__A1 net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14138_ clknet_leaf_20_clk final_design.vga.h_next_count\[7\] net1159 vssd1 vssd1
+ vccd1 vccd1 final_design.VGA_data_control.VGA_request_address\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_1871 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06960_ _01908_ _01910_ vssd1 vssd1 vccd1 vccd1 _01911_ sky130_fd_sc_hd__and2_1
X_14069_ clknet_leaf_15_clk _00039_ net1095 vssd1 vssd1 vccd1 vccd1 final_design.uart.receiving
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_78_1901 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_3_clk clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_3_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_24_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06891_ _01838_ _01839_ _01840_ _01841_ net769 net790 vssd1 vssd1 vccd1 vccd1 _01842_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_20_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08630_ _03102_ _03580_ _03579_ vssd1 vssd1 vccd1 vccd1 _03581_ sky130_fd_sc_hd__a21o_1
XANTENNA__07976__S1 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08561_ net718 _03511_ vssd1 vssd1 vccd1 vccd1 _03512_ sky130_fd_sc_hd__or2_1
XFILLER_0_72_1522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07512_ _01825_ _02460_ _01790_ _01824_ vssd1 vssd1 vccd1 vccd1 _02463_ sky130_fd_sc_hd__o211a_1
XANTENNA__07728__S1 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06538__D _01480_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12779__10_A clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08492_ _03439_ _03440_ _03441_ _03442_ net677 net701 vssd1 vssd1 vccd1 vccd1 _03443_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_65_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07443_ _02391_ _02393_ vssd1 vssd1 vccd1 vccd1 _02394_ sky130_fd_sc_hd__nand2_2
XFILLER_0_58_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10638__A net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_983 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_21_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07374_ net882 _02318_ _02324_ _02311_ _02312_ vssd1 vssd1 vccd1 vccd1 _02325_ sky130_fd_sc_hd__a32oi_4
XFILLER_0_50_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_21_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09113_ _02419_ _02424_ net619 vssd1 vssd1 vccd1 vccd1 _04033_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_73_975 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_2802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11601__A2 net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_2813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout316_A net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1058_A final_design.reqhand.current_client\[3\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09044_ _03973_ _03968_ net259 vssd1 vssd1 vccd1 vccd1 _03974_ sky130_fd_sc_hd__mux2_1
XANTENNA__07947__A _01750_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06851__A net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold420 final_design.cpu.reg_window\[770\] vssd1 vssd1 vccd1 vccd1 net1762 sky130_fd_sc_hd__dlygate4sd3_1
Xhold431 final_design.cpu.reg_window\[598\] vssd1 vssd1 vccd1 vccd1 net1773 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11365__A1 net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08114__Y _03065_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold442 final_design.cpu.reg_window\[371\] vssd1 vssd1 vccd1 vccd1 net1784 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12562__B1 net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold453 final_design.cpu.reg_window\[927\] vssd1 vssd1 vccd1 vccd1 net1795 sky130_fd_sc_hd__dlygate4sd3_1
Xhold464 final_design.uart.working_data\[5\] vssd1 vssd1 vccd1 vccd1 net1806 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11188__B net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold475 final_design.cpu.reg_window\[515\] vssd1 vssd1 vccd1 vccd1 net1817 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold486 final_design.cpu.reg_window\[651\] vssd1 vssd1 vccd1 vccd1 net1828 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout900 net905 vssd1 vssd1 vccd1 vccd1 net900 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout685_A net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout911 net912 vssd1 vssd1 vccd1 vccd1 net911 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_1_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold497 final_design.cpu.reg_window\[79\] vssd1 vssd1 vccd1 vccd1 net1839 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout922 net953 vssd1 vssd1 vccd1 vccd1 net922 sky130_fd_sc_hd__buf_2
X_09946_ net530 net529 _02325_ net528 net452 net460 vssd1 vssd1 vccd1 vccd1 _04865_
+ sky130_fd_sc_hd__mux4_1
Xfanout933 net934 vssd1 vssd1 vccd1 vccd1 net933 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout1013_X net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout944 net945 vssd1 vssd1 vccd1 vccd1 net944 sky130_fd_sc_hd__clkbuf_4
Xfanout955 net957 vssd1 vssd1 vccd1 vccd1 net955 sky130_fd_sc_hd__clkbuf_4
Xfanout966 net967 vssd1 vssd1 vccd1 vccd1 net966 sky130_fd_sc_hd__clkbuf_4
Xfanout977 _06299_ vssd1 vssd1 vccd1 vccd1 net977 sky130_fd_sc_hd__clkbuf_2
XANTENNA__11668__A2 net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout852_A net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1120 final_design.cpu.reg_window\[319\] vssd1 vssd1 vccd1 vccd1 net2462 sky130_fd_sc_hd__dlygate4sd3_1
X_09877_ net529 net456 _04063_ vssd1 vssd1 vccd1 vccd1 _04796_ sky130_fd_sc_hd__a21o_1
Xfanout988 _05167_ vssd1 vssd1 vccd1 vccd1 net988 sky130_fd_sc_hd__clkbuf_4
Xfanout999 _06295_ vssd1 vssd1 vccd1 vccd1 net999 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08533__A2 _03481_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1131 final_design.reqhand.instruction\[10\] vssd1 vssd1 vccd1 vccd1 net2473 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10876__B1 net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1142 final_design.cpu.reg_window\[424\] vssd1 vssd1 vccd1 vccd1 net2484 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1153 final_design.cpu.reg_window\[99\] vssd1 vssd1 vccd1 vccd1 net2495 sky130_fd_sc_hd__dlygate4sd3_1
X_08828_ _03657_ _03778_ _03656_ vssd1 vssd1 vccd1 vccd1 _03779_ sky130_fd_sc_hd__a21o_1
Xhold1164 final_design.cpu.reg_window\[46\] vssd1 vssd1 vccd1 vccd1 net2506 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_79_Right_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1175 final_design.cpu.reg_window\[820\] vssd1 vssd1 vccd1 vccd1 net2517 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1186 final_design.uart.working_data\[4\] vssd1 vssd1 vccd1 vccd1 net2528 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout640_X net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13741__CLK clknet_leaf_48_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08759_ final_design.CPU_instr_adr\[3\] _02330_ vssd1 vssd1 vccd1 vccd1 _03710_ sky130_fd_sc_hd__or2_1
Xhold1197 final_design.cpu.reg_window\[61\] vssd1 vssd1 vccd1 vccd1 net2539 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout738_X net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11770_ _05848_ net568 vssd1 vssd1 vccd1 vccd1 _06228_ sky130_fd_sc_hd__nor2_8
XTAP_TAPCELL_ROW_0_172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12093__A2 _06090_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06585__X _01536_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12747__B net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10721_ _05436_ _05457_ vssd1 vssd1 vccd1 vccd1 _05460_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_0_194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11651__B net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout905_X net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13440_ clknet_leaf_10_clk _00671_ net1097 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[428\]
+ sky130_fd_sc_hd__dfrtp_1
X_10652_ _05389_ _05393_ vssd1 vssd1 vccd1 vccd1 _05394_ sky130_fd_sc_hd__xnor2_1
XANTENNA__11370__C _06057_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11053__B1 _05172_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13371_ clknet_leaf_64_clk _00602_ net1074 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[359\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09797__B2 _04086_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10583_ net1410 net1031 net1003 _05328_ vssd1 vssd1 vccd1 vccd1 _00179_ sky130_fd_sc_hd__a22o_1
X_12322_ net1919 net188 net366 vssd1 vssd1 vccd1 vccd1 _01036_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13121__CLK clknet_leaf_49_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input79_A memory_size[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09549__A1 _04342_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12253_ net573 _06182_ net507 net373 net1597 vssd1 vssd1 vccd1 vccd1 _00969_ sky130_fd_sc_hd__a32o_1
X_11204_ net426 net558 _05911_ net314 net2132 vssd1 vssd1 vccd1 vccd1 _00282_ sky130_fd_sc_hd__a32o_1
XANTENNA__12553__B1 net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12184_ net1870 net198 net382 vssd1 vssd1 vccd1 vccd1 _00903_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_1899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12953__RESET_B net1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13271__CLK clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11135_ _02358_ net803 net805 vssd1 vssd1 vccd1 vccd1 _05850_ sky130_fd_sc_hd__or3b_1
XANTENNA__14177__RESET_B net1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12839__CLK clknet_leaf_19_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input34_X net34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11066_ net959 _05785_ _05788_ _04042_ vssd1 vssd1 vccd1 vccd1 _05789_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__08040__X _02991_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10017_ net594 net659 _03611_ _03617_ vssd1 vssd1 vccd1 vccd1 _04936_ sky130_fd_sc_hd__or4bb_1
XTAP_TAPCELL_ROW_30_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_3006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_3017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10331__A2 net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_3028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_3039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06630__S1 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12497__X _06284_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12608__B2 final_design.data_from_mem\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12084__A2 net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11968_ _06170_ net278 net404 net1966 vssd1 vssd1 vccd1 vccd1 _00701_ sky130_fd_sc_hd__a22o_1
XFILLER_0_73_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_15_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13707_ clknet_leaf_52_clk _00938_ net1183 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[695\]
+ sky130_fd_sc_hd__dfrtp_1
X_10919_ _05647_ _05648_ net1397 net1033 vssd1 vssd1 vccd1 vccd1 _00195_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_15_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12149__S net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11899_ net207 net2042 net272 vssd1 vssd1 vccd1 vccd1 _00641_ sky130_fd_sc_hd__mux2_1
XANTENNA__10458__A _02570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13638_ clknet_leaf_50_clk _00869_ net1172 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[626\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13569_ clknet_leaf_47_clk _00800_ net1203 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[557\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11595__A1 net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07767__A net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07090_ final_design.cpu.reg_window\[204\] final_design.cpu.reg_window\[236\] net895
+ vssd1 vssd1 vccd1 vccd1 _02041_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13614__CLK clknet_leaf_44_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12544__B1 net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1857 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09800_ _03563_ _04718_ _03391_ vssd1 vssd1 vccd1 vccd1 _04719_ sky130_fd_sc_hd__o21ai_1
Xfanout207 net208 vssd1 vssd1 vccd1 vccd1 net207 sky130_fd_sc_hd__buf_2
XANTENNA__09960__A1 _04871_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout218 net219 vssd1 vssd1 vccd1 vccd1 net218 sky130_fd_sc_hd__clkbuf_2
X_07992_ final_design.cpu.reg_window\[80\] final_design.cpu.reg_window\[112\] net846
+ vssd1 vssd1 vccd1 vccd1 _02943_ sky130_fd_sc_hd__mux2_1
Xfanout229 _05864_ vssd1 vssd1 vccd1 vccd1 net229 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06943_ _01890_ _01891_ _01892_ _01893_ net772 net795 vssd1 vssd1 vccd1 vccd1 _01894_
+ sky130_fd_sc_hd__mux4_1
X_09731_ _04220_ _04408_ _04648_ _04649_ vssd1 vssd1 vccd1 vccd1 _04650_ sky130_fd_sc_hd__o211a_1
XANTENNA__13764__CLK clknet_leaf_54_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09662_ net487 _04578_ _04579_ _04580_ _04294_ vssd1 vssd1 vccd1 vccd1 _04581_ sky130_fd_sc_hd__a32o_1
XFILLER_0_74_1606 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06874_ net549 _01823_ vssd1 vssd1 vccd1 vccd1 _01825_ sky130_fd_sc_hd__xor2_1
XANTENNA__10322__A2 net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08613_ _03391_ _03563_ _03562_ vssd1 vssd1 vccd1 vccd1 _03564_ sky130_fd_sc_hd__a21o_1
X_09593_ _02770_ _04281_ _04168_ _02705_ vssd1 vssd1 vccd1 vccd1 _04512_ sky130_fd_sc_hd__o211ai_1
XANTENNA_fanout266_A net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08544_ final_design.cpu.reg_window\[1\] final_design.cpu.reg_window\[33\] net836
+ vssd1 vssd1 vccd1 vccd1 _03495_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_1461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1915 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12075__A2 _05959_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11471__B net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11283__B1 net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08475_ _03359_ _03425_ vssd1 vssd1 vccd1 vccd1 _03426_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout433_A _05847_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1175_A net1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07426_ final_design.cpu.reg_window\[833\] final_design.cpu.reg_window\[865\] net919
+ vssd1 vssd1 vccd1 vccd1 _02377_ sky130_fd_sc_hd__mux2_1
XANTENNA__13144__CLK clknet_leaf_65_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11898__S net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08126__S1 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07357_ final_design.cpu.reg_window\[195\] final_design.cpu.reg_window\[227\] net901
+ vssd1 vssd1 vccd1 vccd1 _02308_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout221_X net221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout600_A net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10389__A2 net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout319_X net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07288_ net882 _02238_ _02227_ _02221_ vssd1 vssd1 vccd1 vccd1 _02239_ sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_33_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09027_ final_design.CPU_instr_adr\[12\] net1017 _03956_ _03958_ vssd1 vssd1 vccd1
+ vccd1 _00223_ sky130_fd_sc_hd__a22o_1
XANTENNA__11199__A net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13294__CLK clknet_leaf_43_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12535__B1 net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold250 final_design.cpu.reg_window\[783\] vssd1 vssd1 vccd1 vccd1 net1592 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07637__S0 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold261 final_design.cpu.reg_window\[153\] vssd1 vssd1 vccd1 vccd1 net1603 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout590_X net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout688_X net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold272 final_design.cpu.reg_window\[975\] vssd1 vssd1 vccd1 vccd1 net1614 sky130_fd_sc_hd__dlygate4sd3_1
Xhold283 final_design.cpu.reg_window\[904\] vssd1 vssd1 vccd1 vccd1 net1625 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10010__A1 _02326_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold294 final_design.cpu.reg_window\[771\] vssd1 vssd1 vccd1 vccd1 net1636 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout730 _01492_ vssd1 vssd1 vccd1 vccd1 net730 sky130_fd_sc_hd__buf_4
Xfanout741 _01477_ vssd1 vssd1 vccd1 vccd1 net741 sky130_fd_sc_hd__clkbuf_4
X_09929_ _04178_ _04829_ _04847_ vssd1 vssd1 vccd1 vccd1 _04848_ sky130_fd_sc_hd__or3b_1
Xfanout752 _01427_ vssd1 vssd1 vccd1 vccd1 net752 sky130_fd_sc_hd__buf_4
Xfanout763 _01426_ vssd1 vssd1 vccd1 vccd1 net763 sky130_fd_sc_hd__buf_4
XANTENNA_fanout855_X net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout774 net778 vssd1 vssd1 vccd1 vccd1 net774 sky130_fd_sc_hd__buf_4
XANTENNA__08506__A2 _03450_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout785 net788 vssd1 vssd1 vccd1 vccd1 net785 sky130_fd_sc_hd__clkbuf_4
Xfanout796 _06333_ vssd1 vssd1 vccd1 vccd1 net796 sky130_fd_sc_hd__clkbuf_4
X_12940_ clknet_leaf_22_clk _00178_ net1163 vssd1 vssd1 vccd1 vccd1 net128 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_77_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11510__A1 net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07562__D net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10977__S net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12871_ clknet_leaf_25_clk _00109_ net1152 vssd1 vssd1 vccd1 vccd1 final_design.data_from_mem\[5\]
+ sky130_fd_sc_hd__dfrtp_4
X_11822_ net215 net2065 net265 vssd1 vssd1 vccd1 vccd1 _00574_ sky130_fd_sc_hd__mux2_1
XANTENNA__08447__S net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07351__S net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11753_ net204 net2154 net418 vssd1 vssd1 vccd1 vccd1 _00516_ sky130_fd_sc_hd__mux2_1
XANTENNA__11274__B1 net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10704_ net1003 _05442_ _05443_ net1032 net1373 vssd1 vssd1 vccd1 vccd1 _00185_ sky130_fd_sc_hd__a32o_1
XFILLER_0_16_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09482__A3 net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11684_ net563 net421 _06200_ net294 net1980 vssd1 vssd1 vccd1 vccd1 _00473_ sky130_fd_sc_hd__a32o_1
XANTENNA__13152__RESET_B net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_42_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10635_ final_design.CPU_instr_adr\[9\] _05377_ net1054 vssd1 vssd1 vccd1 vccd1 _05378_
+ sky130_fd_sc_hd__mux2_1
X_13423_ clknet_leaf_38_clk _00654_ net1190 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[411\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_42_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11577__A1 net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13637__CLK clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13354_ clknet_leaf_51_clk _00585_ net1170 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[342\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1917 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10566_ net96 final_design.VGA_adr\[4\] vssd1 vssd1 vccd1 vccd1 _05312_ sky130_fd_sc_hd__or2_1
XFILLER_0_64_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12305_ net1616 net221 net364 vssd1 vssd1 vccd1 vccd1 _01019_ sky130_fd_sc_hd__mux2_1
X_13285_ clknet_leaf_48_clk _00516_ net1185 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[273\]
+ sky130_fd_sc_hd__dfrtp_1
X_10497_ _05233_ _05246_ vssd1 vssd1 vccd1 vccd1 _05247_ sky130_fd_sc_hd__or2_1
XFILLER_0_62_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12526__B1 net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11329__B2 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12236_ net564 _06166_ net505 net372 net1434 vssd1 vssd1 vccd1 vccd1 _00953_ sky130_fd_sc_hd__a32o_1
XFILLER_0_20_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13787__CLK clknet_leaf_65_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14199__1257 vssd1 vssd1 vccd1 vccd1 _14199__1257/HI net1257 sky130_fd_sc_hd__conb_1
XFILLER_0_27_1685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_1696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12167_ net2282 net226 net381 vssd1 vssd1 vccd1 vccd1 _00886_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_36_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12432__S net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11118_ final_design.uart.bits_received\[0\] final_design.uart.bits_received\[1\]
+ final_design.uart.bits_received\[2\] final_design.uart.bits_received\[3\] vssd1
+ vssd1 vccd1 vccd1 _05835_ sky130_fd_sc_hd__a31o_1
XFILLER_0_78_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11556__B net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12098_ net1974 net226 net389 vssd1 vssd1 vccd1 vccd1 _00822_ sky130_fd_sc_hd__mux2_1
XANTENNA__10460__B net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13017__CLK clknet_leaf_56_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11049_ _01387_ _05772_ vssd1 vssd1 vccd1 vccd1 _05773_ sky130_fd_sc_hd__nor2_1
Xinput7 DAT_I[14] vssd1 vssd1 vccd1 vccd1 net7 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08865__B _01538_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06590_ _01536_ _01539_ vssd1 vssd1 vccd1 vccd1 _01541_ sky130_fd_sc_hd__nand2_1
XANTENNA__13167__CLK clknet_leaf_42_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09042__A net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08356__S1 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11804__A2 net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08260_ _03207_ _03208_ _03209_ _03210_ net675 net697 vssd1 vssd1 vccd1 vccd1 _03211_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__08681__A1 _02545_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07211_ final_design.cpu.reg_window\[456\] final_design.cpu.reg_window\[488\] net891
+ vssd1 vssd1 vccd1 vccd1 _02162_ sky130_fd_sc_hd__mux2_1
X_08191_ final_design.cpu.reg_window\[78\] final_design.cpu.reg_window\[110\] net812
+ vssd1 vssd1 vccd1 vccd1 _03142_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11511__S net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07142_ _01468_ net734 net836 vssd1 vssd1 vccd1 vccd1 _02093_ sky130_fd_sc_hd__and3_1
XANTENNA__08092__S net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08433__B2 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07073_ _02020_ _02021_ _02022_ _02023_ net774 net792 vssd1 vssd1 vccd1 vccd1 _02024_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__12690__X _06333_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12517__B1 net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_691 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_40 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08292__S0 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07975_ final_design.cpu.reg_window\[529\] final_design.cpu.reg_window\[561\] net845
+ vssd1 vssd1 vccd1 vccd1 _02926_ sky130_fd_sc_hd__mux2_1
X_09714_ net72 _04184_ vssd1 vssd1 vccd1 vccd1 _04633_ sky130_fd_sc_hd__nand2_1
X_06926_ final_design.cpu.reg_window\[530\] final_design.cpu.reg_window\[562\] net924
+ vssd1 vssd1 vccd1 vccd1 _01877_ sky130_fd_sc_hd__mux2_1
XANTENNA__07960__A net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09792__S0 net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06857_ net754 _01807_ vssd1 vssd1 vccd1 vccd1 _01808_ sky130_fd_sc_hd__nor2_1
X_09645_ _04218_ _04563_ _04556_ net261 _04558_ vssd1 vssd1 vccd1 vccd1 _04564_ sky130_fd_sc_hd__o2111ai_1
XANTENNA_fanout550_A _01784_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12578__A net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13663__RESET_B net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout269_X net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout648_A _05849_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09576_ _03295_ _03569_ _03576_ vssd1 vssd1 vccd1 vccd1 _04495_ sky130_fd_sc_hd__a21o_1
XFILLER_0_78_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06788_ final_design.cpu.reg_window\[534\] final_design.cpu.reg_window\[566\] net920
+ vssd1 vssd1 vccd1 vccd1 _01739_ sky130_fd_sc_hd__mux2_1
XANTENNA__08267__S net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14092__CLK clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08527_ final_design.cpu.reg_window\[514\] final_design.cpu.reg_window\[546\] net832
+ vssd1 vssd1 vccd1 vccd1 _03478_ sky130_fd_sc_hd__mux2_1
XANTENNA__11256__B1 _05843_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1887 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout436_X net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout815_A net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08458_ final_design.cpu.reg_window\[708\] final_design.cpu.reg_window\[740\] net819
+ vssd1 vssd1 vccd1 vccd1 _03409_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11008__B1 net1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07409_ net740 _02358_ vssd1 vssd1 vccd1 vccd1 _02360_ sky130_fd_sc_hd__nand2_1
XFILLER_0_68_1218 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08389_ net709 _03333_ net722 vssd1 vssd1 vccd1 vccd1 _03340_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout603_X net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11559__A1 net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11421__S net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10420_ net1796 net1031 _05193_ net246 vssd1 vssd1 vccd1 vccd1 _00151_ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10351_ net2 net1023 net1007 final_design.data_from_mem\[0\] vssd1 vssd1 vccd1 vccd1
+ _00104_ sky130_fd_sc_hd__o22a_1
XANTENNA__06986__A1 net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12508__B1 net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08015__B net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13070_ clknet_leaf_45_clk _00301_ net1213 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[58\]
+ sky130_fd_sc_hd__dfrtp_1
X_10282_ net2530 _05138_ net798 vssd1 vssd1 vccd1 vccd1 _05140_ sky130_fd_sc_hd__o21ai_1
X_12021_ _06223_ net292 net402 net2325 vssd1 vssd1 vccd1 vccd1 _00752_ sky130_fd_sc_hd__a22o_1
XFILLER_0_63_1885 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10561__A net1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09127__A net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08669__C _02061_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_1347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout560 net561 vssd1 vssd1 vccd1 vccd1 net560 sky130_fd_sc_hd__buf_2
XFILLER_0_79_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout571 _05868_ vssd1 vssd1 vccd1 vccd1 net571 sky130_fd_sc_hd__buf_4
Xfanout582 net583 vssd1 vssd1 vccd1 vccd1 net582 sky130_fd_sc_hd__clkbuf_4
Xfanout593 _05199_ vssd1 vssd1 vccd1 vccd1 net593 sky130_fd_sc_hd__clkbuf_8
X_13972_ clknet_leaf_8_clk _01203_ net1153 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[960\]
+ sky130_fd_sc_hd__dfrtp_1
X_12923_ clknet_leaf_30_clk _00161_ net1233 vssd1 vssd1 vccd1 vccd1 net146 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_17_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12854_ clknet_leaf_16_clk _00092_ net1096 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.ready_data\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_1801 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08177__S net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13333__RESET_B net1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_1852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11805_ net2362 net414 net291 _06061_ vssd1 vssd1 vccd1 vccd1 _00558_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_48_1863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11247__B1 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1845 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_1889 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11736_ net230 net2508 net416 vssd1 vssd1 vccd1 vccd1 _00499_ sky130_fd_sc_hd__mux2_1
XANTENNA__08663__A1 _01999_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10736__A net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11667_ net176 net632 vssd1 vssd1 vccd1 vccd1 _06191_ sky130_fd_sc_hd__and2_1
X_13406_ clknet_leaf_10_clk _00637_ net1100 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[394\]
+ sky130_fd_sc_hd__dfrtp_1
X_10618_ net66 _05361_ vssd1 vssd1 vccd1 vccd1 _05362_ sky130_fd_sc_hd__and2_1
XFILLER_0_3_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11598_ net179 net636 vssd1 vssd1 vccd1 vccd1 _06155_ sky130_fd_sc_hd__and2_1
XANTENNA__08966__A2 net1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10549_ final_design.CPU_instr_adr\[5\] _05277_ vssd1 vssd1 vccd1 vccd1 _05296_ sky130_fd_sc_hd__or2_1
X_13337_ clknet_leaf_55_clk _00568_ net1148 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[325\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_38_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13268_ clknet_leaf_9_clk _00499_ net1104 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[256\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12219_ net570 _06147_ net507 net377 net1993 vssd1 vssd1 vccd1 vccd1 _00937_ sky130_fd_sc_hd__a32o_1
X_13199_ clknet_leaf_42_clk _00430_ net1220 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[187\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11722__A1 net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09391__A2 _04309_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07760_ final_design.cpu.reg_window\[408\] final_design.cpu.reg_window\[440\] net864
+ vssd1 vssd1 vccd1 vccd1 _02711_ sky130_fd_sc_hd__mux2_1
XANTENNA__08026__S0 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09679__B1 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06711_ _01658_ _01660_ vssd1 vssd1 vccd1 vccd1 _01662_ sky130_fd_sc_hd__and2_1
XFILLER_0_79_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07691_ _02543_ _02544_ _02637_ _02639_ vssd1 vssd1 vccd1 vccd1 _02642_ sky130_fd_sc_hd__o22a_1
XFILLER_0_56_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11506__S net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09430_ net496 _04348_ _04231_ vssd1 vssd1 vccd1 vccd1 _04349_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_56_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06642_ final_design.cpu.reg_window\[539\] final_design.cpu.reg_window\[571\] net941
+ vssd1 vssd1 vccd1 vccd1 _01593_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13802__CLK clknet_leaf_59_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06901__A1 _01468_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08329__S1 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09361_ _04046_ _04255_ _04256_ _04279_ vssd1 vssd1 vccd1 vccd1 _04280_ sky130_fd_sc_hd__a31o_1
X_06573_ final_design.cpu.reg_window\[797\] final_design.cpu.reg_window\[829\] net950
+ vssd1 vssd1 vccd1 vccd1 _01524_ sky130_fd_sc_hd__mux2_1
XANTENNA__10349__C net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08312_ _02186_ net598 vssd1 vssd1 vccd1 vccd1 _03263_ sky130_fd_sc_hd__nand2_1
XANTENNA__11789__B2 net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09292_ _01626_ _01657_ net552 _01717_ net458 net467 vssd1 vssd1 vccd1 vccd1 _04211_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__07001__S1 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1705 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_2241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_9_clk_X clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_2252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_1885 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_12 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_2263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10461__A1 net157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13952__CLK clknet_leaf_11_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_23 _06257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08243_ net598 _03192_ _03168_ vssd1 vssd1 vccd1 vccd1 _03194_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_6_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10461__B2 net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_1749 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12738__B1 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08174_ final_design.cpu.reg_window\[591\] final_design.cpu.reg_window\[623\] net806
+ vssd1 vssd1 vccd1 vccd1 _03125_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07125_ final_design.cpu.reg_window\[139\] final_design.cpu.reg_window\[171\] net915
+ vssd1 vssd1 vccd1 vccd1 _02076_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_1749 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_2181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07056_ _02003_ _02004_ _02005_ _02006_ net772 net791 vssd1 vssd1 vccd1 vccd1 _02007_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_30_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_2192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput130 net130 vssd1 vssd1 vccd1 vccd1 ADR_O[7] sky130_fd_sc_hd__clkbuf_4
Xoutput141 net141 vssd1 vssd1 vccd1 vccd1 DAT_O[16] sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_54_2045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput152 net152 vssd1 vssd1 vccd1 vccd1 DAT_O[26] sky130_fd_sc_hd__buf_2
XANTENNA__09906__A1 _04072_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_2056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout598_A net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput163 net163 vssd1 vssd1 vccd1 vccd1 DAT_O[7] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_54_2067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07068__S1 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput174 net174 vssd1 vssd1 vccd1 vccd1 gpio_out[2] sky130_fd_sc_hd__buf_2
XANTENNA__07166__S net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13332__CLK clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07393__A1 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout386_X net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout765_A net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13844__RESET_B net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07958_ final_design.cpu.reg_window\[401\] final_design.cpu.reg_window\[433\] net848
+ vssd1 vssd1 vccd1 vccd1 _02909_ sky130_fd_sc_hd__mux2_1
X_06909_ final_design.cpu.reg_window\[402\] final_design.cpu.reg_window\[434\] net924
+ vssd1 vssd1 vccd1 vccd1 _01860_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_1905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07889_ final_design.cpu.reg_window\[343\] final_design.cpu.reg_window\[375\] net851
+ vssd1 vssd1 vccd1 vccd1 _02840_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout932_A net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout553_X net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11416__S net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13482__CLK clknet_leaf_51_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09628_ _02898_ _04331_ vssd1 vssd1 vccd1 vccd1 _04547_ sky130_fd_sc_hd__nand2_1
XANTENNA__11229__B1 net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09559_ _04452_ _04455_ _04477_ _04425_ vssd1 vssd1 vccd1 vccd1 _04478_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout720_X net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_7_0_clk_X clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout818_X net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14198__1256 vssd1 vssd1 vccd1 vccd1 _14198__1256/HI net1256 sky130_fd_sc_hd__conb_1
XFILLER_0_77_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12570_ final_design.uart.receiving final_design.uart.working_data\[5\] vssd1 vssd1
+ vccd1 vccd1 _06290_ sky130_fd_sc_hd__and2_1
XFILLER_0_38_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11521_ net1954 net201 net523 vssd1 vssd1 vccd1 vccd1 _00389_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06751__S0 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14240_ net1294 vssd1 vssd1 vccd1 vccd1 gpio_out[18] sky130_fd_sc_hd__buf_2
X_11452_ net239 net638 vssd1 vssd1 vccd1 vccd1 _06099_ sky130_fd_sc_hd__and2_1
XFILLER_0_34_742 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08671__D _01659_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10403_ net2463 net1027 _05184_ net246 vssd1 vssd1 vccd1 vccd1 _00143_ sky130_fd_sc_hd__a22o_1
X_14171_ clknet_leaf_19_clk _01345_ net1157 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.data_to_VGA\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09070__A1 _03655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11383_ net661 _03815_ _01491_ vssd1 vssd1 vccd1 vccd1 _06069_ sky130_fd_sc_hd__o21a_1
XANTENNA__11952__A1 _06153_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input61_A mem_adr_start[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13122_ clknet_leaf_3_clk _00353_ net1068 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[110\]
+ sky130_fd_sc_hd__dfrtp_1
X_10334_ net1529 net1011 net988 final_design.data_from_mem\[19\] vssd1 vssd1 vccd1
+ vccd1 _00091_ sky130_fd_sc_hd__a22o_1
X_13053_ clknet_leaf_2_clk _00284_ net1064 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[41\]
+ sky130_fd_sc_hd__dfrtp_1
X_10265_ final_design.uart.BAUD_counter\[24\] _05128_ vssd1 vssd1 vccd1 vccd1 _05129_
+ sky130_fd_sc_hd__and2_1
XANTENNA__09128__Y _04047_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11704__A1 net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12004_ _06206_ net278 net400 net2340 vssd1 vssd1 vccd1 vccd1 _00735_ sky130_fd_sc_hd__a22o_1
X_10196_ final_design.uart.BAUD_counter\[11\] final_design.uart.BAUD_counter\[10\]
+ final_design.uart.bits_received\[2\] final_design.uart.bits_received\[3\] vssd1
+ vssd1 vccd1 vccd1 _05085_ sky130_fd_sc_hd__or4_1
XANTENNA__08008__S0 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13825__CLK clknet_leaf_47_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09291__S net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout390 net391 vssd1 vssd1 vccd1 vccd1 net390 sky130_fd_sc_hd__clkbuf_8
XANTENNA__09125__A2 net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07804__S net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13955_ clknet_leaf_1_clk _01186_ net1071 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[943\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06487__Y _01438_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12906_ clknet_leaf_61_clk _00144_ net1136 vssd1 vssd1 vccd1 vccd1 net159 sky130_fd_sc_hd__dfrtp_1
XANTENNA__07231__S1 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13886_ clknet_leaf_9_clk _01117_ net1103 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[874\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_801 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13975__CLK clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12837_ clknet_leaf_19_clk _00075_ net1156 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.ready_data\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1030 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_867 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08636__A1 net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12768_ final_design.VGA_adr\[8\] net796 _06402_ net954 vssd1 vssd1 vccd1 vccd1 _01355_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__06944__A net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10757__A2_N net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11719_ net190 net628 vssd1 vssd1 vccd1 vccd1 _06218_ sky130_fd_sc_hd__and2_1
XANTENNA__11640__B1 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10443__B2 net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12157__S net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13205__CLK clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12699_ final_design.VGA_data_control.v_count\[5\] _06339_ vssd1 vssd1 vccd1 vccd1
+ _06340_ sky130_fd_sc_hd__xnor2_1
Xinput10 DAT_I[17] vssd1 vssd1 vccd1 vccd1 net10 sky130_fd_sc_hd__clkbuf_1
Xinput21 DAT_I[27] vssd1 vssd1 vccd1 vccd1 net21 sky130_fd_sc_hd__clkbuf_1
Xinput32 DAT_I[8] vssd1 vssd1 vccd1 vccd1 net32 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_68_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput43 mem_adr_start[16] vssd1 vssd1 vccd1 vccd1 net43 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_1402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput54 mem_adr_start[26] vssd1 vssd1 vccd1 vccd1 net54 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_40_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput65 mem_adr_start[7] vssd1 vssd1 vccd1 vccd1 net65 sky130_fd_sc_hd__clkbuf_1
XANTENNA__09061__A1 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold805 final_design.cpu.reg_window\[498\] vssd1 vssd1 vccd1 vccd1 net2147 sky130_fd_sc_hd__dlygate4sd3_1
Xinput76 memory_size[17] vssd1 vssd1 vccd1 vccd1 net76 sky130_fd_sc_hd__clkbuf_2
Xhold816 final_design.cpu.reg_window\[391\] vssd1 vssd1 vccd1 vccd1 net2158 sky130_fd_sc_hd__dlygate4sd3_1
Xinput87 memory_size[27] vssd1 vssd1 vccd1 vccd1 net87 sky130_fd_sc_hd__buf_1
XANTENNA__10746__A2 _04509_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput98 memory_size[8] vssd1 vssd1 vccd1 vccd1 net98 sky130_fd_sc_hd__buf_1
XFILLER_0_64_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold827 final_design.cpu.reg_window\[582\] vssd1 vssd1 vccd1 vccd1 net2169 sky130_fd_sc_hd__dlygate4sd3_1
Xhold838 final_design.cpu.reg_window\[180\] vssd1 vssd1 vccd1 vccd1 net2180 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13355__CLK clknet_leaf_38_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold849 final_design.cpu.reg_window\[477\] vssd1 vssd1 vccd1 vccd1 net2191 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08930_ _01789_ _02463_ _01759_ vssd1 vssd1 vccd1 vccd1 _03872_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_81_1793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12499__A2 net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08861_ _03802_ _03810_ vssd1 vssd1 vccd1 vccd1 _03811_ sky130_fd_sc_hd__and2_1
XANTENNA__07375__A1 net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_1829 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07812_ _02750_ _02751_ _02762_ net878 vssd1 vssd1 vccd1 vccd1 _02763_ sky130_fd_sc_hd__a22oi_4
X_08792_ _03688_ _03732_ _03742_ _03687_ vssd1 vssd1 vccd1 vccd1 _03743_ sky130_fd_sc_hd__and4b_1
XANTENNA__12620__S _05080_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07714__S net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07743_ final_design.cpu.reg_window\[602\] final_design.cpu.reg_window\[634\] net856
+ vssd1 vssd1 vccd1 vccd1 _02694_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12120__A1 net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08324__B1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout179_A _06081_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09667__A3 _04579_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06838__B _01788_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_2450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07674_ final_design.cpu.reg_window\[798\] final_design.cpu.reg_window\[830\] net855
+ vssd1 vssd1 vccd1 vccd1 _02625_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_66_2461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_66_2472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06625_ _01572_ _01573_ _01574_ _01575_ net776 net793 vssd1 vssd1 vccd1 vccd1 _01576_
+ sky130_fd_sc_hd__mux4_1
X_09413_ _02804_ _04330_ _04131_ _02900_ vssd1 vssd1 vccd1 vccd1 _04332_ sky130_fd_sc_hd__o211ai_1
XTAP_TAPCELL_ROW_62_2314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_2325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_2959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_2336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout346_A net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1088_A net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09344_ _04261_ _04262_ net496 _04097_ vssd1 vssd1 vccd1 vccd1 _04263_ sky130_fd_sc_hd__a211o_1
X_06556_ net741 _01497_ net665 _01506_ vssd1 vssd1 vccd1 vccd1 _01507_ sky130_fd_sc_hd__a211o_4
XANTENNA__12423__A2 _06264_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08545__S net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09275_ net86 net87 _04193_ vssd1 vssd1 vccd1 vccd1 _04194_ sky130_fd_sc_hd__or3_1
XFILLER_0_30_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06487_ net884 vssd1 vssd1 vccd1 vccd1 _01438_ sky130_fd_sc_hd__clkinv_4
XANTENNA_fanout513_A net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14130__CLK clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06733__S0 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08226_ final_design.cpu.reg_window\[139\] final_design.cpu.reg_window\[171\] net836
+ vssd1 vssd1 vccd1 vccd1 _03177_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07850__A2 _02797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_2888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_2899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08157_ final_design.cpu.reg_window\[463\] final_design.cpu.reg_window\[495\] net810
+ vssd1 vssd1 vccd1 vccd1 _03108_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_56_2107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout301_X net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_2118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_2129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07108_ net882 _02051_ _02057_ _02044_ _02045_ vssd1 vssd1 vccd1 vccd1 _02059_ sky130_fd_sc_hd__a32o_4
XANTENNA__07063__B1 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07685__A _01507_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08088_ _01718_ _02839_ _02864_ _02868_ _03038_ vssd1 vssd1 vccd1 vccd1 _03039_ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout882_A net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07039_ final_design.cpu.reg_window\[526\] final_design.cpu.reg_window\[558\] net894
+ vssd1 vssd1 vccd1 vccd1 _01990_ sky130_fd_sc_hd__mux2_1
XANTENNA__11000__A net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10050_ _04919_ _04921_ _04922_ _04968_ _04476_ vssd1 vssd1 vccd1 vccd1 _04969_ sky130_fd_sc_hd__o2111a_1
XANTENNA__08012__C1 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11698__B1 net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout670_X net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11162__A2 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout768_X net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06588__X _01539_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10370__B1 net1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07461__S1 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13998__CLK clknet_leaf_43_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12872__CLK clknet_leaf_25_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout935_X net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13740_ clknet_leaf_46_clk _00971_ net1214 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[728\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10952_ net84 _05651_ _05679_ vssd1 vssd1 vccd1 vccd1 _05680_ sky130_fd_sc_hd__a21o_1
XANTENNA__07213__S1 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13671_ clknet_leaf_63_clk _00902_ net1119 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[659\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11870__B1 net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10883_ _05590_ _05593_ _05611_ _05612_ vssd1 vssd1 vccd1 vccd1 _05614_ sky130_fd_sc_hd__o211ai_1
XANTENNA__13228__CLK clknet_leaf_46_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11670__A net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12622_ final_design.VGA_data_control.state\[1\] _01402_ final_design.VGA_data_control.state\[0\]
+ vssd1 vssd1 vccd1 vccd1 _06297_ sky130_fd_sc_hd__o21a_1
XANTENNA__12414__A2 net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12553_ _06216_ net348 net323 net2148 vssd1 vssd1 vccd1 vccd1 _01257_ sky130_fd_sc_hd__a22o_1
XANTENNA__11622__B1 net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09291__A1 _01657_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11504_ net2005 net242 net522 vssd1 vssd1 vccd1 vccd1 _00373_ sky130_fd_sc_hd__mux2_1
X_12484_ _06144_ net349 net331 net2017 vssd1 vssd1 vccd1 vccd1 _01190_ sky130_fd_sc_hd__a22o_1
XANTENNA__13378__CLK clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12178__A1 net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14223_ final_design.v_out vssd1 vssd1 vccd1 vccd1 net173 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_80_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11669__X _06192_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11435_ net1805 net189 net312 vssd1 vssd1 vccd1 vccd1 _00332_ sky130_fd_sc_hd__mux2_1
XANTENNA__09139__X _04058_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07595__A _01539_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14154_ clknet_leaf_18_clk _01328_ net1108 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.data_to_VGA\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_11366_ net661 _03832_ net733 vssd1 vssd1 vccd1 vccd1 _06054_ sky130_fd_sc_hd__o21a_1
XANTENNA__11388__Y _06074_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06703__S net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10317_ net1487 net1011 net989 final_design.data_from_mem\[2\] vssd1 vssd1 vccd1
+ vccd1 _00074_ sky130_fd_sc_hd__a22o_1
X_13105_ clknet_leaf_34_clk _00336_ net1242 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[93\]
+ sky130_fd_sc_hd__dfrtp_1
X_14085_ clknet_leaf_25_clk _01282_ net1151 vssd1 vssd1 vccd1 vccd1 final_design.reqhand.instruction\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_11297_ final_design.data_from_mem\[18\] net235 net233 vssd1 vssd1 vccd1 vccd1 _05994_
+ sky130_fd_sc_hd__a21o_2
X_10248_ _05118_ net798 _05117_ vssd1 vssd1 vccd1 vccd1 _00014_ sky130_fd_sc_hd__and3b_1
X_13036_ clknet_leaf_46_clk _00267_ net1203 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[24\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1130 net1131 vssd1 vssd1 vccd1 vccd1 net1130 sky130_fd_sc_hd__clkbuf_4
Xfanout1141 net1150 vssd1 vssd1 vccd1 vccd1 net1141 sky130_fd_sc_hd__buf_2
XANTENNA__12440__S net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1152 net1153 vssd1 vssd1 vccd1 vccd1 net1152 sky130_fd_sc_hd__buf_2
X_10179_ final_design.uart.BAUD_counter\[25\] final_design.uart.BAUD_counter\[24\]
+ final_design.uart.BAUD_counter\[27\] final_design.uart.BAUD_counter\[26\] vssd1
+ vssd1 vccd1 vccd1 _05069_ sky130_fd_sc_hd__or4_1
XANTENNA__10361__B1 net1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1163 net1165 vssd1 vssd1 vccd1 vccd1 net1163 sky130_fd_sc_hd__clkbuf_4
Xfanout1174 net1175 vssd1 vssd1 vccd1 vccd1 net1174 sky130_fd_sc_hd__clkbuf_4
Xfanout1185 net1186 vssd1 vssd1 vccd1 vccd1 net1185 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07534__S net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11564__B net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14003__CLK clknet_leaf_40_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1196 net1197 vssd1 vssd1 vccd1 vccd1 net1196 sky130_fd_sc_hd__buf_2
X_13938_ clknet_leaf_44_clk _01169_ net1209 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[926\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11861__B1 net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13869_ clknet_leaf_39_clk _01100_ net1205 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[857\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14153__CLK clknet_leaf_18_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06410_ final_design.CPU_instr_adr\[12\] vssd1 vssd1 vccd1 vccd1 _01365_ sky130_fd_sc_hd__inv_2
XANTENNA__11580__A net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07390_ final_design.cpu.reg_window\[130\] final_design.cpu.reg_window\[162\] net918
+ vssd1 vssd1 vccd1 vccd1 _02341_ sky130_fd_sc_hd__mux2_1
XANTENNA__06674__A net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12405__A2 net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10416__B2 net245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1833 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09282__A1 net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09060_ _03987_ vssd1 vssd1 vccd1 vccd1 _03988_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_13_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_1877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09985__A net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08011_ _01939_ net603 vssd1 vssd1 vccd1 vccd1 _02962_ sky130_fd_sc_hd__nand2_1
XFILLER_0_25_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12615__S _05080_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold602 final_design.cpu.reg_window\[446\] vssd1 vssd1 vccd1 vccd1 net1944 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold613 final_design.cpu.reg_window\[645\] vssd1 vssd1 vccd1 vccd1 net1955 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold624 final_design.cpu.reg_window\[458\] vssd1 vssd1 vccd1 vccd1 net1966 sky130_fd_sc_hd__dlygate4sd3_1
Xhold635 final_design.cpu.reg_window\[669\] vssd1 vssd1 vccd1 vccd1 net1977 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkload33_A clknet_leaf_42_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold646 final_design.cpu.reg_window\[545\] vssd1 vssd1 vccd1 vccd1 net1988 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_70_2605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold657 final_design.cpu.reg_window\[137\] vssd1 vssd1 vccd1 vccd1 net1999 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold668 final_design.cpu.reg_window\[450\] vssd1 vssd1 vccd1 vccd1 net2010 sky130_fd_sc_hd__dlygate4sd3_1
X_09962_ net90 _04880_ vssd1 vssd1 vccd1 vccd1 _04881_ sky130_fd_sc_hd__xnor2_1
Xhold679 final_design.cpu.reg_window\[483\] vssd1 vssd1 vccd1 vccd1 net2021 sky130_fd_sc_hd__dlygate4sd3_1
X_14197__1255 vssd1 vssd1 vccd1 vccd1 _14197__1255/HI net1255 sky130_fd_sc_hd__conb_1
X_08913_ _03768_ _03770_ vssd1 vssd1 vccd1 vccd1 _03857_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12895__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09893_ _03558_ _03559_ _03638_ vssd1 vssd1 vccd1 vccd1 _04812_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_40_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout296_A net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09742__C1 net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08844_ final_design.CPU_instr_adr\[20\] _03794_ vssd1 vssd1 vccd1 vccd1 _03795_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_58_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10352__B1 _05170_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_2512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1003_A _05173_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_68_2523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_2534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_2545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08775_ final_design.CPU_instr_adr\[8\] _02186_ vssd1 vssd1 vccd1 vccd1 _03726_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout463_A net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_64_2409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07726_ final_design.cpu.reg_window\[474\] final_design.cpu.reg_window\[506\] net863
+ vssd1 vssd1 vccd1 vccd1 _02677_ sky130_fd_sc_hd__mux2_1
XANTENNA_hold1209_A net166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout251_X net251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11852__B1 net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout630_A net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07657_ _02605_ _02607_ vssd1 vssd1 vccd1 vccd1 _02608_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout349_X net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout728_A net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06608_ net754 _01558_ vssd1 vssd1 vccd1 vccd1 _01559_ sky130_fd_sc_hd__or2_1
X_07588_ net712 _02538_ net877 vssd1 vssd1 vccd1 vccd1 _02539_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_76_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_1799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13520__CLK clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06539_ _01464_ _01475_ _01483_ vssd1 vssd1 vccd1 vccd1 _01490_ sky130_fd_sc_hd__nor3_1
XANTENNA__10407__B2 net246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09327_ _02641_ _03607_ _04051_ vssd1 vssd1 vccd1 vccd1 _04246_ sky130_fd_sc_hd__or3_1
XANTENNA__08076__A2 _03022_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout516_X net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09258_ net727 _04127_ _04176_ vssd1 vssd1 vccd1 vccd1 _04177_ sky130_fd_sc_hd__or3_2
XFILLER_0_65_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08209_ net874 _03141_ _03147_ _03153_ _03159_ vssd1 vssd1 vccd1 vccd1 _03160_ sky130_fd_sc_hd__o32a_4
X_09189_ net485 _04054_ vssd1 vssd1 vccd1 vccd1 _04108_ sky130_fd_sc_hd__nand2_1
XANTENNA__13670__CLK clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11220_ net645 _05925_ _05924_ net653 vssd1 vssd1 vccd1 vccd1 _05926_ sky130_fd_sc_hd__a211o_1
XFILLER_0_82_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11649__B net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout885_X net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11151_ net648 net228 vssd1 vssd1 vccd1 vccd1 _05865_ sky130_fd_sc_hd__and2_1
XANTENNA__07682__S1 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10102_ final_design.VGA_data_control.v_count\[0\] _05017_ _05007_ vssd1 vssd1 vccd1
+ vccd1 _05018_ sky130_fd_sc_hd__a21boi_1
X_11082_ _05780_ _05802_ _05803_ vssd1 vssd1 vccd1 vccd1 _05804_ sky130_fd_sc_hd__nor3_1
XANTENNA__14026__CLK clknet_leaf_60_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10033_ _04330_ _04951_ net448 vssd1 vssd1 vccd1 vccd1 _04952_ sky130_fd_sc_hd__a21oi_1
XANTENNA__06759__A net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input24_A DAT_I[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13050__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14176__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11984_ _06186_ net291 net407 net1587 vssd1 vssd1 vccd1 vccd1 _00717_ sky130_fd_sc_hd__a22o_1
XFILLER_0_59_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13723_ clknet_leaf_66_clk _00954_ net1063 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[711\]
+ sky130_fd_sc_hd__dfrtp_1
X_10935_ _05662_ _05663_ vssd1 vssd1 vccd1 vccd1 _05664_ sky130_fd_sc_hd__nor2_1
X_13654_ clknet_leaf_61_clk _00885_ net1137 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[642\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08185__S net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10866_ final_design.CPU_instr_adr\[20\] net1000 _05595_ net1042 vssd1 vssd1 vccd1
+ vccd1 _05598_ sky130_fd_sc_hd__o22a_1
XANTENNA__06494__A net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_34_clk_X clknet_leaf_34_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12605_ net1407 net996 net982 final_design.data_from_mem\[23\] vssd1 vssd1 vccd1
+ vccd1 _01298_ sky130_fd_sc_hd__a22o_1
XFILLER_0_13_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13585_ clknet_leaf_34_clk _00816_ net1239 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[573\]
+ sky130_fd_sc_hd__dfrtp_1
X_10797_ _05512_ _05514_ _05531_ vssd1 vssd1 vccd1 vccd1 _05532_ sky130_fd_sc_hd__and3_1
XFILLER_0_53_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_1817 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12536_ _06199_ net348 net323 net2152 vssd1 vssd1 vccd1 vccd1 _01240_ sky130_fd_sc_hd__a22o_1
XFILLER_0_82_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07814__A2 _02763_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_49_clk_X clknet_leaf_49_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12467_ _06127_ net349 net331 net2111 vssd1 vssd1 vccd1 vccd1 _01173_ sky130_fd_sc_hd__a22o_1
XANTENNA__12435__S net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14206_ net1264 vssd1 vssd1 vccd1 vccd1 gpio_oeb[18] sky130_fd_sc_hd__buf_2
XFILLER_0_1_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09567__A2 net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11418_ net1760 net220 net310 vssd1 vssd1 vccd1 vccd1 _00315_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12020__B1 net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12398_ _06096_ net349 net339 net2165 vssd1 vssd1 vccd1 vccd1 _01108_ sky130_fd_sc_hd__a22o_1
X_14137_ clknet_leaf_17_clk final_design.vga.h_next_count\[6\] net1114 vssd1 vssd1
+ vccd1 vccd1 final_design.VGA_data_control.VGA_request_address\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_10_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11349_ net436 net583 _06039_ net316 net1976 vssd1 vssd1 vccd1 vccd1 _00299_ sky130_fd_sc_hd__a32o_1
XFILLER_0_39_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1883 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14068_ clknet_leaf_15_clk _00038_ net1094 vssd1 vssd1 vccd1 vccd1 final_design.uart.BAUD_counter_state
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_78_1913 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13019_ clknet_leaf_0_clk _00250_ net1061 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12170__S net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06890_ final_design.cpu.reg_window\[915\] final_design.cpu.reg_window\[947\] net911
+ vssd1 vssd1 vccd1 vccd1 _01841_ sky130_fd_sc_hd__mux2_1
XANTENNA__10334__B1 net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12087__B1 net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08560_ _03507_ _03508_ _03509_ _03510_ net679 net692 vssd1 vssd1 vccd1 vccd1 _03511_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__07189__S0 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10637__A1 net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13543__CLK clknet_leaf_62_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07511_ _01824_ _02461_ vssd1 vssd1 vccd1 vccd1 _02462_ sky130_fd_sc_hd__nand2_1
XANTENNA__10637__B2 net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08491_ final_design.cpu.reg_window\[899\] final_design.cpu.reg_window\[931\] net823
+ vssd1 vssd1 vccd1 vccd1 _03442_ sky130_fd_sc_hd__mux2_1
XANTENNA__06675__Y _01626_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11514__S net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07442_ net740 _02392_ vssd1 vssd1 vccd1 vccd1 _02393_ sky130_fd_sc_hd__nand2_1
XFILLER_0_58_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09986__Y _04905_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07373_ net758 _02323_ vssd1 vssd1 vccd1 vccd1 _02324_ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_21_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13693__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09112_ _03715_ _04031_ vssd1 vssd1 vccd1 vccd1 _04032_ sky130_fd_sc_hd__nor2_1
XFILLER_0_44_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_2803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11601__A3 _06156_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_2814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09043_ _02444_ net622 _03969_ _03972_ vssd1 vssd1 vccd1 vccd1 _03973_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout309_A _06095_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold410 final_design.cpu.reg_window\[664\] vssd1 vssd1 vccd1 vccd1 net1752 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12011__B1 net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14049__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold421 final_design.cpu.reg_window\[657\] vssd1 vssd1 vccd1 vccd1 net1763 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold432 final_design.cpu.reg_window\[705\] vssd1 vssd1 vccd1 vccd1 net1774 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_1794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11365__A2 net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold443 final_design.cpu.reg_window\[727\] vssd1 vssd1 vccd1 vccd1 net1785 sky130_fd_sc_hd__dlygate4sd3_1
Xhold454 net135 vssd1 vssd1 vccd1 vccd1 net1796 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1120_A net1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold465 final_design.cpu.reg_window\[656\] vssd1 vssd1 vccd1 vccd1 net1807 sky130_fd_sc_hd__dlygate4sd3_1
Xhold476 final_design.cpu.reg_window\[766\] vssd1 vssd1 vccd1 vccd1 net1818 sky130_fd_sc_hd__dlygate4sd3_1
Xhold487 final_design.cpu.reg_window\[562\] vssd1 vssd1 vccd1 vccd1 net1829 sky130_fd_sc_hd__dlygate4sd3_1
Xhold498 final_design.cpu.reg_window\[90\] vssd1 vssd1 vccd1 vccd1 net1840 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout901 net905 vssd1 vssd1 vccd1 vccd1 net901 sky130_fd_sc_hd__clkbuf_4
X_09945_ net725 _04863_ vssd1 vssd1 vccd1 vccd1 _04864_ sky130_fd_sc_hd__nor2_1
Xfanout912 net917 vssd1 vssd1 vccd1 vccd1 net912 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_5_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout923 net927 vssd1 vssd1 vccd1 vccd1 net923 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_42_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout580_A net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout934 net952 vssd1 vssd1 vccd1 vccd1 net934 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08518__B1 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout945 net952 vssd1 vssd1 vccd1 vccd1 net945 sky130_fd_sc_hd__buf_2
XANTENNA_fanout299_X net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout678_A net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13073__CLK clknet_leaf_34_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout956 net957 vssd1 vssd1 vccd1 vccd1 net956 sky130_fd_sc_hd__clkbuf_4
Xfanout967 _04035_ vssd1 vssd1 vccd1 vccd1 net967 sky130_fd_sc_hd__clkbuf_4
X_09876_ net534 net533 net532 net530 net452 net460 vssd1 vssd1 vccd1 vccd1 _04795_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout1006_X net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout978 net981 vssd1 vssd1 vccd1 vccd1 net978 sky130_fd_sc_hd__clkbuf_4
Xhold1110 final_design.cpu.reg_window\[831\] vssd1 vssd1 vccd1 vccd1 net2452 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout989 _05167_ vssd1 vssd1 vccd1 vccd1 net989 sky130_fd_sc_hd__clkbuf_2
Xhold1121 net156 vssd1 vssd1 vccd1 vccd1 net2463 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1132 final_design.cpu.reg_window\[105\] vssd1 vssd1 vccd1 vccd1 net2474 sky130_fd_sc_hd__dlygate4sd3_1
X_08827_ _01358_ _01538_ _03777_ vssd1 vssd1 vccd1 vccd1 _03778_ sky130_fd_sc_hd__a21oi_1
Xhold1143 final_design.cpu.reg_window\[417\] vssd1 vssd1 vccd1 vccd1 net2485 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout845_A net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1154 final_design.cpu.reg_window\[419\] vssd1 vssd1 vccd1 vccd1 net2496 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout466_X net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1165 final_design.cpu.reg_window\[395\] vssd1 vssd1 vccd1 vccd1 net2507 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1176 final_design.uart.BAUD_counter\[4\] vssd1 vssd1 vccd1 vccd1 net2518 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12078__B1 net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1187 _01310_ vssd1 vssd1 vccd1 vccd1 net2529 sky130_fd_sc_hd__dlygate4sd3_1
X_08758_ final_design.CPU_instr_adr\[3\] _02330_ vssd1 vssd1 vccd1 vccd1 _03709_ sky130_fd_sc_hd__and2_1
Xhold1198 net143 vssd1 vssd1 vccd1 vccd1 net2540 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11825__A0 net207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07709_ _02656_ _02657_ _02658_ _02659_ net686 net704 vssd1 vssd1 vccd1 vccd1 _02660_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout633_X net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08689_ net608 _03549_ _03523_ _02419_ vssd1 vssd1 vccd1 vccd1 _03640_ sky130_fd_sc_hd__a211o_1
XANTENNA__06927__S0 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12093__A3 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11424__S net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10720_ _05438_ _05441_ _05457_ _05436_ vssd1 vssd1 vccd1 vccd1 _05459_ sky130_fd_sc_hd__a211o_1
XANTENNA__12910__CLK clknet_leaf_61_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07203__A net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10651_ _05391_ _05392_ vssd1 vssd1 vccd1 vccd1 _05393_ sky130_fd_sc_hd__nand2_1
XANTENNA__09246__A1 _04158_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10582_ _05309_ _05326_ vssd1 vssd1 vccd1 vccd1 _05328_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12250__B1 net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13370_ clknet_leaf_58_clk _00601_ net1125 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[358\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09797__A2 net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12321_ net1673 net191 net367 vssd1 vssd1 vccd1 vccd1 _01035_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_40_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12252_ net580 _06181_ net511 net374 net1642 vssd1 vssd1 vccd1 vccd1 _00968_ sky130_fd_sc_hd__a32o_1
XANTENNA__12002__B1 net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11379__B net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10013__C1 net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11203_ net646 net243 vssd1 vssd1 vccd1 vccd1 _05911_ sky130_fd_sc_hd__and2_1
XANTENNA__09954__C1 net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12183_ net1769 net200 net380 vssd1 vssd1 vccd1 vccd1 _00902_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_1747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_61_clk_A clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13416__CLK clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08969__A net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11134_ net803 net805 _02359_ vssd1 vssd1 vccd1 vccd1 _05849_ sky130_fd_sc_hd__and3b_2
XANTENNA__12305__A1 net221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11065_ _01358_ _03821_ net1060 vssd1 vssd1 vccd1 vccd1 _05788_ sky130_fd_sc_hd__mux2_1
XANTENNA__10316__B1 net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10016_ net263 _04928_ _04934_ vssd1 vssd1 vccd1 vccd1 _04935_ sky130_fd_sc_hd__and3_1
XANTENNA__10867__A1 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input27_X net27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13566__CLK clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10867__B2 net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_3007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_3018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_3029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12069__B1 net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14146__RESET_B net1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12608__A2 net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11816__A0 net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11967_ _06169_ net276 net404 net1794 vssd1 vssd1 vccd1 vccd1 _00700_ sky130_fd_sc_hd__a22o_1
XANTENNA__09485__A1 _02502_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13706_ clknet_leaf_60_clk _00937_ net1141 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[694\]
+ sky130_fd_sc_hd__dfrtp_1
X_10918_ _05624_ _05645_ _05646_ net1005 vssd1 vssd1 vccd1 vccd1 _05648_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_15_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11898_ net209 net2237 net274 vssd1 vssd1 vccd1 vccd1 _00640_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_28_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10458__B net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_15_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_28_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13637_ clknet_leaf_50_clk _00868_ net1181 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[625\]
+ sky130_fd_sc_hd__dfrtp_1
X_14196__1254 vssd1 vssd1 vccd1 vccd1 _14196__1254/HI net1254 sky130_fd_sc_hd__conb_1
X_10849_ _05559_ _05564_ _05581_ vssd1 vssd1 vccd1 vccd1 _05582_ sky130_fd_sc_hd__or3_1
XFILLER_0_67_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12796__27 clknet_leaf_31_clk vssd1 vssd1 vccd1 vccd1 net1337 sky130_fd_sc_hd__inv_2
XANTENNA__07248__B1 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11044__B2 net1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_14_clk_A clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12241__B1 net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13568_ clknet_leaf_11_clk _00799_ net1087 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[556\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13781__RESET_B net1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11595__A2 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12519_ _06181_ net354 net328 net1959 vssd1 vssd1 vccd1 vccd1 _01224_ sky130_fd_sc_hd__a22o_1
XANTENNA__10474__A net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12165__S net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13499_ clknet_leaf_0_clk _00730_ net1071 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[487\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07259__S net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06471__A1 final_design.data_from_mem\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_29_clk_A clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13096__CLK clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08212__A2 _03160_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout208 _05965_ vssd1 vssd1 vccd1 vccd1 net208 sky130_fd_sc_hd__buf_2
Xfanout219 _05928_ vssd1 vssd1 vccd1 vccd1 net219 sky130_fd_sc_hd__clkbuf_2
X_07991_ _02938_ _02939_ _02940_ _02941_ net682 net702 vssd1 vssd1 vccd1 vccd1 _02942_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__13909__CLK clknet_leaf_57_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11509__S net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09730_ net495 _04113_ _04268_ vssd1 vssd1 vccd1 vccd1 _04649_ sky130_fd_sc_hd__or3_1
X_06942_ final_design.cpu.reg_window\[145\] final_design.cpu.reg_window\[177\] net928
+ vssd1 vssd1 vccd1 vccd1 _01893_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_1721 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09661_ net487 _04225_ vssd1 vssd1 vccd1 vccd1 _04580_ sky130_fd_sc_hd__nor2_1
XFILLER_0_78_1765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06873_ net549 _01823_ vssd1 vssd1 vccd1 vccd1 _01824_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_39_1727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_1618 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08612_ net529 net497 vssd1 vssd1 vccd1 vccd1 _03563_ sky130_fd_sc_hd__nor2_1
XANTENNA__12933__CLK clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09592_ net729 _04502_ _04508_ _04482_ vssd1 vssd1 vccd1 vccd1 _04511_ sky130_fd_sc_hd__a31o_1
XFILLER_0_55_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08543_ final_design.cpu.reg_window\[65\] final_design.cpu.reg_window\[97\] net836
+ vssd1 vssd1 vccd1 vccd1 _03494_ sky130_fd_sc_hd__mux2_1
XANTENNA__11807__B1 net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12075__A3 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11283__A1 net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12480__B1 net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08474_ _03387_ _03389_ _03420_ _03422_ vssd1 vssd1 vccd1 vccd1 _03425_ sky130_fd_sc_hd__o22a_1
XFILLER_0_65_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07425_ net752 _02369_ net746 vssd1 vssd1 vccd1 vccd1 _02376_ sky130_fd_sc_hd__o21a_1
XFILLER_0_15_1771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout426_A net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1168_A net1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12232__B1 net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07356_ final_design.cpu.reg_window\[3\] final_design.cpu.reg_window\[35\] net905
+ vssd1 vssd1 vccd1 vccd1 _02307_ sky130_fd_sc_hd__mux2_1
X_07287_ _02232_ _02237_ net751 vssd1 vssd1 vccd1 vccd1 _02238_ sky130_fd_sc_hd__mux2_1
XANTENNA__13439__CLK clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10384__A net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07169__S net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09026_ net259 _03957_ net1013 vssd1 vssd1 vccd1 vccd1 _03958_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout795_A _01418_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold240 final_design.cpu.reg_window\[965\] vssd1 vssd1 vccd1 vccd1 net1582 sky130_fd_sc_hd__dlygate4sd3_1
Xhold251 final_design.cpu.reg_window\[974\] vssd1 vssd1 vccd1 vccd1 net1593 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09400__A1 net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07637__S1 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold262 final_design.cpu.reg_window\[158\] vssd1 vssd1 vccd1 vccd1 net1604 sky130_fd_sc_hd__dlygate4sd3_1
Xhold273 final_design.cpu.reg_window\[749\] vssd1 vssd1 vccd1 vccd1 net1615 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold284 final_design.cpu.reg_window\[561\] vssd1 vssd1 vccd1 vccd1 net1626 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13589__CLK clknet_leaf_58_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold295 final_design.cpu.reg_window\[514\] vssd1 vssd1 vccd1 vccd1 net1637 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout962_A _04036_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout583_X net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout720 net721 vssd1 vssd1 vccd1 vccd1 net720 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11419__S net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout731 net732 vssd1 vssd1 vccd1 vccd1 net731 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_61_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09928_ _04843_ _04845_ net725 _04831_ vssd1 vssd1 vccd1 vccd1 _04847_ sky130_fd_sc_hd__a211o_1
Xfanout742 net743 vssd1 vssd1 vccd1 vccd1 net742 sky130_fd_sc_hd__clkbuf_4
Xfanout753 net755 vssd1 vssd1 vccd1 vccd1 net753 sky130_fd_sc_hd__clkbuf_4
Xfanout764 net766 vssd1 vssd1 vccd1 vccd1 net764 sky130_fd_sc_hd__buf_4
Xfanout775 net777 vssd1 vssd1 vccd1 vccd1 net775 sky130_fd_sc_hd__buf_4
XFILLER_0_77_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout786 net788 vssd1 vssd1 vccd1 vccd1 net786 sky130_fd_sc_hd__clkbuf_4
Xfanout797 net798 vssd1 vssd1 vccd1 vccd1 net797 sky130_fd_sc_hd__clkbuf_2
X_09859_ net538 net537 net535 net534 net452 net461 vssd1 vssd1 vccd1 vccd1 _04778_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout750_X net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12870_ clknet_leaf_20_clk _00108_ net1158 vssd1 vssd1 vccd1 vccd1 final_design.data_from_mem\[4\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_38_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11821_ net217 net2060 net264 vssd1 vssd1 vccd1 vccd1 _00573_ sky130_fd_sc_hd__mux2_1
XANTENNA__12066__A3 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11274__A1 net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11752_ net223 net2242 net418 vssd1 vssd1 vccd1 vccd1 _00515_ sky130_fd_sc_hd__mux2_1
XANTENNA__12471__B1 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09700__X _04619_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10703_ _05438_ _05441_ vssd1 vssd1 vccd1 vccd1 _05443_ sky130_fd_sc_hd__or2_1
X_11683_ net238 net626 vssd1 vssd1 vccd1 vccd1 _06200_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_46_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input91_A memory_size[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1901 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13422_ clknet_leaf_42_clk _00653_ net1222 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[410\]
+ sky130_fd_sc_hd__dfrtp_1
X_10634_ _05351_ _05376_ _05371_ vssd1 vssd1 vccd1 vccd1 _05377_ sky130_fd_sc_hd__o21a_1
XFILLER_0_10_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12223__B1 net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09314__S1 net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08463__S net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_42_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06772__A _01718_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11577__A2 net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08978__B1 net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13353_ clknet_leaf_36_clk _00584_ net1230 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[341\]
+ sky130_fd_sc_hd__dfrtp_1
X_10565_ net96 final_design.VGA_adr\[4\] vssd1 vssd1 vccd1 vccd1 _05311_ sky130_fd_sc_hd__nand2_1
XFILLER_0_23_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12304_ net1802 net244 net364 vssd1 vssd1 vccd1 vccd1 _01018_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07650__B1 net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13284_ clknet_leaf_52_clk _00515_ net1174 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[272\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_62_1500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10496_ _05244_ _05245_ vssd1 vssd1 vccd1 vccd1 _05246_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_66_1680 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11329__A2 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12235_ net569 _06165_ net507 net373 net1583 vssd1 vssd1 vccd1 vccd1 _00952_ sky130_fd_sc_hd__a32o_1
XFILLER_0_62_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_36_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09147__X _04066_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11396__Y _06081_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12166_ net1872 net241 net381 vssd1 vssd1 vccd1 vccd1 _00885_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_36_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11117_ final_design.uart.bits_received\[2\] _05830_ _05831_ _05834_ vssd1 vssd1
+ vccd1 vccd1 _00207_ sky130_fd_sc_hd__a22o_1
XANTENNA__12956__CLK clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12097_ net1624 net241 net389 vssd1 vssd1 vccd1 vccd1 _00821_ sky130_fd_sc_hd__mux2_1
XANTENNA__12799__30_A clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11048_ net670 _05758_ _05771_ vssd1 vssd1 vccd1 vccd1 _05772_ sky130_fd_sc_hd__o21ai_1
Xinput8 DAT_I[15] vssd1 vssd1 vccd1 vccd1 net8 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_56_1304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11572__B net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12999_ net1330 _00230_ net1196 vssd1 vssd1 vccd1 vccd1 final_design.CPU_instr_adr\[19\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_73_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10068__A2 net251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09610__X _04529_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08681__A2 _03610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07210_ final_design.cpu.reg_window\[264\] final_design.cpu.reg_window\[296\] net901
+ vssd1 vssd1 vccd1 vccd1 _02161_ sky130_fd_sc_hd__mux2_1
XANTENNA__12214__B1 net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08190_ net708 _03140_ vssd1 vssd1 vccd1 vccd1 _03141_ sky130_fd_sc_hd__nor2_1
XFILLER_0_43_902 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07141_ _01488_ net728 _01820_ vssd1 vssd1 vccd1 vccd1 _02092_ sky130_fd_sc_hd__or3b_1
XFILLER_0_43_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07072_ final_design.cpu.reg_window\[909\] final_design.cpu.reg_window\[941\] net934
+ vssd1 vssd1 vccd1 vccd1 _02023_ sky130_fd_sc_hd__mux2_1
XANTENNA__09993__A net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13731__CLK clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10932__A net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06621__S net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08292__S1 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07974_ final_design.cpu.reg_window\[593\] final_design.cpu.reg_window\[625\] net845
+ vssd1 vssd1 vccd1 vccd1 _02925_ sky130_fd_sc_hd__mux2_1
XANTENNA__13881__CLK clknet_leaf_55_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09713_ net727 _04631_ vssd1 vssd1 vccd1 vccd1 _04632_ sky130_fd_sc_hd__or2_1
XANTENNA__07018__A net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06925_ final_design.cpu.reg_window\[594\] final_design.cpu.reg_window\[626\] net924
+ vssd1 vssd1 vccd1 vccd1 _01876_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout376_A net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09504__Y _04423_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09644_ _04342_ _04561_ _04562_ _04222_ vssd1 vssd1 vccd1 vccd1 _04563_ sky130_fd_sc_hd__o211a_1
XANTENNA__09792__S1 net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06856_ _01803_ _01804_ _01805_ _01806_ net776 net794 vssd1 vssd1 vccd1 vccd1 _01807_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__06857__A net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13111__CLK clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12578__B net35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09575_ net261 _04484_ _04493_ vssd1 vssd1 vccd1 vccd1 _04494_ sky130_fd_sc_hd__and3_1
XFILLER_0_77_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06787_ final_design.cpu.reg_window\[598\] final_design.cpu.reg_window\[630\] net920
+ vssd1 vssd1 vccd1 vccd1 _01738_ sky130_fd_sc_hd__mux2_1
X_08526_ final_design.cpu.reg_window\[578\] final_design.cpu.reg_window\[610\] net832
+ vssd1 vssd1 vccd1 vccd1 _03477_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08657__C1 _01453_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08457_ _03404_ _03405_ _03406_ _03407_ net677 net701 vssd1 vssd1 vccd1 vccd1 _03408_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout710_A net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout331_X net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13261__CLK clknet_leaf_48_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1410 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout429_X net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13632__RESET_B net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07408_ final_design.data_from_mem\[9\] net970 _02357_ vssd1 vssd1 vccd1 vccd1 _02359_
+ sky130_fd_sc_hd__o21ai_4
XANTENNA__12205__B1 net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08388_ net716 _03338_ vssd1 vssd1 vccd1 vccd1 _03339_ sky130_fd_sc_hd__nor2_1
X_07339_ final_design.cpu.reg_window\[580\] final_design.cpu.reg_window\[612\] net900
+ vssd1 vssd1 vccd1 vccd1 _02290_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_754 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10350_ wb_manage.BUSY_O net1026 wb_manage.prev_BUSY_O vssd1 vssd1 vccd1 vccd1 _05171_
+ sky130_fd_sc_hd__or3b_1
X_09009_ net255 _03940_ _03941_ _03942_ net1017 vssd1 vssd1 vccd1 vccd1 _03943_ sky130_fd_sc_hd__a221o_1
XFILLER_0_42_990 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10281_ final_design.uart.BAUD_counter\[30\] _05138_ vssd1 vssd1 vccd1 vccd1 _05139_
+ sky130_fd_sc_hd__and2_1
XANTENNA__10842__A net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12979__CLK clknet_leaf_25_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09385__A0 net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_3_0_clk_X clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12020_ _06222_ net288 net402 net2387 vssd1 vssd1 vccd1 vccd1 _00751_ sky130_fd_sc_hd__a22o_1
XANTENNA__11657__B net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09127__B _04045_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14195__1253 vssd1 vssd1 vccd1 vccd1 _14195__1253/HI net1253 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_50_1924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout550 _01784_ vssd1 vssd1 vccd1 vccd1 net550 sky130_fd_sc_hd__buf_2
Xfanout561 net562 vssd1 vssd1 vccd1 vccd1 net561 sky130_fd_sc_hd__buf_2
Xfanout572 net573 vssd1 vssd1 vccd1 vccd1 net572 sky130_fd_sc_hd__clkbuf_4
Xfanout583 net587 vssd1 vssd1 vccd1 vccd1 net583 sky130_fd_sc_hd__clkbuf_2
X_13971_ clknet_leaf_40_clk _01202_ net1219 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[959\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout594 _03627_ vssd1 vssd1 vccd1 vccd1 net594 sky130_fd_sc_hd__buf_4
XANTENNA__11673__A net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12922_ clknet_leaf_61_clk _00160_ net1137 vssd1 vssd1 vccd1 vccd1 net144 sky130_fd_sc_hd__dfrtp_1
XANTENNA__12692__B1 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07362__S net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_1619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_17_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12853_ clknet_leaf_14_clk _00091_ net1110 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.ready_data\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_48_1842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11804_ net2391 net415 net291 _06053_ vssd1 vssd1 vccd1 vccd1 _00557_ sky130_fd_sc_hd__a22o_1
XANTENNA__13604__CLK clknet_leaf_54_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08405__A_N _02239_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1857 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11798__A2 net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11735_ net804 _05846_ _05867_ vssd1 vssd1 vccd1 vccd1 _06226_ sky130_fd_sc_hd__or3_1
XFILLER_0_12_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08663__A2 _02061_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11666_ net434 net577 _06190_ net300 net1493 vssd1 vssd1 vccd1 vccd1 _00465_ sky130_fd_sc_hd__a32o_1
XANTENNA__12774__5_A clknet_leaf_25_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13405_ clknet_leaf_5_clk _00636_ net1077 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[393\]
+ sky130_fd_sc_hd__dfrtp_1
X_10617_ net668 _05348_ _05360_ net964 _05359_ vssd1 vssd1 vccd1 vccd1 _05361_ sky130_fd_sc_hd__o221a_1
XANTENNA__12211__A3 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11597_ net437 net584 _06154_ net304 net2130 vssd1 vssd1 vccd1 vccd1 _00432_ sky130_fd_sc_hd__a32o_1
XFILLER_0_3_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13336_ clknet_leaf_63_clk _00567_ net1121 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[324\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10548_ _05293_ _05294_ vssd1 vssd1 vccd1 vccd1 _05295_ sky130_fd_sc_hd__or2_1
XANTENNA__11970__A2 net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13267_ clknet_leaf_40_clk _00498_ net1207 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[255\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12443__S net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10479_ net47 _05223_ _05225_ _05227_ vssd1 vssd1 vccd1 vccd1 _05230_ sky130_fd_sc_hd__nand4_1
XANTENNA__14224__A final_design.pixel_data vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11200__X _05908_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12218_ net580 _06146_ net511 net378 net2117 vssd1 vssd1 vccd1 vccd1 _00936_ sky130_fd_sc_hd__a32o_1
XFILLER_0_62_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13198_ clknet_leaf_45_clk _00429_ net1213 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[186\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11722__A2 net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12149_ net200 net2368 net384 vssd1 vssd1 vccd1 vccd1 _00870_ sky130_fd_sc_hd__mux2_1
XANTENNA__14161__RESET_B net1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13134__CLK clknet_leaf_45_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08026__S1 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12278__A3 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06710_ _01658_ _01660_ vssd1 vssd1 vccd1 vccd1 _01661_ sky130_fd_sc_hd__nor2_1
XFILLER_0_75_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07690_ _02640_ vssd1 vssd1 vccd1 vccd1 _02641_ sky130_fd_sc_hd__inv_2
X_06641_ final_design.cpu.reg_window\[603\] final_design.cpu.reg_window\[635\] net941
+ vssd1 vssd1 vccd1 vccd1 _01592_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13284__CLK clknet_leaf_52_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06901__A2 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09360_ _04056_ _04278_ _04274_ net261 vssd1 vssd1 vccd1 vccd1 _04279_ sky130_fd_sc_hd__o211ai_2
X_06572_ final_design.cpu.reg_window\[861\] final_design.cpu.reg_window\[893\] net949
+ vssd1 vssd1 vccd1 vccd1 _01523_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11789__A2 net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08311_ _03259_ _03260_ vssd1 vssd1 vccd1 vccd1 _03262_ sky130_fd_sc_hd__nor2_2
XFILLER_0_75_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09291_ _01626_ _01657_ net459 vssd1 vssd1 vccd1 vccd1 _04210_ sky130_fd_sc_hd__mux2_1
XANTENNA__12618__S _05080_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_2242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11522__S net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_2253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_1506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_1717 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_13 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08242_ _02097_ net611 vssd1 vssd1 vccd1 vccd1 _03193_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_60_2264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10461__A2 net1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_24 _06257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10646__B net250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08173_ final_design.cpu.reg_window\[655\] final_design.cpu.reg_window\[687\] net806
+ vssd1 vssd1 vccd1 vccd1 _03124_ sky130_fd_sc_hd__mux2_1
XANTENNA__08406__A2 _03352_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12202__A3 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07124_ final_design.cpu.reg_window\[203\] final_design.cpu.reg_window\[235\] net915
+ vssd1 vssd1 vccd1 vccd1 _02075_ sky130_fd_sc_hd__mux2_1
XANTENNA__11410__A1 net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07055_ final_design.cpu.reg_window\[397\] final_design.cpu.reg_window\[429\] net934
+ vssd1 vssd1 vccd1 vccd1 _02006_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11961__A2 net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_2182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput120 net120 vssd1 vssd1 vccd1 vccd1 ADR_O[27] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_2_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_2193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput131 net131 vssd1 vssd1 vccd1 vccd1 ADR_O[8] sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout1033_A net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12780__11 clknet_leaf_28_clk vssd1 vssd1 vccd1 vccd1 net1321 sky130_fd_sc_hd__inv_2
Xoutput142 net142 vssd1 vssd1 vccd1 vccd1 DAT_O[17] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_54_2046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_2057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput153 net153 vssd1 vssd1 vccd1 vccd1 DAT_O[27] sky130_fd_sc_hd__buf_2
XFILLER_0_11_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08132__A net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput164 net164 vssd1 vssd1 vccd1 vccd1 DAT_O[8] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_54_2068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput175 net175 vssd1 vssd1 vccd1 vccd1 gpio_out[3] sky130_fd_sc_hd__buf_2
XANTENNA_fanout493_A _03453_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_1881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07957_ final_design.cpu.reg_window\[465\] final_design.cpu.reg_window\[497\] net848
+ vssd1 vssd1 vccd1 vccd1 _02908_ sky130_fd_sc_hd__mux2_1
XANTENNA__12269__A3 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout281_X net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout660_A _02512_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout758_A net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout379_X net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06908_ final_design.cpu.reg_window\[466\] final_design.cpu.reg_window\[498\] net924
+ vssd1 vssd1 vccd1 vccd1 _01859_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_1917 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07888_ _01722_ net606 vssd1 vssd1 vccd1 vccd1 _02839_ sky130_fd_sc_hd__nand2_1
X_09627_ _04046_ _04545_ _04543_ vssd1 vssd1 vccd1 vccd1 _04546_ sky130_fd_sc_hd__a21o_1
XFILLER_0_69_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06839_ _01785_ _01788_ vssd1 vssd1 vccd1 vccd1 _01790_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout546_X net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13813__RESET_B net1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09558_ _04452_ _04455_ _04476_ vssd1 vssd1 vccd1 vccd1 _04477_ sky130_fd_sc_hd__a21boi_1
XANTENNA__12426__B1 net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_1663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13777__CLK clknet_leaf_34_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08509_ final_design.cpu.reg_window\[450\] final_design.cpu.reg_window\[482\] net832
+ vssd1 vssd1 vccd1 vccd1 _03460_ sky130_fd_sc_hd__mux2_1
X_09489_ net484 _04407_ vssd1 vssd1 vccd1 vccd1 _04408_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout713_X net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11432__S net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11520_ net1743 net204 net523 vssd1 vssd1 vccd1 vccd1 _00388_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06751__S1 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11451_ net227 net2495 net307 vssd1 vssd1 vccd1 vccd1 _00342_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10402_ _03481_ _05181_ vssd1 vssd1 vccd1 vccd1 _05184_ sky130_fd_sc_hd__nor2_1
X_14170_ clknet_leaf_18_clk _01344_ net1114 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.data_to_VGA\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11401__A1 final_design.data_from_mem\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11382_ net435 net586 _06068_ net316 net2342 vssd1 vssd1 vccd1 vccd1 _00303_ sky130_fd_sc_hd__a32o_1
X_13121_ clknet_leaf_49_clk _00352_ net1184 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[109\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11952__A2 net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10333_ net1504 net1010 net987 final_design.data_from_mem\[18\] vssd1 vssd1 vccd1
+ vccd1 _00090_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13157__CLK clknet_leaf_49_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input54_A mem_adr_start[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13052_ clknet_leaf_3_clk _00283_ net1066 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[40\]
+ sky130_fd_sc_hd__dfrtp_1
X_10264_ _05128_ net797 _05127_ vssd1 vssd1 vccd1 vccd1 _00021_ sky130_fd_sc_hd__and3b_1
XANTENNA__11704__A2 net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12003_ _06205_ net284 net401 net2091 vssd1 vssd1 vccd1 vccd1 _00734_ sky130_fd_sc_hd__a22o_1
X_10195_ _05082_ _05083_ vssd1 vssd1 vccd1 vccd1 _05084_ sky130_fd_sc_hd__or2_1
XANTENNA__08008__S1 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout380 net381 vssd1 vssd1 vccd1 vccd1 net380 sky130_fd_sc_hd__buf_6
Xfanout391 _06265_ vssd1 vssd1 vccd1 vccd1 net391 sky130_fd_sc_hd__buf_6
X_13954_ clknet_leaf_4_clk _01185_ net1079 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[942\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_17_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08188__S net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12905_ clknet_leaf_60_clk _00143_ net1140 vssd1 vssd1 vccd1 vccd1 net156 sky130_fd_sc_hd__dfrtp_1
X_13885_ clknet_leaf_1_clk _01116_ net1081 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[873\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_1476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12836_ clknet_leaf_19_clk _00074_ net1156 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.ready_data\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12417__B1 net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_1042 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12767_ _01369_ _01398_ _06383_ _06398_ vssd1 vssd1 vccd1 vccd1 _06402_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__12438__S net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08636__A2 _02961_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06647__A1 final_design.data_from_mem\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10443__A2 net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11718_ net433 net574 _06217_ net297 net1783 vssd1 vssd1 vccd1 vccd1 _00490_ sky130_fd_sc_hd__a32o_1
X_12698_ _01368_ _06334_ _06336_ _06337_ vssd1 vssd1 vccd1 vccd1 _06339_ sky130_fd_sc_hd__o31a_2
XANTENNA__08217__A _02097_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput11 DAT_I[18] vssd1 vssd1 vccd1 vccd1 net11 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11649_ net194 net631 vssd1 vssd1 vccd1 vccd1 _06182_ sky130_fd_sc_hd__and2_1
Xinput22 DAT_I[28] vssd1 vssd1 vccd1 vccd1 net22 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_1761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput33 DAT_I[9] vssd1 vssd1 vccd1 vccd1 net33 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput44 mem_adr_start[17] vssd1 vssd1 vccd1 vccd1 net44 sky130_fd_sc_hd__buf_1
XFILLER_0_3_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput55 mem_adr_start[27] vssd1 vssd1 vccd1 vccd1 net55 sky130_fd_sc_hd__clkbuf_1
Xinput66 mem_adr_start[8] vssd1 vssd1 vccd1 vccd1 net66 sky130_fd_sc_hd__clkbuf_1
XANTENNA__06960__A _01908_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput77 memory_size[18] vssd1 vssd1 vccd1 vccd1 net77 sky130_fd_sc_hd__buf_1
Xhold806 final_design.cpu.reg_window\[1014\] vssd1 vssd1 vccd1 vccd1 net2148 sky130_fd_sc_hd__dlygate4sd3_1
Xhold817 final_design.cpu.reg_window\[447\] vssd1 vssd1 vccd1 vccd1 net2159 sky130_fd_sc_hd__dlygate4sd3_1
Xinput88 memory_size[28] vssd1 vssd1 vccd1 vccd1 net88 sky130_fd_sc_hd__buf_1
XANTENNA__10746__A3 net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13319_ clknet_leaf_59_clk _00550_ net1125 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[307\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11943__A2 net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11578__A net197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold828 final_design.cpu.reg_window\[469\] vssd1 vssd1 vccd1 vccd1 net2170 sky130_fd_sc_hd__dlygate4sd3_1
Xinput99 memory_size[9] vssd1 vssd1 vccd1 vccd1 net99 sky130_fd_sc_hd__buf_1
Xhold839 final_design.cpu.reg_window\[1010\] vssd1 vssd1 vccd1 vccd1 net2181 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12173__S net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1761 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09048__A net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14082__CLK clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11156__B1 net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_72_2680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08860_ final_design.CPU_instr_adr\[30\] _03801_ vssd1 vssd1 vccd1 vccd1 _03810_
+ sky130_fd_sc_hd__or2_1
XANTENNA__09990__B net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07811_ _02756_ _02761_ net713 vssd1 vssd1 vccd1 vccd1 _02762_ sky130_fd_sc_hd__mux2_1
X_08791_ _03683_ _03685_ _03686_ _03739_ vssd1 vssd1 vccd1 vccd1 _03742_ sky130_fd_sc_hd__and4_1
XANTENNA__11517__S net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07742_ final_design.cpu.reg_window\[666\] final_design.cpu.reg_window\[698\] net861
+ vssd1 vssd1 vccd1 vccd1 _02693_ sky130_fd_sc_hd__mux2_1
XANTENNA__08324__A1 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07673_ final_design.cpu.reg_window\[862\] final_design.cpu.reg_window\[894\] net856
+ vssd1 vssd1 vccd1 vccd1 _02624_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_66_2451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_66_2462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09412_ _02802_ _02834_ _04330_ _02900_ _02800_ vssd1 vssd1 vccd1 vccd1 _04331_ sky130_fd_sc_hd__a311o_1
XANTENNA__12408__B1 net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06624_ final_design.cpu.reg_window\[411\] final_design.cpu.reg_window\[443\] net948
+ vssd1 vssd1 vccd1 vccd1 _01575_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_62_2315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_2326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07730__S net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_62_2337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09343_ net472 _04098_ vssd1 vssd1 vccd1 vccd1 _04262_ sky130_fd_sc_hd__or2_2
X_06555_ net744 _01505_ vssd1 vssd1 vccd1 vccd1 _01506_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout241_A net242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout339_A net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1284 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_507 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09274_ net85 _04192_ vssd1 vssd1 vccd1 vccd1 _04193_ sky130_fd_sc_hd__or2_2
XFILLER_0_74_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06486_ final_design.reqhand.instruction\[19\] final_design.data_from_mem\[19\] net971
+ vssd1 vssd1 vccd1 vccd1 _01437_ sky130_fd_sc_hd__mux2_4
X_14194__1252 vssd1 vssd1 vccd1 vccd1 _14194__1252/HI net1252 sky130_fd_sc_hd__conb_1
XANTENNA__06733__S1 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08225_ final_design.cpu.reg_window\[203\] final_design.cpu.reg_window\[235\] net835
+ vssd1 vssd1 vccd1 vccd1 _03176_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout1150_A net1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout506_A net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_2889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09588__B1 net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08156_ final_design.cpu.reg_window\[271\] final_design.cpu.reg_window\[303\] net810
+ vssd1 vssd1 vccd1 vccd1 _03107_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_2108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_2119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11395__B1 net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07063__A1 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07107_ net881 _02051_ _02057_ _02044_ _02045_ vssd1 vssd1 vccd1 vccd1 _02058_ sky130_fd_sc_hd__a32oi_4
X_08087_ _01750_ _02896_ vssd1 vssd1 vccd1 vccd1 _03038_ sky130_fd_sc_hd__and2b_1
XANTENNA__14083__RESET_B net1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1036_X net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07177__S net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07038_ final_design.cpu.reg_window\[590\] final_design.cpu.reg_window\[622\] net894
+ vssd1 vssd1 vccd1 vccd1 _01989_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_1823 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout496_X net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout875_A net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11698__A1 net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08563__A1 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1889 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input1_X net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08989_ net621 _03921_ _03924_ _03655_ vssd1 vssd1 vccd1 vccd1 _03925_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout663_X net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10370__B2 final_design.data_from_mem\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11427__S net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10951_ _05677_ _05678_ _05651_ vssd1 vssd1 vccd1 vccd1 _05679_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_74_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13670_ clknet_leaf_50_clk _00901_ net1172 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[658\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11870__A1 _06017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10882_ _05611_ _05612_ _05590_ _05593_ vssd1 vssd1 vccd1 vccd1 _05613_ sky130_fd_sc_hd__a211o_1
XFILLER_0_32_1903 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09421__A net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12621_ net2022 final_design.reqhand.data_from_UART\[7\] _05080_ vssd1 vssd1 vccd1
+ vccd1 _01314_ sky130_fd_sc_hd__mux2_1
XANTENNA__09815__A1 net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12552_ _06215_ net354 net324 net2410 vssd1 vssd1 vccd1 vccd1 _01256_ sky130_fd_sc_hd__a22o_1
XANTENNA__10286__B net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11503_ net2446 net228 net522 vssd1 vssd1 vccd1 vccd1 _00372_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12483_ _06143_ net351 net333 net1968 vssd1 vssd1 vccd1 vccd1 _01189_ sky130_fd_sc_hd__a22o_1
X_14222_ final_design.h_out vssd1 vssd1 vccd1 vccd1 net172 sky130_fd_sc_hd__clkbuf_1
X_11434_ net2007 net190 net312 vssd1 vssd1 vccd1 vccd1 _00331_ sky130_fd_sc_hd__mux2_1
XANTENNA__06780__A net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09043__A2 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11386__B1 _05947_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11925__A2 net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14153_ clknet_leaf_18_clk _01327_ net1108 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.data_to_VGA\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_11365_ net436 net582 _06053_ net316 net1613 vssd1 vssd1 vccd1 vccd1 _00301_ sky130_fd_sc_hd__a32o_1
XFILLER_0_22_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13104_ clknet_leaf_33_clk _00335_ net1235 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[92\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06801__A1 final_design.data_from_mem\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10316_ net1463 net1011 net988 final_design.data_from_mem\[1\] vssd1 vssd1 vccd1
+ vccd1 _00073_ sky130_fd_sc_hd__a22o_1
X_14084_ clknet_leaf_24_clk _01281_ net1163 vssd1 vssd1 vccd1 vccd1 final_design.reqhand.instruction\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_11296_ _01881_ net641 _05991_ _05992_ net658 vssd1 vssd1 vccd1 vccd1 _05993_ sky130_fd_sc_hd__a221o_1
X_13035_ clknet_leaf_53_clk _00266_ net1187 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_10247_ final_design.uart.BAUD_counter\[17\] final_design.uart.BAUD_counter\[16\]
+ _05114_ vssd1 vssd1 vccd1 vccd1 _05118_ sky130_fd_sc_hd__and3_1
XFILLER_0_20_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1120 net1127 vssd1 vssd1 vccd1 vccd1 net1120 sky130_fd_sc_hd__buf_2
XANTENNA__12350__A2 net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1131 net1167 vssd1 vssd1 vccd1 vccd1 net1131 sky130_fd_sc_hd__clkbuf_2
Xfanout1142 net1150 vssd1 vssd1 vccd1 vccd1 net1142 sky130_fd_sc_hd__clkbuf_4
XANTENNA_clkbuf_leaf_8_clk_X clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10178_ final_design.uart.BAUD_counter\[17\] final_design.uart.BAUD_counter\[16\]
+ final_design.uart.BAUD_counter\[19\] final_design.uart.BAUD_counter\[18\] vssd1
+ vssd1 vccd1 vccd1 _05068_ sky130_fd_sc_hd__or4_1
Xfanout1153 net1162 vssd1 vssd1 vccd1 vccd1 net1153 sky130_fd_sc_hd__clkbuf_4
XANTENNA__13942__CLK clknet_leaf_59_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10361__B2 final_design.data_from_mem\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1164 net1165 vssd1 vssd1 vccd1 vccd1 net1164 sky130_fd_sc_hd__clkbuf_2
Xfanout1175 net1176 vssd1 vssd1 vccd1 vccd1 net1175 sky130_fd_sc_hd__clkbuf_2
XANTENNA__06660__S0 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1186 net1192 vssd1 vssd1 vccd1 vccd1 net1186 sky130_fd_sc_hd__clkbuf_4
Xfanout1197 net1245 vssd1 vssd1 vccd1 vccd1 net1197 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08306__A1 net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13937_ clknet_leaf_34_clk _01168_ net1243 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[925\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11310__B1 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13868_ clknet_leaf_46_clk _01099_ net1217 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[856\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11861__A1 net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12819_ net1367 vssd1 vssd1 vccd1 vccd1 _00260_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__11580__B _06016_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12168__S net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13799_ clknet_leaf_61_clk _01030_ net1124 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[787\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_1801 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09282__A2 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1845 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13322__CLK clknet_leaf_59_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_1891 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_1889 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08010_ _02948_ _02949_ _02960_ net879 vssd1 vssd1 vccd1 vccd1 _02961_ sky130_fd_sc_hd__a22o_4
XFILLER_0_71_189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_74_2720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_1391 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold603 final_design.cpu.reg_window\[934\] vssd1 vssd1 vccd1 vccd1 net1945 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07045__A1 net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_2731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold614 final_design.cpu.reg_window\[1019\] vssd1 vssd1 vccd1 vccd1 net1956 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06479__S0 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_2742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold625 final_design.cpu.reg_window\[328\] vssd1 vssd1 vccd1 vccd1 net1967 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13472__CLK clknet_leaf_11_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold636 final_design.cpu.reg_window\[87\] vssd1 vssd1 vccd1 vccd1 net1978 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold647 final_design.cpu.reg_window\[335\] vssd1 vssd1 vccd1 vccd1 net1989 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_70_2606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold658 final_design.cpu.reg_window\[932\] vssd1 vssd1 vccd1 vccd1 net2000 sky130_fd_sc_hd__dlygate4sd3_1
X_09961_ _04871_ _04876_ _04878_ net725 vssd1 vssd1 vccd1 vccd1 _04880_ sky130_fd_sc_hd__a211o_1
Xhold669 final_design.cpu.reg_window\[800\] vssd1 vssd1 vccd1 vccd1 net2011 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09417__S0 net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08912_ _01692_ _02467_ net621 vssd1 vssd1 vccd1 vccd1 _03856_ sky130_fd_sc_hd__a21oi_1
X_09892_ _02325_ net483 net441 vssd1 vssd1 vccd1 vccd1 _04811_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_42_1586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12341__A2 net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08843_ final_design.CPU_instr_adr\[19\] final_design.CPU_instr_adr\[18\] _03793_
+ vssd1 vssd1 vccd1 vccd1 _03794_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout191_A _06038_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06556__B1 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10352__A1 net13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10352__B2 final_design.data_from_mem\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_2513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout289_A net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_2524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08774_ _03698_ _03724_ _03697_ vssd1 vssd1 vccd1 vccd1 _03725_ sky130_fd_sc_hd__a21o_1
XFILLER_0_20_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_2535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07725_ final_design.cpu.reg_window\[282\] final_design.cpu.reg_window\[314\] net863
+ vssd1 vssd1 vccd1 vccd1 _02676_ sky130_fd_sc_hd__mux2_1
XANTENNA__11301__B1 net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07656_ net607 _02602_ _02577_ _01566_ vssd1 vssd1 vccd1 vccd1 _02607_ sky130_fd_sc_hd__o211a_1
XFILLER_0_71_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07460__S net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06607_ _01554_ _01555_ _01556_ _01557_ net776 net794 vssd1 vssd1 vccd1 vccd1 _01558_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__11490__B net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07587_ _02534_ _02535_ _02536_ _02537_ net685 net703 vssd1 vssd1 vccd1 vccd1 _02538_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_53_1671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout623_A _02506_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout244_X net244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10407__A2 net1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09326_ _04056_ _04243_ _04244_ vssd1 vssd1 vccd1 vccd1 _04245_ sky130_fd_sc_hd__o21a_1
X_06538_ _01456_ _01465_ _01474_ _01480_ vssd1 vssd1 vccd1 vccd1 _01489_ sky130_fd_sc_hd__or4_4
XFILLER_0_35_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09257_ _04175_ net450 _04174_ vssd1 vssd1 vccd1 vccd1 _04176_ sky130_fd_sc_hd__and3b_1
XFILLER_0_8_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout411_X net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06469_ final_design.reqhand.instruction\[15\] final_design.data_from_mem\[15\] net971
+ vssd1 vssd1 vccd1 vccd1 _01420_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1153_X net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13815__CLK clknet_leaf_58_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08208_ net716 _03158_ net874 vssd1 vssd1 vccd1 vccd1 _03159_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_1_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09188_ net489 _04055_ vssd1 vssd1 vccd1 vccd1 _04107_ sky130_fd_sc_hd__nor2_2
X_08139_ final_design.cpu.reg_window\[845\] final_design.cpu.reg_window\[877\] net855
+ vssd1 vssd1 vccd1 vccd1 _03090_ sky130_fd_sc_hd__mux2_1
X_11150_ _04805_ net654 _05843_ _05863_ vssd1 vssd1 vccd1 vccd1 _05864_ sky130_fd_sc_hd__a211oi_2
XANTENNA_fanout780_X net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13965__CLK clknet_leaf_48_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout878_X net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10101_ final_design.vga.h_current_state\[0\] final_design.vga.h_current_state\[1\]
+ _05015_ vssd1 vssd1 vccd1 vccd1 _05017_ sky130_fd_sc_hd__and3_2
X_11081_ net91 net1047 vssd1 vssd1 vccd1 vccd1 _05803_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_8_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07635__S net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12332__A2 net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10032_ _02836_ _04162_ _04158_ vssd1 vssd1 vccd1 vccd1 _04951_ sky130_fd_sc_hd__or3b_1
XANTENNA__11665__B net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10343__B2 final_design.data_from_mem\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09135__B _04053_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input17_A DAT_I[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12096__A1 net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11983_ _06185_ net290 net407 net1764 vssd1 vssd1 vccd1 vccd1 _00716_ sky130_fd_sc_hd__a22o_1
XFILLER_0_19_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11681__A net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13722_ clknet_leaf_64_clk _00953_ net1075 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[710\]
+ sky130_fd_sc_hd__dfrtp_1
X_10934_ _01386_ _05649_ _05658_ _05661_ vssd1 vssd1 vccd1 vccd1 _05663_ sky130_fd_sc_hd__nor4_1
XANTENNA__09422__Y _04341_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13345__CLK clknet_leaf_48_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13653_ clknet_leaf_58_clk _00884_ net1132 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[641\]
+ sky130_fd_sc_hd__dfrtp_1
X_10865_ net962 _05596_ vssd1 vssd1 vccd1 vccd1 _05597_ sky130_fd_sc_hd__or2_1
XFILLER_0_67_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_1793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12399__A2 net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12604_ net1399 net996 net982 final_design.data_from_mem\[22\] vssd1 vssd1 vccd1
+ vccd1 _01297_ sky130_fd_sc_hd__a22o_1
XFILLER_0_66_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13584_ clknet_leaf_36_clk _00815_ net1236 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[572\]
+ sky130_fd_sc_hd__dfrtp_1
X_10796_ net76 _05511_ _05530_ vssd1 vssd1 vccd1 vccd1 _05531_ sky130_fd_sc_hd__a21o_1
XFILLER_0_27_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12535_ _06198_ net346 net322 net2235 vssd1 vssd1 vccd1 vccd1 _01239_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_26_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13495__CLK clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1829 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06714__S net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12466_ _06126_ net349 net331 net2144 vssd1 vssd1 vccd1 vccd1 _01172_ sky130_fd_sc_hd__a22o_1
X_14205_ net1263 vssd1 vssd1 vccd1 vccd1 gpio_oeb[17] sky130_fd_sc_hd__buf_2
XFILLER_0_62_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11417_ net1588 net243 net310 vssd1 vssd1 vccd1 vccd1 _00314_ sky130_fd_sc_hd__mux2_1
XANTENNA__09567__A3 net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12397_ net553 _06268_ net339 net2422 vssd1 vssd1 vccd1 vccd1 _01107_ sky130_fd_sc_hd__a22o_1
X_14136_ clknet_leaf_17_clk final_design.vga.h_next_count\[5\] net1113 vssd1 vssd1
+ vccd1 vccd1 final_design.VGA_data_control.h_count\[5\] sky130_fd_sc_hd__dfrtp_2
X_11348_ net650 net190 vssd1 vssd1 vccd1 vccd1 _06039_ sky130_fd_sc_hd__and2_1
XANTENNA__07983__C1 _01908_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11856__A net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12451__S net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14067_ clknet_leaf_15_clk _00030_ net1093 vssd1 vssd1 vccd1 vccd1 final_design.uart.BAUD_counter\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_11279_ net643 _05977_ _05976_ net658 vssd1 vssd1 vccd1 vccd1 _05978_ sky130_fd_sc_hd__a211o_1
XANTENNA__07545__S net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13018_ clknet_leaf_1_clk _00249_ net1081 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_78_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10334__B2 final_design.data_from_mem\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14120__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07750__A2 _02698_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06553__A3 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12087__A1 net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07189__S1 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07510_ _01825_ _02460_ vssd1 vssd1 vccd1 vccd1 _02461_ sky130_fd_sc_hd__or2_1
X_08490_ final_design.cpu.reg_window\[963\] final_design.cpu.reg_window\[995\] net824
+ vssd1 vssd1 vccd1 vccd1 _03441_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_1557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07441_ final_design.reqhand.instruction\[8\] final_design.data_from_mem\[8\] net972
+ vssd1 vssd1 vccd1 vccd1 _02392_ sky130_fd_sc_hd__mux2_1
XANTENNA__12785__16_A clknet_leaf_28_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13838__CLK clknet_leaf_45_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08138__S0 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10000__A _04918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07372_ _02319_ _02320_ _02321_ _02322_ net768 net781 vssd1 vssd1 vccd1 vccd1 _02323_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_11_1817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09111_ final_design.CPU_instr_adr\[0\] _02425_ vssd1 vssd1 vccd1 vccd1 _04031_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_21_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_2804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11530__S net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_2815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09042_ net622 _03971_ vssd1 vssd1 vccd1 vccd1 _03972_ sky130_fd_sc_hd__nor2_1
XANTENNA__12862__CLK clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13988__CLK clknet_leaf_54_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold400 final_design.cpu.reg_window\[670\] vssd1 vssd1 vccd1 vccd1 net1742 sky130_fd_sc_hd__dlygate4sd3_1
Xhold411 final_design.cpu.reg_window\[644\] vssd1 vssd1 vccd1 vccd1 net1753 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout204_A _05989_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold422 final_design.cpu.reg_window\[473\] vssd1 vssd1 vccd1 vccd1 net1764 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11365__A3 _06053_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12562__A2 net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold433 final_design.cpu.reg_window\[366\] vssd1 vssd1 vccd1 vccd1 net1775 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold444 final_design.cpu.reg_window\[649\] vssd1 vssd1 vccd1 vccd1 net1786 sky130_fd_sc_hd__dlygate4sd3_1
Xhold455 final_design.cpu.reg_window\[47\] vssd1 vssd1 vccd1 vccd1 net1797 sky130_fd_sc_hd__dlygate4sd3_1
Xhold466 final_design.cpu.reg_window\[36\] vssd1 vssd1 vccd1 vccd1 net1808 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_971 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold477 final_design.cpu.reg_window\[838\] vssd1 vssd1 vccd1 vccd1 net1819 sky130_fd_sc_hd__dlygate4sd3_1
Xhold488 final_design.cpu.reg_window\[774\] vssd1 vssd1 vccd1 vccd1 net1830 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout902 net904 vssd1 vssd1 vccd1 vccd1 net902 sky130_fd_sc_hd__clkbuf_4
XANTENNA__13218__CLK clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09944_ _04861_ _04862_ _04858_ _04860_ vssd1 vssd1 vccd1 vccd1 _04863_ sky130_fd_sc_hd__a2bb2o_1
Xfanout913 net917 vssd1 vssd1 vccd1 vccd1 net913 sky130_fd_sc_hd__clkbuf_4
Xhold499 final_design.cpu.reg_window\[697\] vssd1 vssd1 vccd1 vccd1 net1841 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1113_A net1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08518__A1 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout924 net927 vssd1 vssd1 vccd1 vccd1 net924 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_5_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout935 net952 vssd1 vssd1 vccd1 vccd1 net935 sky130_fd_sc_hd__clkbuf_4
Xfanout946 net951 vssd1 vssd1 vccd1 vccd1 net946 sky130_fd_sc_hd__clkbuf_4
XANTENNA_input9_A DAT_I[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout957 _04043_ vssd1 vssd1 vccd1 vccd1 net957 sky130_fd_sc_hd__clkbuf_4
X_09875_ net532 net530 net452 vssd1 vssd1 vccd1 vccd1 _04794_ sky130_fd_sc_hd__mux2_1
Xhold1100 final_design.cpu.reg_window\[306\] vssd1 vssd1 vccd1 vccd1 net2442 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout573_A net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10325__B2 final_design.data_from_mem\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout979 net981 vssd1 vssd1 vccd1 vccd1 net979 sky130_fd_sc_hd__clkbuf_4
Xhold1111 final_design.cpu.reg_window\[109\] vssd1 vssd1 vccd1 vccd1 net2453 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1122 final_design.cpu.reg_window\[480\] vssd1 vssd1 vccd1 vccd1 net2464 sky130_fd_sc_hd__dlygate4sd3_1
X_08826_ final_design.CPU_instr_adr\[29\] _01539_ _03776_ vssd1 vssd1 vccd1 vccd1
+ _03777_ sky130_fd_sc_hd__a21oi_1
Xhold1133 final_design.cpu.reg_window\[310\] vssd1 vssd1 vccd1 vccd1 net2475 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1144 final_design.cpu.reg_window\[34\] vssd1 vssd1 vccd1 vccd1 net2486 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_77_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1155 final_design.cpu.reg_window\[992\] vssd1 vssd1 vccd1 vccd1 net2497 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12078__A1 net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1166 final_design.cpu.reg_window\[256\] vssd1 vssd1 vccd1 vccd1 net2508 sky130_fd_sc_hd__dlygate4sd3_1
X_08757_ _03706_ _03707_ vssd1 vssd1 vccd1 vccd1 _03708_ sky130_fd_sc_hd__nor2_1
Xhold1177 final_design.cpu.reg_window\[124\] vssd1 vssd1 vccd1 vccd1 net2519 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout361_X net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1188 final_design.uart.BAUD_counter\[30\] vssd1 vssd1 vccd1 vccd1 net2530 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1199 final_design.CPU_instr_adr\[25\] vssd1 vssd1 vccd1 vccd1 net2541 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout838_A net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout459_X net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07708_ final_design.cpu.reg_window\[667\] final_design.cpu.reg_window\[699\] net861
+ vssd1 vssd1 vccd1 vccd1 _02659_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08688_ net609 _03550_ _02419_ _02423_ vssd1 vssd1 vccd1 vccd1 _03639_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_0_174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06927__S1 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07639_ final_design.cpu.reg_window\[860\] final_design.cpu.reg_window\[892\] net866
+ vssd1 vssd1 vccd1 vccd1 _02590_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_0_196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout626_X net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07978__X _02929_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10650_ _05368_ _05390_ vssd1 vssd1 vccd1 vccd1 _05392_ sky130_fd_sc_hd__or2_1
XFILLER_0_82_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11589__B1 net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09309_ _04091_ _04227_ vssd1 vssd1 vccd1 vccd1 _04228_ sky130_fd_sc_hd__and2_1
XANTENNA__12250__A1 net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10581_ _05326_ vssd1 vssd1 vccd1 vccd1 _05327_ sky130_fd_sc_hd__inv_2
XFILLER_0_64_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11440__S net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12320_ net1824 net193 net366 vssd1 vssd1 vccd1 vccd1 _01034_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_40_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10564__B net250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12251_ net585 _06180_ net512 net374 net1551 vssd1 vssd1 vccd1 vccd1 _00967_ sky130_fd_sc_hd__a32o_1
X_11202_ _04903_ net651 net588 _05909_ vssd1 vssd1 vccd1 vccd1 _05910_ sky130_fd_sc_hd__o211a_2
XANTENNA__12553__A2 net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12182_ net1846 net202 net382 vssd1 vssd1 vccd1 vccd1 _00901_ sky130_fd_sc_hd__mux2_1
X_11133_ _05840_ _05846_ vssd1 vssd1 vccd1 vccd1 _05848_ sky130_fd_sc_hd__or2_4
XANTENNA__14143__CLK clknet_leaf_19_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11064_ net1056 _05785_ _05786_ vssd1 vssd1 vccd1 vccd1 _05787_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10316__B2 final_design.data_from_mem\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10015_ _04220_ _04693_ _04932_ _04933_ vssd1 vssd1 vccd1 vccd1 _04934_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_34_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_3008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_3019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output123_A net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08368__S0 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09152__Y _04071_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11966_ _06168_ net277 net404 net1986 vssd1 vssd1 vccd1 vccd1 _00699_ sky130_fd_sc_hd__a22o_1
XFILLER_0_25_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10917_ _05624_ _05646_ _05645_ vssd1 vssd1 vccd1 vccd1 _05647_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12962__RESET_B net1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13705_ clknet_leaf_36_clk _00936_ net1229 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[693\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_15_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11897_ net213 net2457 net272 vssd1 vssd1 vccd1 vccd1 _00639_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13636_ clknet_leaf_54_clk _00867_ net1179 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[624\]
+ sky130_fd_sc_hd__dfrtp_1
X_10848_ _05578_ _05579_ vssd1 vssd1 vccd1 vccd1 _05581_ sky130_fd_sc_hd__nor2_1
XANTENNA__12885__CLK clknet_leaf_19_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07248__A1 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11044__A2 net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12446__S net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12241__A1 net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13567_ clknet_leaf_8_clk _00798_ net1153 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[555\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10779_ _05487_ _05489_ _05513_ vssd1 vssd1 vccd1 vccd1 _05515_ sky130_fd_sc_hd__or3b_1
XFILLER_0_70_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08996__A1 net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11203__X _05911_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12518_ _06180_ net357 net328 net1873 vssd1 vssd1 vccd1 vccd1 _01223_ sky130_fd_sc_hd__a22o_1
XANTENNA__11595__A3 _06153_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13498_ clknet_leaf_58_clk _00729_ net1128 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[486\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12449_ net2109 net203 net336 vssd1 vssd1 vccd1 vccd1 _01156_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12544__A2 net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11752__A0 net223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_256 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14119_ clknet_leaf_17_clk final_design.vga.h_next_state\[1\] net1114 vssd1 vssd1
+ vccd1 vccd1 final_design.vga.h_current_state\[1\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__12181__S net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout209 net211 vssd1 vssd1 vccd1 vccd1 net209 sky130_fd_sc_hd__buf_2
X_07990_ final_design.cpu.reg_window\[400\] final_design.cpu.reg_window\[432\] net846
+ vssd1 vssd1 vccd1 vccd1 _02941_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_wire541_A _01995_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06941_ final_design.cpu.reg_window\[209\] final_design.cpu.reg_window\[241\] net928
+ vssd1 vssd1 vccd1 vccd1 _01892_ sky130_fd_sc_hd__mux2_1
XANTENNA__13510__CLK clknet_leaf_51_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1733 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09660_ _04362_ _04363_ net478 vssd1 vssd1 vccd1 vccd1 _04579_ sky130_fd_sc_hd__o21ai_2
XPHY_EDGE_ROW_19_Left_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06872_ _01504_ _01822_ vssd1 vssd1 vccd1 vccd1 _01823_ sky130_fd_sc_hd__nand2_2
XFILLER_0_78_1777 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08611_ net531 _03386_ vssd1 vssd1 vccd1 vccd1 _03562_ sky130_fd_sc_hd__nor2_1
X_09591_ net729 _04482_ _04502_ _04508_ vssd1 vssd1 vccd1 vccd1 _04510_ sky130_fd_sc_hd__nand4_2
XFILLER_0_55_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13660__CLK clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08542_ _03489_ _03490_ _03491_ _03492_ net680 net700 vssd1 vssd1 vccd1 vccd1 _03493_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__11283__A2 net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08473_ _03420_ _03422_ vssd1 vssd1 vccd1 vccd1 _03424_ sky130_fd_sc_hd__or2_1
XFILLER_0_37_1496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07424_ net760 _02374_ vssd1 vssd1 vccd1 vccd1 _02375_ sky130_fd_sc_hd__or2_1
XANTENNA__14016__CLK clknet_leaf_11_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12232__A1 net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07355_ final_design.cpu.reg_window\[67\] final_design.cpu.reg_window\[99\] net905
+ vssd1 vssd1 vccd1 vccd1 _02306_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_28_Left_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout321_A _04047_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1063_A net1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_936 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07286_ _02233_ _02234_ _02235_ _02236_ net767 net787 vssd1 vssd1 vccd1 vccd1 _02237_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__10384__B net1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09025_ final_design.CPU_instr_adr\[12\] _03789_ vssd1 vssd1 vccd1 vccd1 _03957_
+ sky130_fd_sc_hd__xnor2_1
XANTENNA__14166__CLK clknet_leaf_18_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13040__CLK clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout207_X net207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12535__A2 net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09936__B1 net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold230 final_design.cpu.reg_window\[970\] vssd1 vssd1 vccd1 vccd1 net1572 sky130_fd_sc_hd__dlygate4sd3_1
Xhold241 final_design.cpu.reg_window\[709\] vssd1 vssd1 vccd1 vccd1 net1583 sky130_fd_sc_hd__dlygate4sd3_1
Xhold252 final_design.cpu.reg_window\[717\] vssd1 vssd1 vccd1 vccd1 net1594 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11743__A0 net244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout788_A _01418_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold263 final_design.cpu.reg_window\[662\] vssd1 vssd1 vccd1 vccd1 net1605 sky130_fd_sc_hd__dlygate4sd3_1
Xhold274 final_design.cpu.reg_window\[776\] vssd1 vssd1 vccd1 vccd1 net1616 sky130_fd_sc_hd__dlygate4sd3_1
Xhold285 final_design.cpu.reg_window\[186\] vssd1 vssd1 vccd1 vccd1 net1627 sky130_fd_sc_hd__dlygate4sd3_1
Xhold296 final_design.cpu.reg_window\[254\] vssd1 vssd1 vccd1 vccd1 net1638 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1116_X net1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout710 net715 vssd1 vssd1 vccd1 vccd1 net710 sky130_fd_sc_hd__buf_4
XANTENNA_clkbuf_leaf_33_clk_X clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout721 _01720_ vssd1 vssd1 vccd1 vccd1 net721 sky130_fd_sc_hd__clkbuf_4
XANTENNA__13190__CLK clknet_leaf_51_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout732 _01491_ vssd1 vssd1 vccd1 vccd1 net732 sky130_fd_sc_hd__clkbuf_4
X_09927_ _04843_ _04845_ _04831_ vssd1 vssd1 vccd1 vccd1 _04846_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_37_Left_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout743 _01476_ vssd1 vssd1 vccd1 vccd1 net743 sky130_fd_sc_hd__buf_4
XANTENNA_fanout955_A net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout576_X net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout754 net755 vssd1 vssd1 vccd1 vccd1 net754 sky130_fd_sc_hd__clkbuf_2
Xfanout765 net766 vssd1 vssd1 vccd1 vccd1 net765 sky130_fd_sc_hd__buf_4
Xfanout776 net777 vssd1 vssd1 vccd1 vccd1 net776 sky130_fd_sc_hd__buf_4
XFILLER_0_77_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09858_ _03294_ net446 _04775_ _04776_ net263 vssd1 vssd1 vccd1 vccd1 _04777_ sky130_fd_sc_hd__o2111ai_1
Xfanout787 net788 vssd1 vssd1 vccd1 vccd1 net787 sky130_fd_sc_hd__buf_4
XANTENNA__09703__A3 _04579_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout798 net800 vssd1 vssd1 vccd1 vccd1 net798 sky130_fd_sc_hd__buf_2
XFILLER_0_38_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08809_ final_design.CPU_instr_adr\[21\] _01788_ vssd1 vssd1 vccd1 vccd1 _03760_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_57_1839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09789_ _04219_ _04343_ _04221_ vssd1 vssd1 vccd1 vccd1 _04708_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout743_X net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_48_clk_X clknet_leaf_48_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11435__S net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11820_ net219 net1860 net264 vssd1 vssd1 vccd1 vccd1 _00572_ sky130_fd_sc_hd__mux2_1
X_11751_ net206 net2223 net416 vssd1 vssd1 vccd1 vccd1 _00514_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout910_X net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1438 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10702_ _05438_ _05441_ vssd1 vssd1 vccd1 vccd1 _05442_ sky130_fd_sc_hd__nand2_1
X_11682_ net430 net570 _06199_ net295 net1672 vssd1 vssd1 vccd1 vccd1 _00472_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_46_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13421_ clknet_leaf_44_clk _00652_ net1200 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[409\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_23_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10633_ _05354_ _05375_ vssd1 vssd1 vccd1 vccd1 _05376_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_3_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_23_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_1913 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1269 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06772__B _01722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08978__A1 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13352_ clknet_leaf_35_clk _00583_ net1241 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[340\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input84_A memory_size[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10564_ _04724_ net250 vssd1 vssd1 vccd1 vccd1 _05310_ sky130_fd_sc_hd__nor2_1
XANTENNA__10785__A1 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10785__B2 net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12303_ net1830 net238 net364 vssd1 vssd1 vccd1 vccd1 _01017_ sky130_fd_sc_hd__mux2_1
XANTENNA__11982__B1 net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13283_ clknet_leaf_1_clk _00514_ net1074 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[271\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07650__A1 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10495_ _05234_ _05242_ _05243_ net58 vssd1 vssd1 vccd1 vccd1 _05245_ sky130_fd_sc_hd__a31o_1
XANTENNA__12526__A2 net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12234_ net563 _06164_ net505 net372 net1545 vssd1 vssd1 vccd1 vccd1 _00951_ sky130_fd_sc_hd__a32o_1
XFILLER_0_66_1692 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13533__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11734__B1 net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12165_ net2294 net228 net381 vssd1 vssd1 vccd1 vccd1 _00884_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_36_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07095__S net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11116_ final_design.uart.bits_received\[2\] _05832_ vssd1 vssd1 vccd1 vccd1 _05834_
+ sky130_fd_sc_hd__xnor2_1
X_12096_ net2064 net228 net389 vssd1 vssd1 vccd1 vccd1 _00820_ sky130_fd_sc_hd__mux2_1
X_11047_ net966 _05770_ _05768_ vssd1 vssd1 vccd1 vccd1 _05771_ sky130_fd_sc_hd__a21o_1
XANTENNA__13683__CLK clknet_leaf_38_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1917 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput9 DAT_I[16] vssd1 vssd1 vccd1 vccd1 net9 sky130_fd_sc_hd__clkbuf_1
X_12998_ net1329 _00229_ net1195 vssd1 vssd1 vccd1 vccd1 final_design.CPU_instr_adr\[18\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__14039__CLK clknet_leaf_15_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07013__S0 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11949_ _06150_ net290 net411 net2044 vssd1 vssd1 vccd1 vccd1 _00684_ sky130_fd_sc_hd__a22o_1
XFILLER_0_59_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10473__A0 final_design.CPU_instr_adr\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1901 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12214__A1 net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13619_ clknet_leaf_40_clk _00850_ net1206 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[607\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12176__S net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13063__CLK clknet_leaf_62_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07140_ _02078_ _02079_ _02090_ net883 vssd1 vssd1 vccd1 vccd1 _02091_ sky130_fd_sc_hd__a22oi_4
XFILLER_0_55_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11973__B1 net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07071_ final_design.cpu.reg_window\[973\] final_design.cpu.reg_window\[1005\] net934
+ vssd1 vssd1 vccd1 vccd1 _02022_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12517__A2 net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09394__A1 net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12900__CLK clknet_leaf_25_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07973_ final_design.cpu.reg_window\[657\] final_design.cpu.reg_window\[689\] net848
+ vssd1 vssd1 vccd1 vccd1 _02924_ sky130_fd_sc_hd__mux2_1
X_09712_ _04626_ _04630_ vssd1 vssd1 vccd1 vccd1 _04631_ sky130_fd_sc_hd__or2_1
X_06924_ final_design.cpu.reg_window\[658\] final_design.cpu.reg_window\[690\] net925
+ vssd1 vssd1 vccd1 vccd1 _01875_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12150__A0 net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09643_ net486 _04559_ _04560_ _04224_ _04092_ vssd1 vssd1 vccd1 vccd1 _04562_ sky130_fd_sc_hd__a221o_1
X_06855_ final_design.cpu.reg_window\[916\] final_design.cpu.reg_window\[948\] net950
+ vssd1 vssd1 vccd1 vccd1 _01806_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout369_A _06274_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09574_ _04492_ _04488_ net318 _04067_ vssd1 vssd1 vccd1 vccd1 _04493_ sky130_fd_sc_hd__o2bb2a_1
X_06786_ net760 _01736_ vssd1 vssd1 vccd1 vccd1 _01737_ sky130_fd_sc_hd__nor2_1
XFILLER_0_56_1861 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08525_ final_design.cpu.reg_window\[642\] final_design.cpu.reg_window\[674\] net832
+ vssd1 vssd1 vccd1 vccd1 _03476_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_1834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12453__A1 net196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11256__A2 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1180_A net1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_60_clk_A clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_62_clk clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_62_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__13406__CLK clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08456_ final_design.cpu.reg_window\[900\] final_design.cpu.reg_window\[932\] net819
+ vssd1 vssd1 vccd1 vccd1 _03407_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_1567 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07407_ final_design.data_from_mem\[9\] net970 _02357_ vssd1 vssd1 vccd1 vccd1 _02358_
+ sky130_fd_sc_hd__o21a_2
X_08387_ _03334_ _03335_ _03336_ _03337_ net677 net698 vssd1 vssd1 vccd1 vccd1 _03338_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout324_X net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout703_A net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07338_ final_design.cpu.reg_window\[644\] final_design.cpu.reg_window\[676\] net900
+ vssd1 vssd1 vccd1 vccd1 _02289_ sky130_fd_sc_hd__mux2_1
XANTENNA__13556__CLK clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11964__B1 net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07269_ _02216_ _02217_ _02218_ _02219_ net767 net787 vssd1 vssd1 vccd1 vccd1 _02220_
+ sky130_fd_sc_hd__mux4_1
X_09008_ net620 _03938_ net255 vssd1 vssd1 vccd1 vccd1 _03942_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12508__A2 net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11497__Y _06116_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10280_ _05138_ net797 _05137_ vssd1 vssd1 vccd1 vccd1 _00027_ sky130_fd_sc_hd__and3b_1
XFILLER_0_44_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11716__B1 net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout693_X net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout860_X net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout958_X net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout540 _02026_ vssd1 vssd1 vccd1 vccd1 net540 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_50_1914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout551 _01750_ vssd1 vssd1 vccd1 vccd1 net551 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_50_1925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout562 net571 vssd1 vssd1 vccd1 vccd1 net562 sky130_fd_sc_hd__clkbuf_2
Xfanout573 net576 vssd1 vssd1 vccd1 vccd1 net573 sky130_fd_sc_hd__clkbuf_4
X_13970_ clknet_leaf_39_clk _01201_ net1209 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[958\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout584 net585 vssd1 vssd1 vccd1 vccd1 net584 sky130_fd_sc_hd__buf_2
XANTENNA_clkbuf_leaf_13_clk_A clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12769__B net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout595 net596 vssd1 vssd1 vccd1 vccd1 net595 sky130_fd_sc_hd__buf_2
XANTENNA__09424__A net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12921_ clknet_leaf_50_clk _00159_ net1168 vssd1 vssd1 vccd1 vccd1 net143 sky130_fd_sc_hd__dfrtp_1
XANTENNA__11673__B net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12692__A1 _05008_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12852_ clknet_leaf_14_clk _00090_ net1106 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.ready_data\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_17_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11803_ net2516 net415 net290 _06046_ vssd1 vssd1 vccd1 vccd1 _00556_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_48_1843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12444__A1 net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_28_clk_A clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13086__CLK clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_53_clk clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_53_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_44_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_1809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11734_ net579 net423 _06225_ net296 net1697 vssd1 vssd1 vccd1 vccd1 _00498_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_44_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11665_ net178 net632 vssd1 vssd1 vccd1 vccd1 _06190_ sky130_fd_sc_hd__and2_1
XFILLER_0_68_1721 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10616_ net1054 _05356_ net1001 final_design.CPU_instr_adr\[8\] vssd1 vssd1 vccd1
+ vccd1 _05360_ sky130_fd_sc_hd__o2bb2a_1
X_13404_ clknet_leaf_5_clk _00635_ net1078 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[392\]
+ sky130_fd_sc_hd__dfrtp_1
X_11596_ net180 net636 vssd1 vssd1 vccd1 vccd1 _06154_ sky130_fd_sc_hd__and2_1
XANTENNA__10302__S0 net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11955__B1 net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13335_ clknet_leaf_6_clk _00566_ net1134 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[323\]
+ sky130_fd_sc_hd__dfrtp_1
X_10547_ _05273_ _05292_ vssd1 vssd1 vccd1 vccd1 _05294_ sky130_fd_sc_hd__and2_1
XFILLER_0_51_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12923__CLK clknet_leaf_30_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13266_ clknet_leaf_39_clk _00497_ net1205 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[254\]
+ sky130_fd_sc_hd__dfrtp_1
X_10478_ net47 _05223_ _05225_ _05227_ vssd1 vssd1 vccd1 vccd1 _05229_ sky130_fd_sc_hd__and4_1
X_12217_ net585 _06145_ net512 net378 net1842 vssd1 vssd1 vccd1 vccd1 _00935_ sky130_fd_sc_hd__a32o_1
XFILLER_0_27_1473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13197_ clknet_leaf_48_clk _00428_ net1200 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[185\]
+ sky130_fd_sc_hd__dfrtp_1
X_12148_ net202 net2406 net387 vssd1 vssd1 vccd1 vccd1 _00869_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_10_Right_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12079_ net574 _05990_ net508 net395 net1626 vssd1 vssd1 vccd1 vccd1 _00804_ sky130_fd_sc_hd__a32o_1
XFILLER_0_79_1861 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12683__B2 final_design.data_from_mem\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13429__CLK clknet_leaf_56_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10694__B1 net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06640_ final_design.cpu.reg_window\[667\] final_design.cpu.reg_window\[699\] net941
+ vssd1 vssd1 vccd1 vccd1 _01591_ sky130_fd_sc_hd__mux2_1
XANTENNA__12435__A1 net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06571_ net753 _01515_ net747 vssd1 vssd1 vccd1 vccd1 _01522_ sky130_fd_sc_hd__o21a_1
Xclkbuf_leaf_44_clk clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_44_clk sky130_fd_sc_hd__clkbuf_8
X_08310_ net610 _03257_ _03258_ net535 vssd1 vssd1 vccd1 vccd1 _03261_ sky130_fd_sc_hd__a211o_1
X_09290_ _02639_ net442 net438 _02638_ vssd1 vssd1 vccd1 vccd1 _04209_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_64_2390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13579__CLK clknet_leaf_52_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_2243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08241_ _03179_ _03180_ _03191_ net876 vssd1 vssd1 vccd1 vccd1 _03192_ sky130_fd_sc_hd__a22oi_4
XTAP_TAPCELL_ROW_60_2254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_14 net1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_2265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_25 _06257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12199__B1 net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08172_ final_design.cpu.reg_window\[719\] final_design.cpu.reg_window\[751\] net806
+ vssd1 vssd1 vccd1 vccd1 _03123_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09603__A2 net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11946__B1 net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07123_ final_design.cpu.reg_window\[11\] final_design.cpu.reg_window\[43\] net915
+ vssd1 vssd1 vccd1 vccd1 _02074_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07054_ final_design.cpu.reg_window\[461\] final_design.cpu.reg_window\[493\] net931
+ vssd1 vssd1 vccd1 vccd1 _02005_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_58_2172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput110 net110 vssd1 vssd1 vccd1 vccd1 ADR_O[18] sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_58_2183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput121 net121 vssd1 vssd1 vccd1 vccd1 ADR_O[28] sky130_fd_sc_hd__clkbuf_4
XANTENNA__13012__RESET_B net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_2194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput132 net132 vssd1 vssd1 vccd1 vccd1 ADR_O[9] sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_54_2036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput143 net143 vssd1 vssd1 vccd1 vccd1 DAT_O[18] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_54_2047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput154 net154 vssd1 vssd1 vccd1 vccd1 DAT_O[28] sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_54_2058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput165 net165 vssd1 vssd1 vccd1 vccd1 DAT_O[9] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_54_2069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11174__A1 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout486_A net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11774__A net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07956_ final_design.cpu.reg_window\[273\] final_design.cpu.reg_window\[305\] net850
+ vssd1 vssd1 vccd1 vccd1 _02907_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_1893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_1901 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06907_ final_design.cpu.reg_window\[274\] final_design.cpu.reg_window\[306\] net924
+ vssd1 vssd1 vccd1 vccd1 _01858_ sky130_fd_sc_hd__mux2_1
XANTENNA__07225__S0 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07887_ _02800_ _02801_ _02833_ _02835_ vssd1 vssd1 vccd1 vccd1 _02838_ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout274_X net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09626_ _02868_ _04544_ vssd1 vssd1 vccd1 vccd1 _04545_ sky130_fd_sc_hd__xnor2_1
X_06838_ _01785_ _01788_ vssd1 vssd1 vccd1 vccd1 _01789_ sky130_fd_sc_hd__nor2_1
XFILLER_0_78_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09557_ _04474_ _04475_ vssd1 vssd1 vccd1 vccd1 _04476_ sky130_fd_sc_hd__xnor2_1
XANTENNA__11229__A2 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout820_A net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout441_X net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06769_ final_design.data_from_mem\[23\] net969 _01719_ vssd1 vssd1 vccd1 vccd1 _01720_
+ sky130_fd_sc_hd__o21a_4
XANTENNA_fanout918_A net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout539_X net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_35_clk clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_35_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__10437__B1 net1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08508_ final_design.cpu.reg_window\[258\] final_design.cpu.reg_window\[290\] net838
+ vssd1 vssd1 vccd1 vccd1 _03459_ sky130_fd_sc_hd__mux2_1
X_09488_ net477 _04406_ vssd1 vssd1 vccd1 vccd1 _04407_ sky130_fd_sc_hd__nor2_1
X_08439_ _03387_ _03389_ vssd1 vssd1 vccd1 vccd1 _03390_ sky130_fd_sc_hd__nor2_1
XFILLER_0_68_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout706_X net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12946__CLK clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11450_ net227 net638 vssd1 vssd1 vccd1 vccd1 _06098_ sky130_fd_sc_hd__and2_1
XANTENNA__08763__B1_N final_design.CPU_instr_adr\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11937__B1 net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10401_ net1418 net1027 _05183_ net246 vssd1 vssd1 vccd1 vccd1 _00142_ sky130_fd_sc_hd__a22o_1
XFILLER_0_22_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11381_ net649 net182 vssd1 vssd1 vccd1 vccd1 _06068_ sky130_fd_sc_hd__and2_1
XFILLER_0_22_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13120_ clknet_leaf_12_clk _00351_ net1086 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[108\]
+ sky130_fd_sc_hd__dfrtp_1
X_10332_ net1651 net1010 net987 final_design.data_from_mem\[17\] vssd1 vssd1 vccd1
+ vccd1 _00089_ sky130_fd_sc_hd__a22o_1
XANTENNA__08323__A net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13051_ clknet_leaf_0_clk _00282_ net1062 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[39\]
+ sky130_fd_sc_hd__dfrtp_1
X_10263_ final_design.uart.BAUD_counter\[23\] final_design.uart.BAUD_counter\[22\]
+ _05124_ vssd1 vssd1 vccd1 vccd1 _05128_ sky130_fd_sc_hd__and3_1
XANTENNA__12362__B1 net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12002_ _06204_ net278 net400 net2284 vssd1 vssd1 vccd1 vccd1 _00733_ sky130_fd_sc_hd__a22o_1
XANTENNA_input47_A mem_adr_start[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10194_ final_design.uart.BAUD_counter\[1\] final_design.uart.BAUD_counter\[0\] vssd1
+ vssd1 vccd1 vccd1 _05083_ sky130_fd_sc_hd__or2_1
XANTENNA__10912__A1 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10912__B2 net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout370 net371 vssd1 vssd1 vccd1 vccd1 net370 sky130_fd_sc_hd__buf_4
Xfanout381 net383 vssd1 vssd1 vccd1 vccd1 net381 sky130_fd_sc_hd__buf_4
XANTENNA__09154__A net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout392 net393 vssd1 vssd1 vccd1 vccd1 net392 sky130_fd_sc_hd__buf_4
X_13953_ clknet_leaf_47_clk _01184_ net1199 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[941\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12665__B2 final_design.data_from_mem\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12904_ clknet_leaf_61_clk _00142_ net1136 vssd1 vssd1 vccd1 vccd1 net145 sky130_fd_sc_hd__dfrtp_1
X_13884_ clknet_leaf_5_clk _01115_ net1083 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[872\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_1319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_1488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12835_ clknet_leaf_19_clk _00073_ net1111 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.ready_data\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13721__CLK clknet_leaf_56_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_26_clk clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_26_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_57_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12766_ _06383_ _06396_ _06397_ _06400_ _06401_ vssd1 vssd1 vccd1 vccd1 _01354_ sky130_fd_sc_hd__a311o_1
XFILLER_0_33_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10979__A1 net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10979__B2 net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11717_ net192 net629 vssd1 vssd1 vccd1 vccd1 _06217_ sky130_fd_sc_hd__and2_1
X_12697_ final_design.VGA_data_control.v_count\[8\] final_design.VGA_data_control.v_count\[5\]
+ _01398_ _06336_ final_design.VGA_data_control.v_count\[7\] vssd1 vssd1 vccd1 vccd1
+ _06338_ sky130_fd_sc_hd__a32o_1
XFILLER_0_72_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11640__A2 net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13871__CLK clknet_leaf_42_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11648_ net586 net424 _06181_ net300 net2089 vssd1 vssd1 vccd1 vccd1 _00456_ sky130_fd_sc_hd__a32o_1
Xinput12 DAT_I[19] vssd1 vssd1 vccd1 vccd1 net12 sky130_fd_sc_hd__clkbuf_1
Xinput23 DAT_I[29] vssd1 vssd1 vccd1 vccd1 net23 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11928__B1 net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput34 en vssd1 vssd1 vccd1 vccd1 net34 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_29_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput45 mem_adr_start[18] vssd1 vssd1 vccd1 vccd1 net45 sky130_fd_sc_hd__clkbuf_1
XANTENNA__12454__S net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11579_ net436 net585 _06145_ net304 net2180 vssd1 vssd1 vccd1 vccd1 _00423_ sky130_fd_sc_hd__a32o_1
Xinput56 mem_adr_start[28] vssd1 vssd1 vccd1 vccd1 net56 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput67 mem_adr_start[9] vssd1 vssd1 vccd1 vccd1 net67 sky130_fd_sc_hd__buf_1
Xhold807 final_design.cpu.reg_window\[887\] vssd1 vssd1 vccd1 vccd1 net2149 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput78 memory_size[19] vssd1 vssd1 vccd1 vccd1 net78 sky130_fd_sc_hd__buf_1
XANTENNA__07548__S net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput89 memory_size[29] vssd1 vssd1 vccd1 vccd1 net89 sky130_fd_sc_hd__clkbuf_2
X_13318_ clknet_leaf_51_clk _00549_ net1170 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[306\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11578__B net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold818 final_design.cpu.reg_window\[276\] vssd1 vssd1 vccd1 vccd1 net2160 sky130_fd_sc_hd__dlygate4sd3_1
Xhold829 final_design.cpu.reg_window\[376\] vssd1 vssd1 vccd1 vccd1 net2171 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13101__CLK clknet_leaf_45_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12026__Y _06261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1773 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13249_ clknet_leaf_49_clk _00480_ net1186 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[237\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11156__A1 net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12353__B1 net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_2670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07810_ _02757_ _02758_ _02759_ _02760_ net683 net693 vssd1 vssd1 vccd1 vccd1 _02761_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__13251__CLK clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08790_ _03685_ _03686_ vssd1 vssd1 vccd1 vccd1 _03741_ sky130_fd_sc_hd__nand2_1
XANTENNA__08379__S net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08309__C1 net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07741_ final_design.cpu.reg_window\[730\] final_design.cpu.reg_window\[762\] net861
+ vssd1 vssd1 vccd1 vccd1 _02692_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07672_ net713 _02616_ net723 vssd1 vssd1 vccd1 vccd1 _02623_ sky130_fd_sc_hd__o21a_1
XFILLER_0_75_1566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_1905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_2452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09411_ _04158_ _04163_ _02837_ vssd1 vssd1 vccd1 vccd1 _04330_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_66_2463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06623_ final_design.cpu.reg_window\[475\] final_design.cpu.reg_window\[507\] net943
+ vssd1 vssd1 vccd1 vccd1 _01574_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_66_2474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_2316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_17_clk clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_17_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_62_2327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12969__CLK clknet_leaf_15_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11533__S net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09342_ net473 _04260_ vssd1 vssd1 vccd1 vccd1 _04261_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_62_2338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08088__A1 _01718_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06554_ final_design.reqhand.instruction\[30\] final_design.data_from_mem\[30\] net972
+ vssd1 vssd1 vccd1 vccd1 _01505_ sky130_fd_sc_hd__mux2_2
XFILLER_0_74_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12926__Q net149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09273_ net83 net84 _04191_ vssd1 vssd1 vccd1 vccd1 _04192_ sky130_fd_sc_hd__or3_1
XFILLER_0_8_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06485_ net762 _01435_ vssd1 vssd1 vccd1 vccd1 _01436_ sky130_fd_sc_hd__or2_2
XFILLER_0_74_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout234_A _05983_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_519 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08224_ final_design.cpu.reg_window\[11\] final_design.cpu.reg_window\[43\] net835
+ vssd1 vssd1 vccd1 vccd1 _03175_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11919__B1 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08155_ final_design.cpu.reg_window\[335\] final_design.cpu.reg_window\[367\] net820
+ vssd1 vssd1 vccd1 vccd1 _03106_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout401_A _06257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12364__S net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_2109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1143_A net1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07106_ net757 _02056_ vssd1 vssd1 vccd1 vccd1 _02057_ sky130_fd_sc_hd__or2_1
XANTENNA__07458__S net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12592__B1 net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11488__B _06093_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08086_ _03035_ _03036_ _02901_ vssd1 vssd1 vccd1 vccd1 _03037_ sky130_fd_sc_hd__o21a_1
X_07037_ net750 _01987_ vssd1 vssd1 vccd1 vccd1 _01988_ sky130_fd_sc_hd__or2_1
XANTENNA__11147__A1 final_design.data_from_mem\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1835 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1029_X net1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12344__B1 net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08012__A1 net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11698__A2 net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout391_X net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout770_A net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout868_A net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08988_ net623 _03923_ vssd1 vssd1 vccd1 vccd1 _03924_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_3_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07939_ final_design.cpu.reg_window\[598\] final_design.cpu.reg_window\[630\] net839
+ vssd1 vssd1 vccd1 vccd1 _02890_ sky130_fd_sc_hd__mux2_1
XANTENNA__13744__CLK clknet_leaf_36_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12647__B2 final_design.data_from_mem\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout656_X net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10950_ net84 net1046 vssd1 vssd1 vccd1 vccd1 _05678_ sky130_fd_sc_hd__or2_1
XANTENNA__07206__B _01537_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07921__S net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09609_ _04513_ _04527_ vssd1 vssd1 vccd1 vccd1 _04528_ sky130_fd_sc_hd__nor2_1
XFILLER_0_79_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10881_ net81 _05589_ vssd1 vssd1 vccd1 vccd1 _05612_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout823_X net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11870__A2 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13894__CLK clknet_leaf_52_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1915 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12620_ net2423 final_design.reqhand.data_from_UART\[6\] _05080_ vssd1 vssd1 vccd1
+ vccd1 _01313_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12551_ _06214_ net357 net324 net2306 vssd1 vssd1 vccd1 vccd1 _01255_ sky130_fd_sc_hd__a22o_1
XANTENNA__11622__A2 net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11502_ net2020 net232 net521 vssd1 vssd1 vccd1 vccd1 _00371_ sky130_fd_sc_hd__mux2_1
X_12482_ _06142_ net351 net333 net2430 vssd1 vssd1 vccd1 vccd1 _01188_ sky130_fd_sc_hd__a22o_1
XANTENNA__13124__CLK clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14221_ net1279 vssd1 vssd1 vccd1 vccd1 gpio_oeb[33] sky130_fd_sc_hd__buf_2
X_11433_ net1978 net192 net313 vssd1 vssd1 vccd1 vccd1 _00330_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11386__B2 _01538_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14152_ clknet_leaf_14_clk _01326_ net1106 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.data_to_VGA\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_11364_ net650 net187 vssd1 vssd1 vccd1 vccd1 _06053_ sky130_fd_sc_hd__and2_1
XANTENNA__12987__RESET_B net1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10315_ net1478 net1012 net989 final_design.data_from_mem\[0\] vssd1 vssd1 vccd1
+ vccd1 _00072_ sky130_fd_sc_hd__a22o_1
X_13103_ clknet_leaf_43_clk _00334_ net1218 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[91\]
+ sky130_fd_sc_hd__dfrtp_1
X_14083_ clknet_leaf_20_clk _01280_ net1161 vssd1 vssd1 vccd1 vccd1 final_design.reqhand.instruction\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13274__CLK clknet_leaf_58_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11295_ net738 _03909_ vssd1 vssd1 vccd1 vccd1 _05992_ sky130_fd_sc_hd__nand2_1
XANTENNA__12335__B1 net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13034_ clknet_leaf_60_clk _00265_ net1140 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_10246_ final_design.uart.BAUD_counter\[15\] final_design.uart.BAUD_counter\[16\]
+ _05113_ final_design.uart.BAUD_counter\[17\] vssd1 vssd1 vccd1 vccd1 _05117_ sky130_fd_sc_hd__a31o_1
Xfanout1110 net1112 vssd1 vssd1 vccd1 vccd1 net1110 sky130_fd_sc_hd__clkbuf_4
Xfanout1121 net1127 vssd1 vssd1 vccd1 vccd1 net1121 sky130_fd_sc_hd__clkbuf_4
Xfanout1132 net1135 vssd1 vssd1 vccd1 vccd1 net1132 sky130_fd_sc_hd__clkbuf_4
X_10177_ final_design.uart.BAUD_counter\[21\] final_design.uart.BAUD_counter\[20\]
+ final_design.uart.BAUD_counter\[23\] final_design.uart.BAUD_counter\[22\] vssd1
+ vssd1 vccd1 vccd1 _05067_ sky130_fd_sc_hd__or4_1
XFILLER_0_59_1506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1143 net1150 vssd1 vssd1 vccd1 vccd1 net1143 sky130_fd_sc_hd__buf_2
XANTENNA__10361__A2 net1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1154 net1162 vssd1 vssd1 vccd1 vccd1 net1154 sky130_fd_sc_hd__clkbuf_4
Xfanout1165 net1166 vssd1 vssd1 vccd1 vccd1 net1165 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_59_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1176 net1192 vssd1 vssd1 vccd1 vccd1 net1176 sky130_fd_sc_hd__clkbuf_2
XANTENNA__06660__S1 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1187 net1191 vssd1 vssd1 vccd1 vccd1 net1187 sky130_fd_sc_hd__clkbuf_4
Xfanout1198 net1201 vssd1 vssd1 vccd1 vccd1 net1198 sky130_fd_sc_hd__clkbuf_4
X_13936_ clknet_leaf_34_clk _01167_ net1239 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[924\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11310__A1 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09612__A _04529_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10758__A net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12449__S net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13867_ clknet_leaf_53_clk _01098_ net1186 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[855\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11861__A2 _05965_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12818_ net1369 vssd1 vssd1 vccd1 vccd1 _00259_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__11580__C net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_2950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13798_ clknet_leaf_51_clk _01029_ net1175 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[786\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08228__A net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12749_ _06381_ _06383_ _06384_ _06387_ vssd1 vssd1 vccd1 vccd1 _01351_ sky130_fd_sc_hd__a31o_1
XANTENNA__09282__A3 net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09019__B1 net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_1857 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10493__A net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12184__S net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11377__A1 final_design.data_from_mem\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13617__CLK clknet_leaf_34_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07278__S net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_74_2721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold604 final_design.cpu.reg_window\[383\] vssd1 vssd1 vccd1 vccd1 net1946 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06479__S1 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold615 final_design.cpu.reg_window\[923\] vssd1 vssd1 vccd1 vccd1 net1957 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold626 final_design.cpu.reg_window\[946\] vssd1 vssd1 vccd1 vccd1 net1968 sky130_fd_sc_hd__dlygate4sd3_1
Xhold637 final_design.cpu.reg_window\[772\] vssd1 vssd1 vccd1 vccd1 net1979 sky130_fd_sc_hd__dlygate4sd3_1
Xhold648 final_design.cpu.reg_window\[495\] vssd1 vssd1 vccd1 vccd1 net1990 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_70_2607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold659 final_design.cpu.reg_window\[513\] vssd1 vssd1 vccd1 vccd1 net2001 sky130_fd_sc_hd__dlygate4sd3_1
X_09960_ _04871_ _04876_ _04878_ vssd1 vssd1 vccd1 vccd1 _04879_ sky130_fd_sc_hd__a21oi_1
Xclkbuf_leaf_6_clk clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_6_clk sky130_fd_sc_hd__clkbuf_8
X_08911_ net2541 net1014 _03851_ _03855_ vssd1 vssd1 vccd1 vccd1 _00236_ sky130_fd_sc_hd__a22o_1
XANTENNA__13767__CLK clknet_leaf_62_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09891_ _04147_ _04809_ net447 vssd1 vssd1 vccd1 vccd1 _04810_ sky130_fd_sc_hd__a21o_1
XANTENNA__11528__S net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload19_A clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10888__B1 net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08842_ final_design.CPU_instr_adr\[17\] _03792_ vssd1 vssd1 vccd1 vccd1 _03793_
+ sky130_fd_sc_hd__and2_1
XANTENNA__10352__A2 net1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_2514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08773_ _03701_ _03722_ _03700_ vssd1 vssd1 vccd1 vccd1 _03724_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_68_2525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_2536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout184_A _06060_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07724_ final_design.cpu.reg_window\[346\] final_design.cpu.reg_window\[378\] net863
+ vssd1 vssd1 vccd1 vccd1 _02675_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11301__A1 net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08702__C1 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07655_ _01567_ _02604_ vssd1 vssd1 vccd1 vccd1 _02606_ sky130_fd_sc_hd__nand2_1
XANTENNA__07600__S0 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout351_A net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11852__A2 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1093_A net1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06606_ final_design.cpu.reg_window\[924\] final_design.cpu.reg_window\[956\] net946
+ vssd1 vssd1 vccd1 vccd1 _01557_ sky130_fd_sc_hd__mux2_1
X_07586_ final_design.cpu.reg_window\[927\] final_design.cpu.reg_window\[959\] net867
+ vssd1 vssd1 vccd1 vccd1 _02537_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09325_ net261 _04217_ _04230_ vssd1 vssd1 vccd1 vccd1 _04244_ sky130_fd_sc_hd__and3_1
X_06537_ _01456_ _01465_ net880 _01481_ vssd1 vssd1 vccd1 vccd1 _01488_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_48_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_1667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09256_ _02638_ _04173_ _02545_ vssd1 vssd1 vccd1 vccd1 _04175_ sky130_fd_sc_hd__a21boi_1
X_06468_ final_design.data_from_mem\[17\] net969 _01417_ vssd1 vssd1 vccd1 vccd1 _01419_
+ sky130_fd_sc_hd__o21ai_4
XFILLER_0_1_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08207_ _03154_ _03155_ _03156_ _03157_ net675 net691 vssd1 vssd1 vccd1 vccd1 _03158_
+ sky130_fd_sc_hd__mux4_1
X_09187_ net462 _04104_ _04105_ _04098_ net473 vssd1 vssd1 vccd1 vccd1 _04106_ sky130_fd_sc_hd__o2111a_1
XANTENNA__13297__CLK clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout404_X net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11368__A1 final_design.data_from_mem\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08138_ _03085_ _03086_ _03087_ _03088_ net684 net703 vssd1 vssd1 vccd1 vccd1 _03089_
+ sky130_fd_sc_hd__mux4_1
X_08069_ _03016_ _03017_ _03018_ _03019_ net682 net693 vssd1 vssd1 vccd1 vccd1 _03020_
+ sky130_fd_sc_hd__mux4_1
X_10100_ _05015_ vssd1 vssd1 vccd1 vccd1 _05016_ sky130_fd_sc_hd__inv_2
X_11080_ net1047 net91 vssd1 vssd1 vccd1 vccd1 _05802_ sky130_fd_sc_hd__and2b_1
XFILLER_0_41_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout773_X net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11438__S net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08536__A2 _03481_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10031_ _04047_ _04949_ _04948_ _04947_ vssd1 vssd1 vccd1 vccd1 _04950_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_8_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10343__A2 net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1097 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout940_X net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11982_ _06184_ net291 net406 net2137 vssd1 vssd1 vccd1 vccd1 _00715_ sky130_fd_sc_hd__a22o_1
XANTENNA__09497__B1 _04415_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1403 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11681__B net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13721_ clknet_leaf_56_clk _00952_ net1147 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[709\]
+ sky130_fd_sc_hd__dfrtp_1
X_10933_ _05649_ _05658_ _05661_ _01386_ vssd1 vssd1 vccd1 vccd1 _05662_ sky130_fd_sc_hd__o31a_1
XFILLER_0_19_1578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09151__B _04053_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10864_ net956 _05585_ _05595_ net959 vssd1 vssd1 vccd1 vccd1 _05596_ sky130_fd_sc_hd__o22a_1
X_13652_ clknet_leaf_10_clk _00883_ net1153 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[640\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_71_1761 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14072__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12603_ net1400 net996 net982 final_design.data_from_mem\[21\] vssd1 vssd1 vccd1
+ vccd1 _01296_ sky130_fd_sc_hd__a22o_1
X_10795_ _05528_ _05529_ _05511_ vssd1 vssd1 vccd1 vccd1 _05530_ sky130_fd_sc_hd__o21ba_1
X_13583_ clknet_leaf_42_clk _00814_ net1218 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[571\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11901__S net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12534_ _06197_ net346 net323 net2231 vssd1 vssd1 vccd1 vccd1 _01238_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_26_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12465_ net671 net635 _06268_ net330 net2081 vssd1 vssd1 vccd1 vccd1 _01171_ sky130_fd_sc_hd__a32o_1
XANTENNA__12556__B1 net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07098__S net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14204_ net1262 vssd1 vssd1 vccd1 vccd1 gpio_oeb[16] sky130_fd_sc_hd__buf_2
X_11416_ net2162 net237 net310 vssd1 vssd1 vccd1 vccd1 _00313_ sky130_fd_sc_hd__mux2_1
X_12396_ net553 net508 vssd1 vssd1 vccd1 vccd1 _06279_ sky130_fd_sc_hd__nand2_1
XANTENNA__12020__A2 net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10031__A1 _04047_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14135_ clknet_leaf_17_clk final_design.vga.h_next_count\[4\] net1113 vssd1 vssd1
+ vccd1 vccd1 final_design.VGA_data_control.h_count\[4\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11347_ _06034_ _06036_ _06037_ net589 vssd1 vssd1 vccd1 vccd1 _06038_ sky130_fd_sc_hd__o211a_2
XFILLER_0_39_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06730__S net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11856__B net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11278_ final_design.data_from_mem\[16\] _05177_ _05912_ _05917_ vssd1 vssd1 vccd1
+ vccd1 _05977_ sky130_fd_sc_hd__a31o_2
X_14066_ clknet_leaf_15_clk _00029_ net1093 vssd1 vssd1 vccd1 vccd1 final_design.uart.BAUD_counter\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_10229_ net2394 _05104_ _05106_ vssd1 vssd1 vccd1 vccd1 _00007_ sky130_fd_sc_hd__a21oi_1
X_13017_ clknet_leaf_56_clk _00248_ net1146 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10334__A2 net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07735__B1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07127__A net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1 wb_manage.BUSY_O vssd1 vssd1 vccd1 vccd1 net1343 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12087__A2 _06046_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10098__A1 net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13919_ clknet_leaf_4_clk _01150_ net1084 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[907\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10488__A net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12179__S net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07440_ _01489_ net731 _01495_ net681 vssd1 vssd1 vccd1 vccd1 _02391_ sky130_fd_sc_hd__a31o_1
XPHY_EDGE_ROW_8_Right_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08138__S1 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07371_ final_design.cpu.reg_window\[515\] final_design.cpu.reg_window\[547\] net906
+ vssd1 vssd1 vccd1 vccd1 _02322_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09110_ _04030_ final_design.CPU_instr_adr\[1\] _03812_ vssd1 vssd1 vccd1 vccd1 _00210_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__11811__S net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_21_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_1889 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08392__S net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_2805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09041_ _03730_ _03970_ vssd1 vssd1 vccd1 vccd1 _03971_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_76_2816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12547__B1 net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12011__A2 net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold401 final_design.cpu.reg_window\[145\] vssd1 vssd1 vccd1 vccd1 net1743 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07649__S0 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold412 final_design.cpu.reg_window\[835\] vssd1 vssd1 vccd1 vccd1 net1754 sky130_fd_sc_hd__dlygate4sd3_1
Xhold423 final_design.cpu.reg_window\[778\] vssd1 vssd1 vccd1 vccd1 net1765 sky130_fd_sc_hd__dlygate4sd3_1
Xhold434 final_design.uart.BAUD_counter\[16\] vssd1 vssd1 vccd1 vccd1 net1776 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold445 final_design.cpu.reg_window\[782\] vssd1 vssd1 vccd1 vccd1 net1787 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold456 final_design.cpu.reg_window\[991\] vssd1 vssd1 vccd1 vccd1 net1798 sky130_fd_sc_hd__dlygate4sd3_1
Xhold467 final_design.cpu.reg_window\[785\] vssd1 vssd1 vccd1 vccd1 net1809 sky130_fd_sc_hd__dlygate4sd3_1
Xhold478 final_design.cpu.reg_window\[587\] vssd1 vssd1 vccd1 vccd1 net1820 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_1903 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09943_ _03390_ _03421_ _04149_ net447 vssd1 vssd1 vccd1 vccd1 _04862_ sky130_fd_sc_hd__a31o_1
Xhold489 final_design.cpu.reg_window\[746\] vssd1 vssd1 vccd1 vccd1 net1831 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout903 net904 vssd1 vssd1 vccd1 vccd1 net903 sky130_fd_sc_hd__clkbuf_2
Xfanout914 net917 vssd1 vssd1 vccd1 vccd1 net914 sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_39_Right_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout925 net926 vssd1 vssd1 vccd1 vccd1 net925 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout399_A _06261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout936 net952 vssd1 vssd1 vccd1 vccd1 net936 sky130_fd_sc_hd__buf_2
X_09874_ _04460_ _04465_ _04727_ _04461_ _04222_ vssd1 vssd1 vccd1 vccd1 _04793_ sky130_fd_sc_hd__o32a_1
Xfanout947 net951 vssd1 vssd1 vccd1 vccd1 net947 sky130_fd_sc_hd__clkbuf_4
Xfanout958 _04041_ vssd1 vssd1 vccd1 vccd1 net958 sky130_fd_sc_hd__clkbuf_4
Xhold1101 final_design.cpu.reg_window\[546\] vssd1 vssd1 vccd1 vccd1 net2443 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout969 net970 vssd1 vssd1 vccd1 vccd1 net969 sky130_fd_sc_hd__buf_4
XANTENNA__07037__A net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09804__X _04723_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1112 final_design.cpu.reg_window\[544\] vssd1 vssd1 vccd1 vccd1 net2454 sky130_fd_sc_hd__dlygate4sd3_1
X_08825_ final_design.CPU_instr_adr\[28\] _01570_ _03775_ vssd1 vssd1 vccd1 vccd1
+ _03776_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_13_Left_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1123 final_design.cpu.reg_window\[637\] vssd1 vssd1 vccd1 vccd1 net2465 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1134 final_design.cpu.reg_window\[307\] vssd1 vssd1 vccd1 vccd1 net2476 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout187_X net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout566_A net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1145 final_design.cpu.reg_window\[316\] vssd1 vssd1 vccd1 vccd1 net2487 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1156 final_design.cpu.reg_window\[428\] vssd1 vssd1 vccd1 vccd1 net2498 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1167 final_design.cpu.reg_window\[426\] vssd1 vssd1 vccd1 vccd1 net2509 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1178 final_design.cpu.reg_window\[290\] vssd1 vssd1 vccd1 vccd1 net2520 sky130_fd_sc_hd__dlygate4sd3_1
X_08756_ _01366_ _02297_ vssd1 vssd1 vccd1 vccd1 _03707_ sky130_fd_sc_hd__and2_1
Xhold1189 final_design.cpu.reg_window\[164\] vssd1 vssd1 vccd1 vccd1 net2531 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14095__CLK clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07707_ final_design.cpu.reg_window\[731\] final_design.cpu.reg_window\[763\] net861
+ vssd1 vssd1 vccd1 vccd1 _02658_ sky130_fd_sc_hd__mux2_1
XANTENNA__11286__B1 net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout733_A _01491_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10398__A net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08687_ _03456_ _03457_ vssd1 vssd1 vccd1 vccd1 _03638_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout354_X net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1096_X net1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07638_ net719 _02588_ vssd1 vssd1 vccd1 vccd1 _02589_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_0_197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1188 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_48_Right_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout900_A net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout521_X net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07569_ _02516_ _02517_ _02518_ _02519_ net685 net706 vssd1 vssd1 vccd1 vccd1 _02520_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__11589__A1 net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09308_ net527 net492 vssd1 vssd1 vccd1 vccd1 _04227_ sky130_fd_sc_hd__nand2_1
X_10580_ net64 _05324_ vssd1 vssd1 vccd1 vccd1 _05326_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_64_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_7_clk_X clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13932__CLK clknet_leaf_46_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09239_ _02936_ _04135_ _04143_ _04157_ vssd1 vssd1 vccd1 vccd1 _04158_ sky130_fd_sc_hd__or4_4
XFILLER_0_1_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12538__B1 net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12250_ net567 _06179_ net506 net373 net1499 vssd1 vssd1 vccd1 vccd1 _00966_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_40_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout890_X net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout988_X net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10013__A1 net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11201_ _05855_ _05906_ _05908_ net653 vssd1 vssd1 vccd1 vccd1 _05909_ sky130_fd_sc_hd__a211o_1
XANTENNA__11957__A net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12181_ net1763 net203 net382 vssd1 vssd1 vccd1 vccd1 _00900_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_57_Right_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11132_ _05840_ _05846_ vssd1 vssd1 vccd1 vccd1 _05847_ sky130_fd_sc_hd__nor2_4
XANTENNA__06550__S net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold990 final_design.cpu.reg_window\[288\] vssd1 vssd1 vccd1 vccd1 net2332 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11168__S net247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11063_ final_design.CPU_instr_adr\[29\] _01371_ net802 vssd1 vssd1 vccd1 vccd1 _05786_
+ sky130_fd_sc_hd__a21o_1
XANTENNA__10316__A2 net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11513__A1 net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10014_ net489 _04779_ _04341_ vssd1 vssd1 vccd1 vccd1 _04933_ sky130_fd_sc_hd__a21o_1
XANTENNA__08914__C1 net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13312__CLK clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_3009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10800__S net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12069__A2 _05911_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06786__A net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07234__X _02185_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08368__S1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11965_ _06167_ net276 net404 net1704 vssd1 vssd1 vccd1 vccd1 _00698_ sky130_fd_sc_hd__a22o_1
XFILLER_0_58_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_66_Right_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13462__CLK clknet_leaf_59_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13704_ clknet_leaf_40_clk _00935_ net1220 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[692\]
+ sky130_fd_sc_hd__dfrtp_1
X_10916_ net49 _05620_ _05625_ vssd1 vssd1 vccd1 vccd1 _05646_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_15_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11896_ net215 net2507 net273 vssd1 vssd1 vccd1 vccd1 _00638_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_15_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13635_ clknet_leaf_0_clk _00866_ net1061 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[623\]
+ sky130_fd_sc_hd__dfrtp_1
X_10847_ _05579_ vssd1 vssd1 vccd1 vccd1 _05580_ sky130_fd_sc_hd__inv_2
XFILLER_0_82_742 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06725__S net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13566_ clknet_leaf_13_clk _00797_ net1089 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[554\]
+ sky130_fd_sc_hd__dfrtp_1
X_10778_ _05487_ _05489_ _05513_ vssd1 vssd1 vccd1 vccd1 _05514_ sky130_fd_sc_hd__o21bai_1
XANTENNA__09101__S net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12517_ _06179_ net347 net327 net1759 vssd1 vssd1 vccd1 vccd1 _01222_ sky130_fd_sc_hd__a22o_1
XFILLER_0_67_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13497_ clknet_leaf_56_clk _00728_ net1146 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[485\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12529__B1 net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12448_ net1663 net222 net335 vssd1 vssd1 vccd1 vccd1 _01155_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_75_Right_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11201__B1 _05908_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12462__S net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12379_ net1553 net206 net268 vssd1 vssd1 vccd1 vccd1 _01090_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_268 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14118_ clknet_leaf_17_clk final_design.vga.h_next_state\[0\] net1113 vssd1 vssd1
+ vccd1 vccd1 final_design.vga.h_current_state\[0\] sky130_fd_sc_hd__dfrtp_2
XANTENNA__11586__B net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06940_ final_design.cpu.reg_window\[17\] final_design.cpu.reg_window\[49\] net930
+ vssd1 vssd1 vccd1 vccd1 _01891_ sky130_fd_sc_hd__mux2_1
X_14049_ clknet_leaf_16_clk _00010_ net1094 vssd1 vssd1 vccd1 vccd1 final_design.uart.BAUD_counter\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_78_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11504__A1 net242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1745 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06871_ net742 _01498_ _01819_ _01821_ vssd1 vssd1 vccd1 vccd1 _01822_ sky130_fd_sc_hd__o211a_1
XFILLER_0_59_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08610_ _03455_ _03557_ _03560_ _03457_ vssd1 vssd1 vccd1 vccd1 _03561_ sky130_fd_sc_hd__o31a_1
XFILLER_0_78_1789 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09590_ _04502_ _04508_ vssd1 vssd1 vccd1 vccd1 _04509_ sky130_fd_sc_hd__nand2_4
XANTENNA__13805__CLK clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10489__Y _05239_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07144__X _02095_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11268__B1 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08541_ final_design.cpu.reg_window\[385\] final_design.cpu.reg_window\[417\] net838
+ vssd1 vssd1 vccd1 vccd1 _03492_ sky130_fd_sc_hd__mux2_1
XANTENNA__11807__A2 net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08133__B1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08472_ _03420_ _03422_ vssd1 vssd1 vccd1 vccd1 _03423_ sky130_fd_sc_hd__nor2_1
XANTENNA__12480__A2 net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09881__B1 net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07423_ _02370_ _02371_ _02372_ _02373_ net769 net790 vssd1 vssd1 vccd1 vccd1 _02374_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__10491__A1 net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13955__CLK clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10491__B2 _04042_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10946__A _04918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09859__S1 net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12787__18 clknet_leaf_27_clk vssd1 vssd1 vccd1 vccd1 net1328 sky130_fd_sc_hd__inv_2
X_07354_ _02301_ _02302_ _02303_ _02304_ net769 net790 vssd1 vssd1 vccd1 vccd1 _02305_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__06635__S net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07285_ final_design.cpu.reg_window\[646\] final_design.cpu.reg_window\[678\] net902
+ vssd1 vssd1 vccd1 vccd1 _02236_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout314_A net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09024_ net620 _03955_ _03954_ net259 vssd1 vssd1 vccd1 vccd1 _03956_ sky130_fd_sc_hd__a211o_1
XFILLER_0_66_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold220 final_design.cpu.reg_window\[836\] vssd1 vssd1 vccd1 vccd1 net1562 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12372__S net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold231 final_design.cpu.reg_window\[972\] vssd1 vssd1 vccd1 vccd1 net1573 sky130_fd_sc_hd__dlygate4sd3_1
Xhold242 net137 vssd1 vssd1 vccd1 vccd1 net1584 sky130_fd_sc_hd__dlygate4sd3_1
Xhold253 final_design.cpu.reg_window\[251\] vssd1 vssd1 vccd1 vccd1 net1595 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold264 final_design.cpu.reg_window\[374\] vssd1 vssd1 vccd1 vccd1 net1606 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13335__CLK clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold275 final_design.cpu.reg_window\[169\] vssd1 vssd1 vccd1 vccd1 net1617 sky130_fd_sc_hd__dlygate4sd3_1
Xhold286 final_design.VGA_data_control.ready_data\[25\] vssd1 vssd1 vccd1 vccd1 net1628
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout683_A net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout700 net701 vssd1 vssd1 vccd1 vccd1 net700 sky130_fd_sc_hd__clkbuf_4
Xhold297 final_design.cpu.reg_window\[702\] vssd1 vssd1 vccd1 vccd1 net1639 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout711 net713 vssd1 vssd1 vccd1 vccd1 net711 sky130_fd_sc_hd__clkbuf_4
Xfanout722 net724 vssd1 vssd1 vccd1 vccd1 net722 sky130_fd_sc_hd__buf_4
X_09926_ _04124_ _04718_ _04844_ vssd1 vssd1 vccd1 vccd1 _04845_ sky130_fd_sc_hd__or3_1
XANTENNA_fanout1011_X net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout733 _01491_ vssd1 vssd1 vccd1 vccd1 net733 sky130_fd_sc_hd__clkbuf_4
Xfanout744 _01476_ vssd1 vssd1 vccd1 vccd1 net744 sky130_fd_sc_hd__clkbuf_4
Xfanout755 net756 vssd1 vssd1 vccd1 vccd1 net755 sky130_fd_sc_hd__buf_2
Xfanout766 net771 vssd1 vssd1 vccd1 vccd1 net766 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout850_A net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09857_ _03292_ net441 net438 _03291_ vssd1 vssd1 vccd1 vccd1 _04776_ sky130_fd_sc_hd__o22a_1
Xfanout777 net778 vssd1 vssd1 vccd1 vccd1 net777 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_77_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout788 _01418_ vssd1 vssd1 vccd1 vccd1 net788 sky130_fd_sc_hd__buf_2
XANTENNA__07175__A1 net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout799 net800 vssd1 vssd1 vccd1 vccd1 net799 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout569_X net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout948_A net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13485__CLK clknet_leaf_44_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08808_ _03757_ _03758_ vssd1 vssd1 vccd1 vccd1 _03759_ sky130_fd_sc_hd__and2_1
XFILLER_0_38_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09788_ _03358_ _04705_ vssd1 vssd1 vccd1 vccd1 _04707_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_77_1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08739_ final_design.CPU_instr_adr\[10\] _02128_ vssd1 vssd1 vccd1 vccd1 _03690_
+ sky130_fd_sc_hd__and2_1
XANTENNA_fanout736_X net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11750_ net207 net1950 net416 vssd1 vssd1 vccd1 vccd1 _00513_ sky130_fd_sc_hd__mux2_1
XANTENNA__08675__A1 _02061_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12471__A2 net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09872__B1 net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10701_ _05404_ _05439_ _05440_ vssd1 vssd1 vccd1 vccd1 _05441_ sky130_fd_sc_hd__o21ai_2
XANTENNA__10482__B2 net1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11681_ net224 net627 vssd1 vssd1 vccd1 vccd1 _06199_ sky130_fd_sc_hd__and2_1
XANTENNA__11451__S net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_46_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_46_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13420_ clknet_leaf_45_clk _00651_ net1215 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[408\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_23_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10632_ _05372_ _05374_ vssd1 vssd1 vccd1 vccd1 _05375_ sky130_fd_sc_hd__nor2_1
XFILLER_0_14_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_42_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_42_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10563_ _05268_ _05305_ _05307_ _05302_ vssd1 vssd1 vccd1 vccd1 _05309_ sky130_fd_sc_hd__a211o_1
X_13351_ clknet_leaf_58_clk _00582_ net1125 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[339\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14192__1251 vssd1 vssd1 vccd1 vccd1 _14192__1251/HI net1251 sky130_fd_sc_hd__conb_1
XANTENNA__14110__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12302_ net1694 net224 net365 vssd1 vssd1 vccd1 vccd1 _01016_ sky130_fd_sc_hd__mux2_1
XANTENNA_input77_A memory_size[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10494_ net58 _05234_ _05242_ _05243_ vssd1 vssd1 vccd1 vccd1 _05244_ sky130_fd_sc_hd__and4_1
X_13282_ clknet_leaf_10_clk _00513_ net1101 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[270\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11687__A net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12233_ net565 _06163_ net516 net373 net1548 vssd1 vssd1 vccd1 vccd1 _00950_ sky130_fd_sc_hd__a32o_1
XANTENNA__08286__S0 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11734__A1 net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12164_ net1771 net230 net380 vssd1 vssd1 vccd1 vccd1 _00883_ sky130_fd_sc_hd__mux2_1
XANTENNA__08699__C net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11115_ final_design.uart.bits_received\[1\] _05830_ _05831_ _05833_ vssd1 vssd1
+ vccd1 vccd1 _00206_ sky130_fd_sc_hd__a22o_1
XANTENNA__13548__RESET_B net1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08038__S0 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12095_ net1659 net230 net388 vssd1 vssd1 vccd1 vccd1 _00819_ sky130_fd_sc_hd__mux2_1
XANTENNA__13828__CLK clknet_leaf_51_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input32_X net32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11046_ net959 _05767_ _05769_ net956 vssd1 vssd1 vccd1 vccd1 _05770_ sky130_fd_sc_hd__o22a_1
XFILLER_0_40_1877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12852__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09538__S0 net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13978__CLK clknet_leaf_58_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12997_ net1328 _00228_ net1195 vssd1 vssd1 vccd1 vccd1 final_design.CPU_instr_adr\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07013__S1 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11948_ _06149_ net293 net410 net1939 vssd1 vssd1 vccd1 vccd1 _00683_ sky130_fd_sc_hd__a22o_1
XFILLER_0_74_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12457__S net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13208__CLK clknet_leaf_65_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11879_ _06113_ net292 net519 net2470 vssd1 vssd1 vccd1 vccd1 _00623_ sky130_fd_sc_hd__a22o_1
XFILLER_0_12_1913 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11214__X _05921_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13618_ clknet_leaf_38_clk _00849_ net1189 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[606\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_1793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13549_ clknet_leaf_53_clk _00780_ net1185 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[537\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07070_ final_design.cpu.reg_window\[781\] final_design.cpu.reg_window\[813\] net935
+ vssd1 vssd1 vccd1 vccd1 _02021_ sky130_fd_sc_hd__mux2_1
XANTENNA__13358__CLK clknet_leaf_42_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10772__Y _05508_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1880 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12192__S net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07972_ final_design.cpu.reg_window\[721\] final_design.cpu.reg_window\[753\] net848
+ vssd1 vssd1 vccd1 vccd1 _02923_ sky130_fd_sc_hd__mux2_1
X_09711_ _04628_ _04629_ vssd1 vssd1 vccd1 vccd1 _04630_ sky130_fd_sc_hd__nor2_1
X_06923_ final_design.cpu.reg_window\[722\] final_design.cpu.reg_window\[754\] net925
+ vssd1 vssd1 vccd1 vccd1 _01874_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09642_ net486 _04559_ _04560_ _04262_ vssd1 vssd1 vccd1 vccd1 _04561_ sky130_fd_sc_hd__a22o_1
X_06854_ final_design.cpu.reg_window\[980\] final_design.cpu.reg_window\[1012\] net948
+ vssd1 vssd1 vccd1 vccd1 _01805_ sky130_fd_sc_hd__mux2_1
X_06785_ _01732_ _01733_ _01734_ _01735_ net770 net789 vssd1 vssd1 vccd1 vccd1 _01736_
+ sky130_fd_sc_hd__mux4_1
X_09573_ net496 net486 _04491_ _04409_ _04101_ vssd1 vssd1 vccd1 vccd1 _04492_ sky130_fd_sc_hd__o32a_1
XANTENNA_fanout264_A net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08524_ final_design.cpu.reg_window\[706\] final_design.cpu.reg_window\[738\] net832
+ vssd1 vssd1 vccd1 vccd1 _03475_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_19_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08201__S0 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09530__A net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08455_ final_design.cpu.reg_window\[964\] final_design.cpu.reg_window\[996\] net819
+ vssd1 vssd1 vccd1 vccd1 _03406_ sky130_fd_sc_hd__mux2_1
XANTENNA__12367__S net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10676__A net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout431_A _05847_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14133__CLK clknet_leaf_18_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout529_A _02294_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07406_ final_design.reqhand.instruction\[9\] net972 vssd1 vssd1 vccd1 vccd1 _02357_
+ sky130_fd_sc_hd__or2_1
X_08386_ final_design.cpu.reg_window\[134\] final_design.cpu.reg_window\[166\] net823
+ vssd1 vssd1 vccd1 vccd1 _03337_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_1579 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08146__A net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07050__A _01996_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07337_ final_design.cpu.reg_window\[708\] final_design.cpu.reg_window\[740\] net900
+ vssd1 vssd1 vccd1 vccd1 _02288_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout317_X net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1059_X net1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07268_ final_design.cpu.reg_window\[390\] final_design.cpu.reg_window\[422\] net904
+ vssd1 vssd1 vccd1 vccd1 _02219_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout898_A net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09007_ _02451_ net620 _03937_ vssd1 vssd1 vccd1 vccd1 _03941_ sky130_fd_sc_hd__or3_1
X_07199_ final_design.cpu.reg_window\[521\] final_design.cpu.reg_window\[553\] net889
+ vssd1 vssd1 vccd1 vccd1 _02150_ sky130_fd_sc_hd__mux2_1
XANTENNA__11716__A1 net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11300__A net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12774__5 clknet_leaf_25_clk vssd1 vssd1 vccd1 vccd1 net1315 sky130_fd_sc_hd__inv_2
XANTENNA_fanout686_X net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout530 net531 vssd1 vssd1 vccd1 vccd1 net530 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_50_1904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12875__CLK clknet_leaf_17_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09909_ _04806_ _04807_ _04827_ vssd1 vssd1 vccd1 vccd1 _04828_ sky130_fd_sc_hd__and3_1
Xfanout552 _01686_ vssd1 vssd1 vccd1 vccd1 net552 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_50_1926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout563 net564 vssd1 vssd1 vccd1 vccd1 net563 sky130_fd_sc_hd__buf_2
Xfanout574 net576 vssd1 vssd1 vccd1 vccd1 net574 sky130_fd_sc_hd__clkbuf_4
Xfanout585 net586 vssd1 vssd1 vccd1 vccd1 net585 sky130_fd_sc_hd__buf_2
X_12920_ clknet_leaf_61_clk _00158_ net1136 vssd1 vssd1 vccd1 vccd1 net142 sky130_fd_sc_hd__dfrtp_1
Xfanout596 net601 vssd1 vssd1 vccd1 vccd1 net596 sky130_fd_sc_hd__buf_2
XFILLER_0_77_1052 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12851_ clknet_leaf_14_clk _00089_ net1110 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.ready_data\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_17_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11802_ net2376 net415 net293 _06039_ vssd1 vssd1 vccd1 vccd1 _00555_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_29_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_44_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10455__B2 net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11652__B1 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11733_ net176 net628 vssd1 vssd1 vccd1 vccd1 _06225_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_44_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11664_ net436 net584 _06189_ net300 net1692 vssd1 vssd1 vccd1 vccd1 _00464_ sky130_fd_sc_hd__a32o_1
XFILLER_0_37_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13500__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13403_ clknet_leaf_0_clk _00634_ net1071 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[391\]
+ sky130_fd_sc_hd__dfrtp_1
X_10615_ net964 _05358_ vssd1 vssd1 vccd1 vccd1 _05359_ sky130_fd_sc_hd__nand2_1
XFILLER_0_68_1733 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11595_ net435 net586 _06153_ net304 net1878 vssd1 vssd1 vccd1 vccd1 _00431_ sky130_fd_sc_hd__a32o_1
XANTENNA__10302__S1 net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11955__A1 _06156_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13334_ clknet_leaf_59_clk _00565_ net1142 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[322\]
+ sky130_fd_sc_hd__dfrtp_1
X_10546_ _05273_ _05292_ vssd1 vssd1 vccd1 vccd1 _05293_ sky130_fd_sc_hd__nor2_1
XFILLER_0_68_1777 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08490__S net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13265_ clknet_leaf_34_clk _00496_ net1242 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[253\]
+ sky130_fd_sc_hd__dfrtp_1
X_10477_ _05223_ _05225_ _05227_ net47 vssd1 vssd1 vccd1 vccd1 _05228_ sky130_fd_sc_hd__a31o_1
XANTENNA__13650__CLK clknet_leaf_38_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12216_ net567 _06144_ net505 net376 net1657 vssd1 vssd1 vccd1 vccd1 _00934_ sky130_fd_sc_hd__a32o_1
X_13196_ clknet_leaf_45_clk _00427_ net1213 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[184\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12147_ net203 net2367 net387 vssd1 vssd1 vccd1 vccd1 _00868_ sky130_fd_sc_hd__mux2_1
XANTENNA__14006__CLK clknet_leaf_59_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12078_ net573 _05981_ net508 net395 net1601 vssd1 vssd1 vccd1 vccd1 _00803_ sky130_fd_sc_hd__a32o_1
XFILLER_0_79_1873 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11029_ _05752_ vssd1 vssd1 vccd1 vccd1 _05753_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08431__S0 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09902__X _04821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06898__B1 net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_56_Left_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13030__CLK clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14156__CLK clknet_leaf_18_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06570_ net761 _01520_ vssd1 vssd1 vccd1 vccd1 _01521_ sky130_fd_sc_hd__or2_1
XFILLER_0_75_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12187__S net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_2380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_2391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08240_ _03185_ _03190_ net709 vssd1 vssd1 vccd1 vccd1 _03191_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_60_2244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_60_2255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13180__CLK clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_15 _04870_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_2266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12199__A1 net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_26 _06257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08171_ _03118_ _03119_ _03120_ _03121_ net676 net696 vssd1 vssd1 vccd1 vccd1 _03122_
+ sky130_fd_sc_hd__mux4_1
X_07122_ final_design.cpu.reg_window\[75\] final_design.cpu.reg_window\[107\] net916
+ vssd1 vssd1 vccd1 vccd1 _02073_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_65_Left_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07053_ final_design.cpu.reg_window\[269\] final_design.cpu.reg_window\[301\] net930
+ vssd1 vssd1 vccd1 vccd1 _02004_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_47_clk_X clknet_leaf_47_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_2173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput111 net111 vssd1 vssd1 vccd1 vccd1 ADR_O[19] sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_58_2184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput122 net122 vssd1 vssd1 vccd1 vccd1 ADR_O[29] sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_58_2195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput133 net133 vssd1 vssd1 vccd1 vccd1 CYC_O sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_54_2037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12898__CLK clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_2048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput144 net144 vssd1 vssd1 vccd1 vccd1 DAT_O[19] sky130_fd_sc_hd__buf_2
Xoutput155 net155 vssd1 vssd1 vccd1 vccd1 DAT_O[29] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_2059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput166 net166 vssd1 vssd1 vccd1 vccd1 SEL_O[0] sky130_fd_sc_hd__buf_2
XANTENNA__12371__A1 net244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10382__B1 net1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1019_A _06298_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11774__B net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07955_ final_design.cpu.reg_window\[337\] final_design.cpu.reg_window\[369\] net848
+ vssd1 vssd1 vccd1 vccd1 _02906_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout381_A net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06868__B net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1913 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06906_ final_design.cpu.reg_window\[338\] final_design.cpu.reg_window\[370\] net924
+ vssd1 vssd1 vccd1 vccd1 _01857_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07225__S1 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07886_ _02836_ vssd1 vssd1 vccd1 vccd1 _02837_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_74_Left_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11331__C1 net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14191__1250 vssd1 vssd1 vccd1 vccd1 _14191__1250/HI net1250 sky130_fd_sc_hd__conb_1
X_09625_ _02900_ _04353_ _03038_ vssd1 vssd1 vccd1 vccd1 _04544_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11882__B1 net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06837_ _01477_ net681 _01504_ vssd1 vssd1 vccd1 vccd1 _01788_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_74_1247 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout646_A net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout267_X net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06984__S0 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09556_ net76 _04187_ vssd1 vssd1 vccd1 vccd1 _04475_ sky130_fd_sc_hd__xor2_1
X_06768_ final_design.reqhand.instruction\[23\] net971 vssd1 vssd1 vccd1 vccd1 _01719_
+ sky130_fd_sc_hd__or2_1
XANTENNA__12426__A2 net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13523__CLK clknet_leaf_39_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08507_ final_design.cpu.reg_window\[322\] final_design.cpu.reg_window\[354\] net838
+ vssd1 vssd1 vccd1 vccd1 _03458_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12097__S net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11634__B1 net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06699_ net755 _01649_ vssd1 vssd1 vccd1 vccd1 _01650_ sky130_fd_sc_hd__or2_1
X_09487_ _04404_ _04405_ vssd1 vssd1 vccd1 vccd1 _04406_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout434_X net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1176_X net1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08438_ net597 _03384_ _03360_ net530 vssd1 vssd1 vccd1 vccd1 _03389_ sky130_fd_sc_hd__o211a_1
XFILLER_0_34_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08369_ _03314_ _03319_ net707 vssd1 vssd1 vccd1 vccd1 _03320_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout601_X net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1887 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13673__CLK clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07919__S net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10400_ _03513_ _05181_ vssd1 vssd1 vccd1 vccd1 _05183_ sky130_fd_sc_hd__nor2_1
XFILLER_0_65_1917 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11380_ _06063_ _06065_ _06066_ net589 vssd1 vssd1 vccd1 vccd1 _06067_ sky130_fd_sc_hd__o211a_1
XANTENNA__07161__S0 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10331_ net1519 net1011 net988 final_design.data_from_mem\[16\] vssd1 vssd1 vccd1
+ vccd1 _00088_ sky130_fd_sc_hd__a22o_1
XFILLER_0_15_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10262_ final_design.uart.BAUD_counter\[21\] final_design.uart.BAUD_counter\[22\]
+ _05123_ final_design.uart.BAUD_counter\[23\] vssd1 vssd1 vccd1 vccd1 _05127_ sky130_fd_sc_hd__a31o_1
XANTENNA__14029__CLK clknet_leaf_48_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13050_ clknet_leaf_5_clk _00281_ net1082 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[38\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_1603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout970_X net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1051 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14114__Q final_design.reqhand.data_from_UART\[4\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_12001_ _06203_ net276 net400 net2008 vssd1 vssd1 vccd1 vccd1 _00732_ sky130_fd_sc_hd__a22o_1
XANTENNA__12362__B2 _06090_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10193_ final_design.uart.bits_received\[0\] final_design.uart.bits_received\[1\]
+ vssd1 vssd1 vccd1 vccd1 _05082_ sky130_fd_sc_hd__or2_1
XANTENNA__10373__B1 net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout360 net361 vssd1 vssd1 vccd1 vccd1 net360 sky130_fd_sc_hd__buf_4
XANTENNA__13053__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout371 _06274_ vssd1 vssd1 vccd1 vccd1 net371 sky130_fd_sc_hd__clkbuf_4
XANTENNA__14179__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout382 net383 vssd1 vssd1 vccd1 vccd1 net382 sky130_fd_sc_hd__buf_6
Xfanout393 _06263_ vssd1 vssd1 vccd1 vccd1 net393 sky130_fd_sc_hd__buf_4
X_13952_ clknet_leaf_11_clk _01183_ net1098 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[940\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12903_ clknet_leaf_61_clk _00141_ net1136 vssd1 vssd1 vccd1 vccd1 net134 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_1445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13883_ clknet_leaf_64_clk _01114_ net1074 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[871\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11904__S net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12834_ clknet_leaf_19_clk _00072_ net1157 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.ready_data\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_33_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12417__A2 net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_1_Left_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10428__B2 net245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12765_ final_design.VGA_adr\[7\] net796 vssd1 vssd1 vccd1 vccd1 _06401_ sky130_fd_sc_hd__and2_1
XANTENNA__11205__A net245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11716_ net431 net570 _06216_ net295 net1732 vssd1 vssd1 vccd1 vccd1 _00489_ sky130_fd_sc_hd__a32o_1
XFILLER_0_56_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12696_ final_design.VGA_data_control.v_count\[8\] _01398_ vssd1 vssd1 vccd1 vccd1
+ _06337_ sky130_fd_sc_hd__nand2_1
XFILLER_0_72_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11647_ net589 net196 net632 vssd1 vssd1 vccd1 vccd1 _06181_ sky130_fd_sc_hd__and3_1
Xinput13 DAT_I[1] vssd1 vssd1 vccd1 vccd1 net13 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_68_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput24 DAT_I[2] vssd1 vssd1 vccd1 vccd1 net24 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_3_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09169__X _04088_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput35 gpio_in[5] vssd1 vssd1 vccd1 vccd1 net35 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09141__S1 net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput46 mem_adr_start[19] vssd1 vssd1 vccd1 vccd1 net46 sky130_fd_sc_hd__buf_1
X_11578_ net197 net636 vssd1 vssd1 vccd1 vccd1 _06145_ sky130_fd_sc_hd__and2_1
Xinput57 mem_adr_start[29] vssd1 vssd1 vccd1 vccd1 net57 sky130_fd_sc_hd__buf_1
Xinput68 memory_size[0] vssd1 vssd1 vccd1 vccd1 net68 sky130_fd_sc_hd__buf_2
X_13317_ clknet_leaf_49_clk _00548_ net1184 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[305\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold808 final_design.cpu.reg_window\[1001\] vssd1 vssd1 vccd1 vccd1 net2150 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06804__B1 _01504_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput79 memory_size[1] vssd1 vssd1 vccd1 vccd1 net79 sky130_fd_sc_hd__buf_1
X_10529_ net1057 _03784_ vssd1 vssd1 vccd1 vccd1 _05277_ sky130_fd_sc_hd__nand2_1
Xhold819 final_design.cpu.reg_window\[676\] vssd1 vssd1 vccd1 vccd1 net2161 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13248_ clknet_leaf_11_clk _00479_ net1087 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[236\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_72_2660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11875__A net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_2671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10364__B1 net1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13179_ clknet_leaf_66_clk _00410_ net1063 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[167\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11594__B net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11086__S net1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07780__B2 net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07740_ _02687_ _02688_ _02689_ _02690_ net686 net704 vssd1 vssd1 vccd1 vccd1 _02691_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_79_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11313__C1 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13546__CLK clknet_leaf_60_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07671_ net720 _02621_ vssd1 vssd1 vccd1 vccd1 _02622_ sky130_fd_sc_hd__or2_1
XANTENNA__06966__S0 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09410_ _04289_ _04290_ _04327_ _04328_ vssd1 vssd1 vccd1 vccd1 _04329_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_66_2453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11814__S net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_2464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1917 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06622_ final_design.cpu.reg_window\[283\] final_design.cpu.reg_window\[315\] net950
+ vssd1 vssd1 vccd1 vccd1 _01573_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_66_2475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12408__A2 net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_2317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_2328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11616__B1 net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09341_ _04258_ _04259_ vssd1 vssd1 vccd1 vccd1 _04260_ sky130_fd_sc_hd__nor2_1
XFILLER_0_48_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06553_ _01485_ _01489_ net731 _01495_ _01502_ vssd1 vssd1 vccd1 vccd1 _01504_ sky130_fd_sc_hd__a41o_4
XTAP_TAPCELL_ROW_62_2339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09285__A1 net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13696__CLK clknet_leaf_11_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09272_ net82 _04190_ vssd1 vssd1 vccd1 vccd1 _04191_ sky130_fd_sc_hd__or2_2
X_06484_ _01431_ _01432_ _01433_ _01434_ net774 net792 vssd1 vssd1 vccd1 vccd1 _01435_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__09380__S1 net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07391__S0 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08223_ final_design.cpu.reg_window\[75\] final_design.cpu.reg_window\[107\] net835
+ vssd1 vssd1 vccd1 vccd1 _03174_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11402__X _06086_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_12_clk_A clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08245__C1 net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08154_ _01967_ net599 vssd1 vssd1 vccd1 vccd1 _03105_ sky130_fd_sc_hd__nand2_1
XFILLER_0_15_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07105_ _02052_ _02053_ _02054_ _02055_ net765 net780 vssd1 vssd1 vccd1 vccd1 _02056_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__12592__B2 final_design.data_from_mem\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08085_ _01785_ _02799_ vssd1 vssd1 vccd1 vccd1 _03036_ sky130_fd_sc_hd__and2_1
XFILLER_0_28_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07036_ _01983_ _01984_ _01985_ _01986_ net768 net787 vssd1 vssd1 vccd1 vccd1 _01987_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout596_A net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_27_clk_A clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12344__B2 _05959_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13076__CLK clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12380__S net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1847 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08012__A2 _02961_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10355__B1 net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07220__B1 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09255__A _02545_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08987_ _03747_ _03922_ vssd1 vssd1 vccd1 vccd1 _03923_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout763_A _01426_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout384_X net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07938_ final_design.cpu.reg_window\[662\] final_design.cpu.reg_window\[694\] net839
+ vssd1 vssd1 vccd1 vccd1 _02889_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_3_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11855__B1 net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout930_A net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout551_X net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07869_ final_design.cpu.reg_window\[980\] final_design.cpu.reg_window\[1012\] net869
+ vssd1 vssd1 vccd1 vccd1 _02820_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14092__RESET_B net1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout649_X net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12913__CLK clknet_leaf_28_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09608_ _04254_ _04514_ _04526_ vssd1 vssd1 vccd1 vccd1 _04527_ sky130_fd_sc_hd__o21a_1
X_10880_ _05609_ _05610_ _05589_ vssd1 vssd1 vccd1 vccd1 _05611_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_39_804 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11870__A3 net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09539_ net552 _01717_ net551 _01784_ net453 net462 vssd1 vssd1 vccd1 vccd1 _04458_
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_32_1927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12550_ _06213_ net346 net323 net2297 vssd1 vssd1 vccd1 vccd1 _01254_ sky130_fd_sc_hd__a22o_1
XANTENNA__12280__B1 net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11501_ net523 vssd1 vssd1 vccd1 vccd1 _06120_ sky130_fd_sc_hd__inv_2
X_12481_ _06141_ net350 net331 net2037 vssd1 vssd1 vccd1 vccd1 _01187_ sky130_fd_sc_hd__a22o_1
XFILLER_0_34_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11312__X _06007_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14220_ net1278 vssd1 vssd1 vccd1 vccd1 gpio_oeb[32] sky130_fd_sc_hd__buf_2
XFILLER_0_34_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1861 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11432_ net1833 net194 net311 vssd1 vssd1 vccd1 vccd1 _00329_ sky130_fd_sc_hd__mux2_1
XANTENNA__11679__B net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12127__Y _06266_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12583__B2 final_design.data_from_mem\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14151_ clknet_leaf_14_clk _01325_ net1106 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.data_to_VGA\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13419__CLK clknet_leaf_38_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11363_ _04528_ _05143_ net589 _06051_ vssd1 vssd1 vccd1 vccd1 _06052_ sky130_fd_sc_hd__o211a_1
XFILLER_0_46_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13102_ clknet_leaf_45_clk _00333_ net1215 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[90\]
+ sky130_fd_sc_hd__dfrtp_1
X_10314_ _05165_ net1012 vssd1 vssd1 vccd1 vccd1 _05167_ sky130_fd_sc_hd__nor2_2
X_14082_ clknet_leaf_24_clk _01279_ net1161 vssd1 vssd1 vccd1 vccd1 final_design.reqhand.instruction\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_11294_ net660 _03906_ net733 vssd1 vssd1 vccd1 vccd1 _05991_ sky130_fd_sc_hd__o21ai_1
X_13033_ clknet_leaf_40_clk _00264_ net1229 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11695__A net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10245_ net1776 _05114_ _05116_ vssd1 vssd1 vccd1 vccd1 _00013_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_28_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1100 net1105 vssd1 vssd1 vccd1 vccd1 net1100 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09165__A net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1111 net1112 vssd1 vssd1 vccd1 vccd1 net1111 sky130_fd_sc_hd__clkbuf_4
Xfanout1122 net1127 vssd1 vssd1 vccd1 vccd1 net1122 sky130_fd_sc_hd__clkbuf_2
XANTENNA__13569__CLK clknet_leaf_47_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09751__A2 _04222_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10176_ net1052 _05065_ vssd1 vssd1 vccd1 vccd1 _05066_ sky130_fd_sc_hd__and2_2
XANTENNA__12956__RESET_B net1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1133 net1135 vssd1 vssd1 vccd1 vccd1 net1133 sky130_fd_sc_hd__clkbuf_2
Xfanout1144 net1145 vssd1 vssd1 vccd1 vccd1 net1144 sky130_fd_sc_hd__clkbuf_4
Xfanout1155 net1162 vssd1 vssd1 vccd1 vccd1 net1155 sky130_fd_sc_hd__clkbuf_2
Xfanout1166 net1167 vssd1 vssd1 vccd1 vccd1 net1166 sky130_fd_sc_hd__buf_2
XFILLER_0_76_1821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1177 net1178 vssd1 vssd1 vccd1 vccd1 net1177 sky130_fd_sc_hd__clkbuf_4
Xfanout190 _06038_ vssd1 vssd1 vccd1 vccd1 net190 sky130_fd_sc_hd__buf_2
Xfanout1188 net1191 vssd1 vssd1 vccd1 vccd1 net1188 sky130_fd_sc_hd__clkbuf_2
Xfanout1199 net1201 vssd1 vssd1 vccd1 vccd1 net1199 sky130_fd_sc_hd__clkbuf_2
XANTENNA__11846__B1 net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13935_ clknet_leaf_42_clk _01166_ net1226 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[923\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_72_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkload5_A clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09612__B _04530_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13866_ clknet_leaf_59_clk _01097_ net1142 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[854\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11861__A3 net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12817_ net1368 vssd1 vssd1 vccd1 vccd1 _00258_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_80_2940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13797_ clknet_leaf_52_clk _01028_ net1175 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[785\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_80_2951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12748_ net954 _05058_ _06359_ _06372_ _06386_ vssd1 vssd1 vccd1 vccd1 _06387_ sky130_fd_sc_hd__a41o_1
XANTENNA__12271__B1 net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10821__A1 net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10821__B2 _04042_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09019__A1 net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12679_ final_design.VGA_data_control.ready_data\[27\] net1020 net975 final_design.data_from_mem\[27\]
+ vssd1 vssd1 vccd1 vccd1 _06327_ sky130_fd_sc_hd__a22o_1
XFILLER_0_71_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_13_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_13_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1901 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11222__X _05928_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12023__B1 net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13099__CLK clknet_leaf_38_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_2880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_74_2722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold605 final_design.cpu.reg_window\[696\] vssd1 vssd1 vccd1 vccd1 net1947 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10585__B1 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold616 final_design.cpu.reg_window\[939\] vssd1 vssd1 vccd1 vccd1 net1958 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_74_2744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold627 final_design.cpu.reg_window\[175\] vssd1 vssd1 vccd1 vccd1 net1969 sky130_fd_sc_hd__dlygate4sd3_1
Xhold638 final_design.cpu.reg_window\[230\] vssd1 vssd1 vccd1 vccd1 net1980 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold649 final_design.cpu.reg_window\[993\] vssd1 vssd1 vccd1 vccd1 net1991 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_70_2608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_99 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08910_ net257 _03853_ net1014 vssd1 vssd1 vccd1 vccd1 _03855_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10713__S net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09890_ _03638_ _04146_ vssd1 vssd1 vccd1 vccd1 _04809_ sky130_fd_sc_hd__or2_1
XANTENNA__06699__A net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07294__S net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08841_ final_design.CPU_instr_adr\[16\] final_design.CPU_instr_adr\[15\] _03791_
+ vssd1 vssd1 vccd1 vccd1 _03792_ sky130_fd_sc_hd__and3_1
XANTENNA__12936__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_2515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08772_ _03702_ _03722_ vssd1 vssd1 vccd1 vccd1 _03723_ sky130_fd_sc_hd__nand2_1
XFILLER_0_58_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_68_2526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_2537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07723_ _01630_ net605 vssd1 vssd1 vccd1 vccd1 _02674_ sky130_fd_sc_hd__nand2_1
XANTENNA__09803__A net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11301__A2 net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07654_ net616 _02602_ _02603_ _01566_ vssd1 vssd1 vccd1 vccd1 _02605_ sky130_fd_sc_hd__a211oi_1
XANTENNA__07600__S1 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12937__Q net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06605_ final_design.cpu.reg_window\[988\] final_design.cpu.reg_window\[1020\] net946
+ vssd1 vssd1 vccd1 vccd1 _01556_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07585_ final_design.cpu.reg_window\[991\] final_design.cpu.reg_window\[1023\] net859
+ vssd1 vssd1 vccd1 vccd1 _02536_ sky130_fd_sc_hd__mux2_1
XANTENNA__10020__Y _04939_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout344_A net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1086_A net1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09324_ _04234_ _04242_ net491 vssd1 vssd1 vccd1 vccd1 _04243_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12262__B1 net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06536_ _01456_ _01465_ _01474_ vssd1 vssd1 vccd1 vccd1 _01487_ sky130_fd_sc_hd__or3_4
XFILLER_0_76_987 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09255_ _02545_ _02637_ _04173_ vssd1 vssd1 vccd1 vccd1 _04174_ sky130_fd_sc_hd__or3b_1
XANTENNA__12375__S net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout511_A net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06467_ final_design.data_from_mem\[17\] net969 _01417_ vssd1 vssd1 vccd1 vccd1 _01418_
+ sky130_fd_sc_hd__o21a_4
XFILLER_0_1_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout609_A net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08206_ final_design.cpu.reg_window\[526\] final_design.cpu.reg_window\[558\] net813
+ vssd1 vssd1 vccd1 vccd1 _03157_ sky130_fd_sc_hd__mux2_1
XANTENNA__12014__B1 net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09186_ _01452_ net467 net454 vssd1 vssd1 vccd1 vccd1 _04105_ sky130_fd_sc_hd__or3_1
X_08137_ final_design.cpu.reg_window\[653\] final_design.cpu.reg_window\[685\] net854
+ vssd1 vssd1 vccd1 vccd1 _03088_ sky130_fd_sc_hd__mux2_1
XANTENNA__09430__A1 net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08068_ final_design.cpu.reg_window\[530\] final_design.cpu.reg_window\[562\] net844
+ vssd1 vssd1 vccd1 vccd1 _03019_ sky130_fd_sc_hd__mux2_1
XANTENNA__13711__CLK clknet_leaf_40_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12317__A1 net197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout978_A net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout599_X net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07019_ net542 _01968_ vssd1 vssd1 vccd1 vccd1 _01970_ sky130_fd_sc_hd__or2_1
X_10030_ _02837_ _04352_ vssd1 vssd1 vccd1 vccd1 _04949_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_8_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout766_X net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13861__CLK clknet_leaf_52_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09713__A net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11981_ _06183_ net285 net406 net1898 vssd1 vssd1 vccd1 vccd1 _00714_ sky130_fd_sc_hd__a22o_1
XANTENNA__09497__A1 net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13720_ clknet_leaf_65_clk _00951_ net1076 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[708\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_1415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11307__X _06003_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10932_ net963 _05660_ vssd1 vssd1 vccd1 vccd1 _05661_ sky130_fd_sc_hd__nor2_1
XFILLER_0_79_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13651_ clknet_leaf_38_clk _00882_ net1206 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[639\]
+ sky130_fd_sc_hd__dfrtp_1
X_10863_ _05593_ _05594_ vssd1 vssd1 vccd1 vccd1 _05595_ sky130_fd_sc_hd__and2b_1
X_12602_ net2336 net999 net985 final_design.data_from_mem\[20\] vssd1 vssd1 vccd1
+ vccd1 _01295_ sky130_fd_sc_hd__a22o_1
XFILLER_0_71_1773 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12253__B1 net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13582_ clknet_leaf_45_clk _00813_ net1213 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[570\]
+ sky130_fd_sc_hd__dfrtp_1
X_10794_ net76 net1044 vssd1 vssd1 vccd1 vccd1 _05529_ sky130_fd_sc_hd__nor2_1
XANTENNA__10803__A1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12533_ _06258_ net500 net323 net2088 vssd1 vssd1 vccd1 vccd1 _01237_ sky130_fd_sc_hd__a22o_1
XANTENNA__10803__B2 net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13241__CLK clknet_leaf_56_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12005__B1 net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12464_ net673 _06124_ _06260_ vssd1 vssd1 vccd1 vccd1 _06283_ sky130_fd_sc_hd__or3_4
XFILLER_0_53_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14203_ net1261 vssd1 vssd1 vccd1 vccd1 gpio_oeb[15] sky130_fd_sc_hd__buf_2
X_11415_ net1792 net224 net311 vssd1 vssd1 vccd1 vccd1 _00312_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12395_ net2205 net177 net271 vssd1 vssd1 vccd1 vccd1 _01106_ sky130_fd_sc_hd__mux2_1
X_14134_ clknet_leaf_18_clk final_design.vga.h_next_count\[3\] net1113 vssd1 vssd1
+ vccd1 vccd1 final_design.VGA_data_control.h_count\[3\] sky130_fd_sc_hd__dfrtp_2
XANTENNA__09447__X _04366_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11346_ _04917_ net657 vssd1 vssd1 vccd1 vccd1 _06037_ sky130_fd_sc_hd__nand2_1
XANTENNA__13391__CLK clknet_leaf_42_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07983__A1 net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14065_ clknet_leaf_15_clk _00027_ net1091 vssd1 vssd1 vccd1 vccd1 final_design.uart.BAUD_counter\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10319__B1 net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11277_ _01939_ _05947_ _05974_ _05975_ vssd1 vssd1 vccd1 vccd1 _05976_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__09607__B _04516_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13016_ clknet_leaf_62_clk _00247_ net1119 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_10228_ final_design.uart.BAUD_counter\[10\] _05104_ net798 vssd1 vssd1 vccd1 vccd1
+ _05106_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07735__A1 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10159_ net1048 _05050_ final_design.VGA_data_control.h_count\[5\] vssd1 vssd1 vccd1
+ vccd1 _05055_ sky130_fd_sc_hd__a21oi_1
Xhold2 final_design.cpu.reg_window\[8\] vssd1 vssd1 vccd1 vccd1 net1344 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11819__A0 net221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11872__B net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12087__A3 net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12492__B1 net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13918_ clknet_leaf_13_clk _01149_ net1099 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[906\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10488__B net1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13849_ clknet_leaf_55_clk _01080_ net1178 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[837\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11047__A1 net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12244__B1 net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07370_ final_design.cpu.reg_window\[579\] final_design.cpu.reg_window\[611\] net908
+ vssd1 vssd1 vccd1 vccd1 _02321_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12195__S net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09040_ _03694_ _03729_ _03692_ vssd1 vssd1 vccd1 vccd1 _03970_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_2_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_2806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_2817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13734__CLK clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold402 final_design.cpu.reg_window\[73\] vssd1 vssd1 vccd1 vccd1 net1744 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07649__S1 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold413 final_design.cpu.reg_window\[911\] vssd1 vssd1 vccd1 vccd1 net1755 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_1775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold424 final_design.cpu.reg_window\[588\] vssd1 vssd1 vccd1 vccd1 net1766 sky130_fd_sc_hd__dlygate4sd3_1
Xhold435 final_design.cpu.reg_window\[454\] vssd1 vssd1 vccd1 vccd1 net1777 sky130_fd_sc_hd__dlygate4sd3_1
Xhold446 final_design.cpu.reg_window\[595\] vssd1 vssd1 vccd1 vccd1 net1788 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkload31_A clknet_leaf_55_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold457 final_design.cpu.reg_window\[755\] vssd1 vssd1 vccd1 vccd1 net1799 sky130_fd_sc_hd__dlygate4sd3_1
Xhold468 final_design.cpu.reg_window\[961\] vssd1 vssd1 vccd1 vccd1 net1810 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11539__S net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09942_ _03421_ _04149_ _03390_ vssd1 vssd1 vccd1 vccd1 _04861_ sky130_fd_sc_hd__a21oi_1
Xhold479 final_design.cpu.reg_window\[459\] vssd1 vssd1 vccd1 vccd1 net1821 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09517__B _04435_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout904 net905 vssd1 vssd1 vccd1 vccd1 net904 sky130_fd_sc_hd__clkbuf_4
XANTENNA__13884__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1915 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout915 net917 vssd1 vssd1 vccd1 vccd1 net915 sky130_fd_sc_hd__buf_4
XFILLER_0_0_483 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout926 net927 vssd1 vssd1 vccd1 vccd1 net926 sky130_fd_sc_hd__clkbuf_4
X_09873_ net475 _04109_ _04308_ vssd1 vssd1 vccd1 vccd1 _04792_ sky130_fd_sc_hd__or3_1
Xfanout937 net940 vssd1 vssd1 vccd1 vccd1 net937 sky130_fd_sc_hd__clkbuf_4
Xfanout948 net950 vssd1 vssd1 vccd1 vccd1 net948 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout294_A net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout959 _04041_ vssd1 vssd1 vccd1 vccd1 net959 sky130_fd_sc_hd__clkbuf_4
X_08824_ _03660_ _03773_ _03661_ _03659_ vssd1 vssd1 vccd1 vccd1 _03775_ sky130_fd_sc_hd__o211a_1
Xhold1102 final_design.cpu.reg_window\[120\] vssd1 vssd1 vccd1 vccd1 net2444 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1113 final_design.cpu.reg_window\[305\] vssd1 vssd1 vccd1 vccd1 net2455 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1001_A _05239_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1124 final_design.cpu.reg_window\[616\] vssd1 vssd1 vccd1 vccd1 net2466 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1135 final_design.cpu.reg_window\[261\] vssd1 vssd1 vccd1 vccd1 net2477 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1146 final_design.cpu.reg_window\[173\] vssd1 vssd1 vccd1 vccd1 net2488 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13114__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09533__A net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1157 final_design.cpu.reg_window\[369\] vssd1 vssd1 vccd1 vccd1 net2499 sky130_fd_sc_hd__dlygate4sd3_1
X_08755_ _01366_ _02297_ vssd1 vssd1 vccd1 vccd1 _03706_ sky130_fd_sc_hd__nor2_1
Xhold1168 final_design.cpu.reg_window\[289\] vssd1 vssd1 vccd1 vccd1 net2510 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout461_A _03519_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12078__A3 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1179 final_design.cpu.reg_window\[309\] vssd1 vssd1 vccd1 vccd1 net2521 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout559_A net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11286__A1 final_design.data_from_mem\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07706_ final_design.cpu.reg_window\[539\] final_design.cpu.reg_window\[571\] net861
+ vssd1 vssd1 vccd1 vccd1 _02657_ sky130_fd_sc_hd__mux2_1
XANTENNA__12483__B1 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08686_ _02325_ net483 vssd1 vssd1 vccd1 vccd1 _03637_ sky130_fd_sc_hd__nor2_1
XFILLER_0_7_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10398__B _05181_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07637_ _02584_ _02585_ _02586_ _02587_ net687 net705 vssd1 vssd1 vccd1 vccd1 _02588_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_0_176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout726_A _01493_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13264__CLK clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout347_X net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12235__B1 net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06892__A net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1588 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07568_ final_design.cpu.reg_window\[415\] final_design.cpu.reg_window\[447\] net859
+ vssd1 vssd1 vccd1 vccd1 _02519_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11589__A2 net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09307_ net492 _04225_ _04205_ vssd1 vssd1 vccd1 vccd1 _04226_ sky130_fd_sc_hd__or3b_1
X_06519_ final_design.reqhand.instruction\[0\] final_design.reqhand.instruction\[1\]
+ vssd1 vssd1 vccd1 vccd1 _01470_ sky130_fd_sc_hd__nand2_1
XFILLER_0_36_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout514_X net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09651__A1 net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07499_ _02032_ _02449_ vssd1 vssd1 vccd1 vccd1 _02450_ sky130_fd_sc_hd__or2_1
XANTENNA__12250__A3 net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09238_ _04144_ _04153_ _04154_ _04156_ vssd1 vssd1 vccd1 vccd1 _04157_ sky130_fd_sc_hd__a31oi_4
XTAP_TAPCELL_ROW_40_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09169_ _03631_ net659 vssd1 vssd1 vccd1 vccd1 _04088_ sky130_fd_sc_hd__or2_4
XFILLER_0_31_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11200_ _03995_ _05907_ net732 vssd1 vssd1 vccd1 vccd1 _05908_ sky130_fd_sc_hd__mux2_1
X_12180_ _06121_ net501 _06270_ net1807 vssd1 vssd1 vccd1 vccd1 _00899_ sky130_fd_sc_hd__a22o_1
XANTENNA__09954__A2 net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11957__B net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout883_X net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11449__S net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11131_ _05841_ net588 vssd1 vssd1 vccd1 vccd1 _05846_ sky130_fd_sc_hd__nand2_2
XFILLER_0_8_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold980 final_design.cpu.reg_window\[297\] vssd1 vssd1 vccd1 vccd1 net2322 sky130_fd_sc_hd__dlygate4sd3_1
Xhold991 final_design.cpu.reg_window\[32\] vssd1 vssd1 vccd1 vccd1 net2333 sky130_fd_sc_hd__dlygate4sd3_1
X_11062_ _05783_ _05784_ vssd1 vssd1 vccd1 vccd1 _05785_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_38_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07717__A1 net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10013_ net470 _04834_ _04931_ net483 vssd1 vssd1 vccd1 vccd1 _04932_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_34_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07662__S net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input22_A DAT_I[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09443__A net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12069__A3 net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11184__S net247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13607__CLK clknet_leaf_62_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12474__B1 net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11964_ _06166_ net280 net404 net1777 vssd1 vssd1 vccd1 vccd1 _00697_ sky130_fd_sc_hd__a22o_1
XFILLER_0_59_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13703_ clknet_leaf_63_clk _00934_ net1120 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[691\]
+ sky130_fd_sc_hd__dfrtp_1
X_10915_ _05643_ _05644_ vssd1 vssd1 vccd1 vccd1 _05645_ sky130_fd_sc_hd__or2_1
X_11895_ net217 net2253 net272 vssd1 vssd1 vccd1 vccd1 _00637_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_15_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11912__S net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13634_ clknet_leaf_3_clk _00865_ net1067 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[622\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12226__B1 net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10846_ net46 _05566_ _05575_ _05577_ vssd1 vssd1 vccd1 vccd1 _05579_ sky130_fd_sc_hd__and4_1
XFILLER_0_71_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13757__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13565_ clknet_leaf_2_clk _00796_ net1065 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[553\]
+ sky130_fd_sc_hd__dfrtp_1
X_10777_ net75 _05486_ _05512_ vssd1 vssd1 vccd1 vccd1 _05513_ sky130_fd_sc_hd__a21bo_1
XANTENNA__10528__S net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12241__A3 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12516_ _06178_ net351 net329 net1702 vssd1 vssd1 vccd1 vccd1 _01221_ sky130_fd_sc_hd__a22o_1
X_13496_ clknet_leaf_65_clk _00727_ net1119 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[484\]
+ sky130_fd_sc_hd__dfrtp_1
X_12447_ net1755 net206 net334 vssd1 vssd1 vccd1 vccd1 _01154_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12378_ net1714 net207 net268 vssd1 vssd1 vccd1 vccd1 _01089_ sky130_fd_sc_hd__mux2_1
XANTENNA__08602__C1 _02419_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14117_ clknet_leaf_13_clk _01314_ net1089 vssd1 vssd1 vccd1 vccd1 final_design.reqhand.data_from_UART\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_11329_ _01756_ net641 _06021_ net643 _06020_ vssd1 vssd1 vccd1 vccd1 _06022_ sky130_fd_sc_hd__a221o_1
XFILLER_0_5_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12900__RESET_B net1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13137__CLK clknet_leaf_34_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14048_ clknet_leaf_16_clk _00009_ net1092 vssd1 vssd1 vccd1 vccd1 final_design.uart.BAUD_counter\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_66_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11883__A net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06870_ _01485_ _01489_ _01495_ _01820_ _01502_ vssd1 vssd1 vccd1 vccd1 _01821_ sky130_fd_sc_hd__a41o_4
XFILLER_0_78_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13287__CLK clknet_leaf_63_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11268__A1 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08540_ final_design.cpu.reg_window\[449\] final_design.cpu.reg_window\[481\] net833
+ vssd1 vssd1 vccd1 vccd1 _03491_ sky130_fd_sc_hd__mux2_1
XANTENNA__12465__B1 net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08133__A1 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09640__X _04559_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08471_ net596 _03415_ _03417_ _02294_ vssd1 vssd1 vccd1 vccd1 _03422_ sky130_fd_sc_hd__o211a_1
XANTENNA__09881__A1 net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11822__S net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07422_ final_design.cpu.reg_window\[129\] final_design.cpu.reg_window\[161\] net916
+ vssd1 vssd1 vccd1 vccd1 _02373_ sky130_fd_sc_hd__mux2_1
XANTENNA__13077__RESET_B net1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12217__B1 net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12768__A1 final_design.VGA_adr\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10946__B net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13006__RESET_B net1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07353_ final_design.cpu.reg_window\[387\] final_design.cpu.reg_window\[419\] net915
+ vssd1 vssd1 vccd1 vccd1 _02304_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09094__C1 net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12232__A3 net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11123__A net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07284_ final_design.cpu.reg_window\[710\] final_design.cpu.reg_window\[742\] net901
+ vssd1 vssd1 vccd1 vccd1 _02235_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09023_ _03687_ _03733_ vssd1 vssd1 vccd1 vccd1 _03955_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout307_A _06095_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold210 final_design.cpu.reg_window\[966\] vssd1 vssd1 vccd1 vccd1 net1552 sky130_fd_sc_hd__dlygate4sd3_1
Xhold221 final_design.cpu.reg_window\[216\] vssd1 vssd1 vccd1 vccd1 net1563 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09936__A2 net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold232 final_design.cpu.reg_window\[845\] vssd1 vssd1 vccd1 vccd1 net1574 sky130_fd_sc_hd__dlygate4sd3_1
Xhold243 net124 vssd1 vssd1 vccd1 vccd1 net1585 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold254 final_design.cpu.reg_window\[569\] vssd1 vssd1 vccd1 vccd1 net1596 sky130_fd_sc_hd__dlygate4sd3_1
Xhold265 net148 vssd1 vssd1 vccd1 vccd1 net1607 sky130_fd_sc_hd__dlygate4sd3_1
Xhold276 final_design.cpu.reg_window\[678\] vssd1 vssd1 vccd1 vccd1 net1618 sky130_fd_sc_hd__dlygate4sd3_1
Xhold287 final_design.cpu.reg_window\[244\] vssd1 vssd1 vccd1 vccd1 net1629 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout701 _01752_ vssd1 vssd1 vccd1 vccd1 net701 sky130_fd_sc_hd__clkbuf_4
Xhold298 final_design.cpu.reg_window\[583\] vssd1 vssd1 vccd1 vccd1 net1640 sky130_fd_sc_hd__dlygate4sd3_1
X_09925_ _03424_ _03561_ vssd1 vssd1 vccd1 vccd1 _04844_ sky130_fd_sc_hd__nor2_1
Xfanout712 net713 vssd1 vssd1 vccd1 vccd1 net712 sky130_fd_sc_hd__buf_2
XANTENNA__14062__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout723 net724 vssd1 vssd1 vccd1 vccd1 net723 sky130_fd_sc_hd__clkbuf_8
Xfanout734 net736 vssd1 vssd1 vccd1 vccd1 net734 sky130_fd_sc_hd__buf_2
Xfanout745 net746 vssd1 vssd1 vccd1 vccd1 net745 sky130_fd_sc_hd__buf_4
XANTENNA_fanout297_X net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout676_A net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout756 _01427_ vssd1 vssd1 vccd1 vccd1 net756 sky130_fd_sc_hd__buf_4
Xfanout767 net768 vssd1 vssd1 vccd1 vccd1 net767 sky130_fd_sc_hd__buf_4
X_09856_ _04773_ _04774_ _04220_ vssd1 vssd1 vccd1 vccd1 _04775_ sky130_fd_sc_hd__a21o_1
Xfanout778 net779 vssd1 vssd1 vccd1 vccd1 net778 sky130_fd_sc_hd__clkbuf_4
Xfanout789 net790 vssd1 vssd1 vccd1 vccd1 net789 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_52_1990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08807_ final_design.CPU_instr_adr\[22\] _01755_ vssd1 vssd1 vccd1 vccd1 _03758_
+ sky130_fd_sc_hd__xnor2_1
X_09787_ _03388_ _03421_ _04149_ _03389_ _03358_ vssd1 vssd1 vccd1 vccd1 _04706_ sky130_fd_sc_hd__a311o_1
X_06999_ final_design.cpu.reg_window\[207\] final_design.cpu.reg_window\[239\] net889
+ vssd1 vssd1 vccd1 vccd1 _01950_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout843_A net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout464_X net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11259__A1 final_design.data_from_mem\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08738_ final_design.CPU_instr_adr\[11\] _02097_ vssd1 vssd1 vccd1 vccd1 _03689_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_16_1527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout631_X net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08669_ _01999_ _02029_ _02061_ vssd1 vssd1 vccd1 vccd1 _03620_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout729_X net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10700_ _05400_ _05418_ _05419_ vssd1 vssd1 vccd1 vccd1 _05440_ sky130_fd_sc_hd__a21o_1
XANTENNA__12208__B1 net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11680_ net427 net564 _06198_ net294 net1709 vssd1 vssd1 vccd1 vccd1 _00471_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_46_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10631_ _05349_ _05368_ _05369_ vssd1 vssd1 vccd1 vccd1 _05374_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_46_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12223__A3 net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1295 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13350_ clknet_leaf_51_clk _00581_ net1171 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[338\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11431__A1 _06017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10562_ _05306_ _05308_ net1402 net1029 vssd1 vssd1 vccd1 vccd1 _00178_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_49_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12301_ net1979 net240 net364 vssd1 vssd1 vccd1 vccd1 _01015_ sky130_fd_sc_hd__mux2_1
XANTENNA__11982__A2 net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14117__Q final_design.reqhand.data_from_UART\[7\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_13281_ clknet_leaf_48_clk _00512_ net1185 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[269\]
+ sky130_fd_sc_hd__dfrtp_1
X_10493_ net964 _05240_ vssd1 vssd1 vccd1 vccd1 _05243_ sky130_fd_sc_hd__or2_1
XFILLER_0_66_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11320__X _06014_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12232_ net566 _06162_ net506 net373 net1537 vssd1 vssd1 vccd1 vccd1 _00949_ sky130_fd_sc_hd__a32o_1
XANTENNA__11687__B net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06561__S net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08286__S1 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09483__S0 net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11195__B1 net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11734__A2 net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14209__1267 vssd1 vssd1 vccd1 vccd1 _14209__1267/HI net1267 sky130_fd_sc_hd__conb_1
X_12163_ _06117_ _06260_ vssd1 vssd1 vccd1 vccd1 _06270_ sky130_fd_sc_hd__or2_4
XTAP_TAPCELL_ROW_36_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11114_ _05065_ _05082_ _05832_ vssd1 vssd1 vccd1 vccd1 _05833_ sky130_fd_sc_hd__and3b_1
X_12094_ net673 _06091_ net507 vssd1 vssd1 vccd1 vccd1 _06265_ sky130_fd_sc_hd__and3_2
XANTENNA__08038__S1 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11907__S net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11045_ final_design.CPU_instr_adr\[28\] _03829_ net1059 vssd1 vssd1 vccd1 vccd1
+ _05769_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1889 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09173__A _03635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input25_X net25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11990__X _06257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1610 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09538__S1 net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12996_ net1327 _00227_ net1195 vssd1 vssd1 vccd1 vccd1 final_design.CPU_instr_adr\[16\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__07549__S0 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1020 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09901__A _04124_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11947_ _06148_ net285 net410 net2116 vssd1 vssd1 vccd1 vccd1 _00682_ sky130_fd_sc_hd__a22o_1
XANTENNA__06677__A1 final_design.data_from_mem\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11878_ _06112_ net291 net519 net2045 vssd1 vssd1 vccd1 vccd1 _00622_ sky130_fd_sc_hd__a22o_1
XFILLER_0_39_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08517__A net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13617_ clknet_leaf_34_clk _00848_ net1237 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[605\]
+ sky130_fd_sc_hd__dfrtp_1
X_10829_ _01385_ _05539_ _05544_ vssd1 vssd1 vccd1 vccd1 _05563_ sky130_fd_sc_hd__o21ba_1
XANTENNA__09615__A1 _03418_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1761 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11422__A1 net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13548_ clknet_leaf_45_clk _00779_ net1204 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[536\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09091__A2 net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11973__A2 net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13479_ clknet_leaf_63_clk _00710_ net1123 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[467\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_971 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14085__CLK clknet_leaf_25_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1892 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07971_ _02918_ _02919_ _02920_ _02921_ net682 net693 vssd1 vssd1 vccd1 vccd1 _02922_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__11817__S net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09710_ _03068_ _03101_ _04627_ net447 vssd1 vssd1 vccd1 vccd1 _04629_ sky130_fd_sc_hd__a31o_1
X_06922_ _01869_ _01870_ _01871_ _01872_ net773 net791 vssd1 vssd1 vccd1 vccd1 _01873_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__12061__X _06264_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08398__S net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_6_clk_X clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09641_ net478 _04258_ _04259_ net492 vssd1 vssd1 vccd1 vccd1 _04560_ sky130_fd_sc_hd__o31a_2
X_06853_ final_design.cpu.reg_window\[788\] final_design.cpu.reg_window\[820\] net948
+ vssd1 vssd1 vccd1 vccd1 _01804_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06500__A net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13922__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09572_ net473 _04260_ _04490_ vssd1 vssd1 vccd1 vccd1 _04491_ sky130_fd_sc_hd__o21a_1
XANTENNA__10022__A net68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06784_ final_design.cpu.reg_window\[150\] final_design.cpu.reg_window\[182\] net918
+ vssd1 vssd1 vccd1 vccd1 _01735_ sky130_fd_sc_hd__mux2_1
X_08523_ _03470_ _03471_ _03472_ _03473_ net679 net699 vssd1 vssd1 vccd1 vccd1 _03474_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_52_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08201__S1 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08657__A2 _02635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout257_A net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08454_ final_design.cpu.reg_window\[772\] final_design.cpu.reg_window\[804\] net824
+ vssd1 vssd1 vccd1 vccd1 _03405_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07405_ _02343_ _02344_ _02355_ net883 vssd1 vssd1 vccd1 vccd1 _02356_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_50_1451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08385_ final_design.cpu.reg_window\[198\] final_design.cpu.reg_window\[230\] net820
+ vssd1 vssd1 vccd1 vccd1 _03336_ sky130_fd_sc_hd__mux2_1
XANTENNA__09606__A1 _04222_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout424_A _05877_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12205__A3 net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1166_A net1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08146__B _03096_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07336_ _02283_ _02284_ _02285_ _02286_ net767 net787 vssd1 vssd1 vccd1 vccd1 _02287_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_11_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13302__CLK clknet_leaf_59_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11964__A2 net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11788__A net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12383__S net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07267_ final_design.cpu.reg_window\[454\] final_design.cpu.reg_window\[486\] net904
+ vssd1 vssd1 vccd1 vccd1 _02218_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout212_X net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09006_ _03791_ _03939_ vssd1 vssd1 vccd1 vccd1 _03940_ sky130_fd_sc_hd__or2_1
XFILLER_0_42_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09258__A net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07198_ final_design.cpu.reg_window\[585\] final_design.cpu.reg_window\[617\] net888
+ vssd1 vssd1 vccd1 vccd1 _02149_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout793_A net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13452__CLK clknet_leaf_45_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout960_A _04040_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout520 _06239_ vssd1 vssd1 vccd1 vccd1 net520 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout679_X net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout531 _02266_ vssd1 vssd1 vccd1 vccd1 net531 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_50_1905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout542 net543 vssd1 vssd1 vccd1 vccd1 net542 sky130_fd_sc_hd__buf_2
X_09908_ _04808_ _04826_ vssd1 vssd1 vccd1 vccd1 _04827_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_50_1916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout553 _06238_ vssd1 vssd1 vccd1 vccd1 net553 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_50_1927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout564 net565 vssd1 vssd1 vccd1 vccd1 net564 sky130_fd_sc_hd__clkbuf_4
Xfanout575 net576 vssd1 vssd1 vccd1 vccd1 net575 sky130_fd_sc_hd__clkbuf_2
Xfanout586 net587 vssd1 vssd1 vccd1 vccd1 net586 sky130_fd_sc_hd__clkbuf_4
X_09839_ _04754_ _04757_ vssd1 vssd1 vccd1 vccd1 _04758_ sky130_fd_sc_hd__nand2_1
Xfanout597 net601 vssd1 vssd1 vccd1 vccd1 net597 sky130_fd_sc_hd__buf_2
X_12850_ clknet_leaf_19_clk _00088_ net1112 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.ready_data\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07940__S net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11801_ net2533 net414 net285 _06032_ vssd1 vssd1 vccd1 vccd1 _00554_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_29_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_1856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11315__X _06010_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10455__A2 net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11732_ net587 net423 _06224_ net296 net1638 vssd1 vssd1 vccd1 vccd1 _00497_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_44_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11652__A1 net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11663_ net180 net632 vssd1 vssd1 vccd1 vccd1 _06189_ sky130_fd_sc_hd__and2_1
XFILLER_0_0_1901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13402_ clknet_leaf_6_clk _00633_ net1129 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[390\]
+ sky130_fd_sc_hd__dfrtp_1
X_10614_ _05357_ net955 net960 _05356_ vssd1 vssd1 vccd1 vccd1 _05358_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_36_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11594_ net182 net636 vssd1 vssd1 vccd1 vccd1 _06153_ sky130_fd_sc_hd__and2_1
XFILLER_0_68_1745 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07703__S0 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11955__A2 net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13333_ clknet_leaf_56_clk _00564_ net1145 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[321\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_36_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10545_ _05290_ _05291_ vssd1 vssd1 vccd1 vccd1 _05292_ sky130_fd_sc_hd__nor2_1
XFILLER_0_52_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_1789 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13264_ clknet_leaf_33_clk _00495_ net1232 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[252\]
+ sky130_fd_sc_hd__dfrtp_1
X_10476_ net961 _05226_ vssd1 vssd1 vccd1 vccd1 _05227_ sky130_fd_sc_hd__or2_1
X_12215_ net572 _06143_ net508 net379 net2103 vssd1 vssd1 vccd1 vccd1 _00933_ sky130_fd_sc_hd__a32o_1
XFILLER_0_20_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13195_ clknet_leaf_38_clk _00426_ net1191 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[183\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_62_1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12146_ net222 net2301 net387 vssd1 vssd1 vccd1 vccd1 _00867_ sky130_fd_sc_hd__mux2_1
XANTENNA__13945__CLK clknet_leaf_54_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12077_ net558 _05973_ net502 net392 net1750 vssd1 vssd1 vccd1 vccd1 _00802_ sky130_fd_sc_hd__a32o_1
XFILLER_0_79_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08336__B2 net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11028_ _05731_ _05749_ vssd1 vssd1 vccd1 vccd1 _05752_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_75_1705 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11209__Y _05916_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1885 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08431__S1 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_1749 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06898__A1 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09631__A net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12979_ clknet_leaf_25_clk _00004_ net1156 vssd1 vssd1 vccd1 vccd1 wb_manage.curr_state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11225__X _05930_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08195__S0 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13325__CLK clknet_leaf_44_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_2381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_2392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_2245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_2256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_16 _06228_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_2267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_27 _06257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08170_ final_design.cpu.reg_window\[911\] final_design.cpu.reg_window\[943\] net811
+ vssd1 vssd1 vccd1 vccd1 _03121_ sky130_fd_sc_hd__mux2_1
XANTENNA__08534__X _03485_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06990__A _01937_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11946__A2 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07121_ _02068_ _02069_ _02070_ _02071_ net769 net790 vssd1 vssd1 vccd1 vccd1 _02072_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_67_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13475__CLK clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07052_ final_design.cpu.reg_window\[333\] final_design.cpu.reg_window\[365\] net934
+ vssd1 vssd1 vccd1 vccd1 _02003_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_11_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput101 net101 vssd1 vssd1 vccd1 vccd1 ADR_O[0] sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_58_2174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput112 net112 vssd1 vssd1 vccd1 vccd1 ADR_O[1] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_2_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_58_2185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput123 net123 vssd1 vssd1 vccd1 vccd1 ADR_O[2] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_58_2196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput134 net134 vssd1 vssd1 vccd1 vccd1 DAT_O[0] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_54_2038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput145 net145 vssd1 vssd1 vccd1 vccd1 DAT_O[1] sky130_fd_sc_hd__buf_2
XANTENNA__10017__A net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_2049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput156 net156 vssd1 vssd1 vccd1 vccd1 DAT_O[2] sky130_fd_sc_hd__buf_2
XFILLER_0_80_1466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput167 net167 vssd1 vssd1 vccd1 vccd1 SEL_O[1] sky130_fd_sc_hd__buf_2
XANTENNA__10382__B2 final_design.data_from_mem\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07783__C1 _01686_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13439__RESET_B net1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07954_ _01909_ net603 vssd1 vssd1 vccd1 vccd1 _02905_ sky130_fd_sc_hd__nand2_1
XANTENNA__11774__C net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06905_ net548 _01854_ vssd1 vssd1 vccd1 vccd1 _01856_ sky130_fd_sc_hd__or2_1
XFILLER_0_39_1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07885_ _02833_ _02835_ vssd1 vssd1 vccd1 vccd1 _02836_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout374_A net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09624_ _04072_ _04540_ _04541_ _04542_ vssd1 vssd1 vccd1 vccd1 _04543_ sky130_fd_sc_hd__or4_1
XANTENNA__14100__CLK clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06836_ final_design.data_from_mem\[21\] net971 _01786_ vssd1 vssd1 vccd1 vccd1 _01787_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_39_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07760__S net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06984__S1 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09555_ net448 _04472_ _04470_ net729 vssd1 vssd1 vccd1 vccd1 _04474_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_6_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06767_ net886 _01710_ _01716_ _01703_ _01704_ vssd1 vssd1 vccd1 vccd1 _01718_ sky130_fd_sc_hd__a32o_1
XANTENNA__12378__S net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09288__C1 _01535_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout639_A _06093_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08506_ net608 _03450_ _03451_ _02326_ vssd1 vssd1 vccd1 vccd1 _03457_ sky130_fd_sc_hd__a211o_1
XFILLER_0_78_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11634__A1 net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09486_ _01566_ net453 _04207_ net467 vssd1 vssd1 vccd1 vccd1 _04405_ sky130_fd_sc_hd__a211o_1
X_14208__1266 vssd1 vssd1 vccd1 vccd1 _14208__1266/HI net1266 sky130_fd_sc_hd__conb_1
X_06698_ _01645_ _01646_ _01647_ _01648_ net774 net792 vssd1 vssd1 vccd1 vccd1 _01649_
+ sky130_fd_sc_hd__mux4_1
X_08437_ net530 _03386_ vssd1 vssd1 vccd1 vccd1 _03388_ sky130_fd_sc_hd__nand2b_1
XANTENNA_fanout427_X net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13818__CLK clknet_leaf_63_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08368_ _03315_ _03316_ _03317_ _03318_ net674 net691 vssd1 vssd1 vccd1 vccd1 _03319_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_34_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11398__B1 net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11937__A2 net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1899 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07319_ _02268_ _02269_ vssd1 vssd1 vccd1 vccd1 _02270_ sky130_fd_sc_hd__and2b_1
X_08299_ net716 _03249_ vssd1 vssd1 vccd1 vccd1 _03250_ sky130_fd_sc_hd__nor2_1
XFILLER_0_46_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11311__A net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10330_ net1509 net1010 net987 final_design.data_from_mem\[15\] vssd1 vssd1 vccd1
+ vccd1 _00087_ sky130_fd_sc_hd__a22o_1
XANTENNA__07161__S1 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout796_X net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12842__CLK clknet_leaf_15_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13968__CLK clknet_leaf_34_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10261_ net1568 _05124_ _05126_ vssd1 vssd1 vccd1 vccd1 _00020_ sky130_fd_sc_hd__a21oi_1
XANTENNA__06899__X _01850_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12000_ _06202_ net277 net400 net2318 vssd1 vssd1 vccd1 vccd1 _00731_ sky130_fd_sc_hd__a22o_1
XANTENNA__12362__A2 net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1063 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10192_ final_design.uart.BAUD_counter\[2\] final_design.uart.BAUD_counter\[7\] final_design.uart.BAUD_counter\[6\]
+ final_design.uart.BAUD_counter\[3\] vssd1 vssd1 vccd1 vccd1 _05081_ sky130_fd_sc_hd__or4b_1
XANTENNA__08620__A _02127_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout963_X net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10373__B2 final_design.data_from_mem\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11457__S net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout350 _06277_ vssd1 vssd1 vccd1 vccd1 net350 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09515__A0 net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout361 net363 vssd1 vssd1 vccd1 vccd1 net361 sky130_fd_sc_hd__buf_4
XANTENNA__07236__A _02185_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13109__RESET_B net1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout372 net373 vssd1 vssd1 vccd1 vccd1 net372 sky130_fd_sc_hd__buf_4
Xfanout383 _06269_ vssd1 vssd1 vccd1 vccd1 net383 sky130_fd_sc_hd__clkbuf_8
X_13951_ clknet_leaf_7_clk _01182_ net1130 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[939\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_17_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout394 net395 vssd1 vssd1 vccd1 vccd1 net394 sky130_fd_sc_hd__buf_4
X_12902_ clknet_leaf_25_clk _00140_ net1155 vssd1 vssd1 vccd1 vccd1 net169 sky130_fd_sc_hd__dfrtp_4
X_13882_ clknet_leaf_58_clk _01113_ net1125 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[870\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11873__B2 net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13348__CLK clknet_leaf_52_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12833_ net1351 vssd1 vssd1 vccd1 vccd1 _00274_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_1891 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09818__A1 _04222_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12764_ net954 _06382_ _06399_ vssd1 vssd1 vccd1 vccd1 _06400_ sky130_fd_sc_hd__and3_1
XFILLER_0_55_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11715_ net194 net627 vssd1 vssd1 vccd1 vccd1 _06216_ sky130_fd_sc_hd__and2_1
X_12695_ final_design.VGA_data_control.v_count\[5\] _06335_ vssd1 vssd1 vccd1 vccd1
+ _06336_ sky130_fd_sc_hd__nor2_1
XANTENNA__13498__CLK clknet_leaf_58_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11920__S net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11646_ net435 net585 _06180_ net300 net1506 vssd1 vssd1 vccd1 vccd1 _00455_ sky130_fd_sc_hd__a32o_1
Xinput14 DAT_I[20] vssd1 vssd1 vccd1 vccd1 net14 sky130_fd_sc_hd__buf_1
XANTENNA__11928__A2 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput25 DAT_I[30] vssd1 vssd1 vccd1 vccd1 net25 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_25_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput36 mem_adr_start[0] vssd1 vssd1 vccd1 vccd1 net36 sky130_fd_sc_hd__buf_1
X_11577_ net567 net422 _06144_ net303 net2006 vssd1 vssd1 vccd1 vccd1 _00422_ sky130_fd_sc_hd__a32o_1
XFILLER_0_24_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput47 mem_adr_start[1] vssd1 vssd1 vccd1 vccd1 net47 sky130_fd_sc_hd__buf_1
XFILLER_0_68_1575 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13316_ clknet_leaf_52_clk _00547_ net1174 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[304\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput58 mem_adr_start[2] vssd1 vssd1 vccd1 vccd1 net58 sky130_fd_sc_hd__clkbuf_2
XANTENNA__11221__A _04744_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput69 memory_size[10] vssd1 vssd1 vccd1 vccd1 net69 sky130_fd_sc_hd__clkbuf_2
X_10528_ final_design.CPU_instr_adr\[4\] _05275_ net1053 vssd1 vssd1 vccd1 vccd1 _05276_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold809 final_design.cpu.reg_window\[484\] vssd1 vssd1 vccd1 vccd1 net2151 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13247_ clknet_leaf_7_clk _00478_ net1134 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[235\]
+ sky130_fd_sc_hd__dfrtp_1
X_10459_ net1800 net1033 _05213_ net248 vssd1 vssd1 vccd1 vccd1 _00170_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_72_2650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12353__A2 net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11156__A3 net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07845__S net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_2661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_72_2672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13178_ clknet_leaf_6_clk _00409_ net1128 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[166\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11875__B net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10364__B2 final_design.data_from_mem\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11561__B1 net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12129_ _05840_ _05841_ net231 vssd1 vssd1 vccd1 vccd1 _06268_ sky130_fd_sc_hd__and3_2
XANTENNA__14123__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07670_ _02617_ _02618_ _02619_ _02620_ net684 net703 vssd1 vssd1 vccd1 vccd1 _02621_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_75_1546 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11864__B2 net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06985__A net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06966__S1 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06621_ final_design.cpu.reg_window\[347\] final_design.cpu.reg_window\[379\] net950
+ vssd1 vssd1 vccd1 vccd1 _01572_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_66_2454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_2318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09340_ _04078_ _04102_ net467 vssd1 vssd1 vccd1 vccd1 _04259_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_73_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11616__A1 net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06552_ _01484_ _01488_ net734 _01494_ _01501_ vssd1 vssd1 vccd1 vccd1 _01503_ sky130_fd_sc_hd__o41a_4
XTAP_TAPCELL_ROW_62_2329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09271_ net80 net81 _04189_ vssd1 vssd1 vccd1 vccd1 _04190_ sky130_fd_sc_hd__or3_1
X_06483_ final_design.cpu.reg_window\[158\] final_design.cpu.reg_window\[190\] net933
+ vssd1 vssd1 vccd1 vccd1 _01434_ sky130_fd_sc_hd__mux2_1
XANTENNA__11830__S net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08222_ _03169_ _03170_ _03171_ _03172_ net681 net699 vssd1 vssd1 vccd1 vccd1 _03173_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__07391__S1 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12865__CLK clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11919__A2 _06248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07048__A1 final_design.data_from_mem\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12041__A1 net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08153_ _01968_ net612 vssd1 vssd1 vccd1 vccd1 _03104_ sky130_fd_sc_hd__nor2_1
XFILLER_0_71_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07104_ final_design.cpu.reg_window\[524\] final_design.cpu.reg_window\[556\] net893
+ vssd1 vssd1 vccd1 vccd1 _02055_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11395__A3 _06079_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12592__A2 net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08084_ _02803_ _03034_ vssd1 vssd1 vccd1 vccd1 _03035_ sky130_fd_sc_hd__nor2_1
XFILLER_0_82_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_941 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07035_ final_design.cpu.reg_window\[910\] final_design.cpu.reg_window\[942\] net906
+ vssd1 vssd1 vccd1 vccd1 _01986_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout1031_A net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12344__A2 net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10355__B2 final_design.data_from_mem\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout491_A net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1859 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07220__A1 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout589_A net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08986_ _03745_ _03746_ vssd1 vssd1 vccd1 vccd1 _03922_ sky130_fd_sc_hd__nor2_1
X_07937_ final_design.cpu.reg_window\[726\] final_design.cpu.reg_window\[758\] net839
+ vssd1 vssd1 vccd1 vccd1 _02888_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_3_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout756_A _01427_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout377_X net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07868_ final_design.cpu.reg_window\[788\] final_design.cpu.reg_window\[820\] net869
+ vssd1 vssd1 vccd1 vccd1 _02819_ sky130_fd_sc_hd__mux2_1
XANTENNA__08586__S net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08181__C1 net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09607_ net262 _04516_ _04522_ _04525_ vssd1 vssd1 vccd1 vccd1 _04526_ sky130_fd_sc_hd__and4_1
X_06819_ _01766_ _01767_ _01768_ _01769_ net778 net795 vssd1 vssd1 vccd1 vccd1 _01770_
+ sky130_fd_sc_hd__mux4_1
X_07799_ net719 _02749_ vssd1 vssd1 vccd1 vccd1 _02750_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout923_A net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout544_X net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08159__S0 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09538_ net549 net548 net546 net545 net454 net464 vssd1 vssd1 vccd1 vccd1 _04457_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__13640__CLK clknet_leaf_40_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09469_ _04385_ _04387_ vssd1 vssd1 vccd1 vccd1 _04388_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout711_X net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12280__A1 net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11740__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11500_ _05840_ _05842_ _06117_ vssd1 vssd1 vccd1 vccd1 _06119_ sky130_fd_sc_hd__nor3_1
X_12480_ _06140_ net342 net330 net2277 vssd1 vssd1 vccd1 vccd1 _01186_ sky130_fd_sc_hd__a22o_1
XANTENNA__13790__CLK clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11431_ net2052 _06017_ net312 vssd1 vssd1 vccd1 vccd1 _00328_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_1873 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14150_ clknet_leaf_15_clk _01324_ net1107 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.data_to_VGA\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_62_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11362_ net656 _06048_ _06050_ vssd1 vssd1 vccd1 vccd1 _06051_ sky130_fd_sc_hd__or3_1
XFILLER_0_22_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06798__B1 net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11791__B1 net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13101_ clknet_leaf_45_clk _00332_ net1202 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[89\]
+ sky130_fd_sc_hd__dfrtp_1
X_10313_ final_design.VGA_data_control.state\[0\] net1039 final_design.VGA_data_control.state\[1\]
+ vssd1 vssd1 vccd1 vccd1 _05166_ sky130_fd_sc_hd__a21o_2
XFILLER_0_0_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14081_ clknet_leaf_24_clk _01278_ net1161 vssd1 vssd1 vccd1 vccd1 final_design.reqhand.instruction\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13020__CLK clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14146__CLK clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11293_ net433 net575 _05990_ net317 net1646 vssd1 vssd1 vccd1 vccd1 _00292_ sky130_fd_sc_hd__a32o_1
XANTENNA__12335__A2 net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13032_ clknet_leaf_35_clk _00263_ net1240 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input52_A mem_adr_start[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10244_ final_design.uart.BAUD_counter\[16\] _05114_ net798 vssd1 vssd1 vccd1 vccd1
+ _05116_ sky130_fd_sc_hd__o21ai_1
XANTENNA__11695__B net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10346__B2 final_design.data_from_mem\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11543__B1 net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1101 net1105 vssd1 vssd1 vccd1 vccd1 net1101 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_24_1478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1112 net1115 vssd1 vssd1 vccd1 vccd1 net1112 sky130_fd_sc_hd__buf_2
X_10175_ final_design.uart.bits_received\[1\] final_design.uart.bits_received\[2\]
+ _05064_ vssd1 vssd1 vccd1 vccd1 _05065_ sky130_fd_sc_hd__nor3_1
Xfanout1123 net1127 vssd1 vssd1 vccd1 vccd1 net1123 sky130_fd_sc_hd__clkbuf_4
Xfanout1134 net1135 vssd1 vssd1 vccd1 vccd1 net1134 sky130_fd_sc_hd__clkbuf_4
Xfanout1145 net1149 vssd1 vssd1 vccd1 vccd1 net1145 sky130_fd_sc_hd__clkbuf_4
XANTENNA__13170__CLK clknet_leaf_39_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12099__A1 net240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1156 net1157 vssd1 vssd1 vccd1 vccd1 net1156 sky130_fd_sc_hd__clkbuf_4
Xfanout1167 net100 vssd1 vssd1 vccd1 vccd1 net1167 sky130_fd_sc_hd__buf_4
Xfanout180 _06074_ vssd1 vssd1 vccd1 vccd1 net180 sky130_fd_sc_hd__buf_2
Xfanout1178 net1192 vssd1 vssd1 vccd1 vccd1 net1178 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_76_1833 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout191 _06038_ vssd1 vssd1 vccd1 vccd1 net191 sky130_fd_sc_hd__clkbuf_2
Xfanout1189 net1190 vssd1 vssd1 vccd1 vccd1 net1189 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_57_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13934_ clknet_leaf_45_clk _01165_ net1215 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[922\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12996__RESET_B net1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08496__S net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_1877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13865_ clknet_leaf_33_clk _01096_ net1231 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[853\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_46_clk_X clknet_leaf_46_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12816_ net1347 vssd1 vssd1 vccd1 vccd1 _00257_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_80_2930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13796_ clknet_leaf_51_clk _01027_ net1171 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[784\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_80_2941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12888__CLK clknet_leaf_17_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_2952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12271__A1 net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12747_ final_design.VGA_adr\[4\] net796 vssd1 vssd1 vccd1 vccd1 _06386_ sky130_fd_sc_hd__and2_1
XFILLER_0_45_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12678_ _06326_ net1388 net978 vssd1 vssd1 vccd1 vccd1 _01341_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_13_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11629_ net213 net630 vssd1 vssd1 vccd1 vccd1 _06172_ sky130_fd_sc_hd__and2_1
XFILLER_0_48_1913 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08322__S0 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_2870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_2881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_74_2723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10585__A1 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold606 final_design.cpu.reg_window\[418\] vssd1 vssd1 vccd1 vccd1 net1948 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_55_2100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_2734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11782__B1 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold617 final_design.cpu.reg_window\[981\] vssd1 vssd1 vccd1 vccd1 net1959 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold628 final_design.cpu.reg_window\[747\] vssd1 vssd1 vccd1 vccd1 net1970 sky130_fd_sc_hd__dlygate4sd3_1
Xhold639 final_design.cpu.reg_window\[344\] vssd1 vssd1 vccd1 vccd1 net1981 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_70_2609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13513__CLK clknet_leaf_36_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14207__1265 vssd1 vssd1 vccd1 vccd1 _14207__1265/HI net1265 sky130_fd_sc_hd__conb_1
XANTENNA__10337__B2 final_design.data_from_mem\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08840_ final_design.CPU_instr_adr\[14\] _03790_ vssd1 vssd1 vccd1 vccd1 _03791_
+ sky130_fd_sc_hd__and2_1
X_08771_ _03704_ _03721_ _03703_ vssd1 vssd1 vccd1 vccd1 _03722_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_68_2516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06986__Y _01937_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_2527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11825__S net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_2538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07722_ _02670_ _02671_ vssd1 vssd1 vccd1 vccd1 _02673_ sky130_fd_sc_hd__or2_2
XANTENNA__13663__CLK clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1917 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08702__A1 _03635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07653_ net607 _02602_ _02577_ vssd1 vssd1 vccd1 vccd1 _02604_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_36_1327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06604_ final_design.cpu.reg_window\[796\] final_design.cpu.reg_window\[828\] net946
+ vssd1 vssd1 vccd1 vccd1 _01555_ sky130_fd_sc_hd__mux2_1
X_07584_ final_design.cpu.reg_window\[799\] final_design.cpu.reg_window\[831\] net859
+ vssd1 vssd1 vccd1 vccd1 _02535_ sky130_fd_sc_hd__mux2_1
XANTENNA__14019__CLK clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09323_ _04241_ vssd1 vssd1 vccd1 vccd1 _04242_ sky130_fd_sc_hd__inv_2
X_06535_ _01456_ _01465_ _01474_ vssd1 vssd1 vccd1 vccd1 _01486_ sky130_fd_sc_hd__nor3_2
XANTENNA__12262__A1 net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09254_ _02574_ _02606_ _04171_ _02641_ _02575_ vssd1 vssd1 vccd1 vccd1 _04173_ sky130_fd_sc_hd__a311o_1
XANTENNA__06654__S net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06466_ final_design.reqhand.instruction\[17\] net971 vssd1 vssd1 vccd1 vccd1 _01417_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_35_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08205_ final_design.cpu.reg_window\[590\] final_design.cpu.reg_window\[622\] net813
+ vssd1 vssd1 vccd1 vccd1 _03156_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11132__Y _05847_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13043__CLK clknet_leaf_40_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09185_ _04102_ _04103_ vssd1 vssd1 vccd1 vccd1 _04104_ sky130_fd_sc_hd__nand2_1
XANTENNA__14169__CLK clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout504_A net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08154__B net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10025__B1 net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08136_ final_design.cpu.reg_window\[717\] final_design.cpu.reg_window\[749\] net854
+ vssd1 vssd1 vccd1 vccd1 _03087_ sky130_fd_sc_hd__mux2_1
XANTENNA__10576__A1 net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09430__A2 _04348_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10576__B2 net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11796__A net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07441__A1 final_design.data_from_mem\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08067_ final_design.cpu.reg_window\[594\] final_design.cpu.reg_window\[626\] net844
+ vssd1 vssd1 vccd1 vccd1 _03018_ sky130_fd_sc_hd__mux2_1
XANTENNA__12391__S net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13193__CLK clknet_leaf_36_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07018_ net543 _01968_ vssd1 vssd1 vccd1 vccd1 _01969_ sky130_fd_sc_hd__and2_1
XANTENNA__10328__B2 final_design.data_from_mem\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout873_A _01818_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout494_X net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout661_X net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08969_ net625 _03906_ vssd1 vssd1 vccd1 vccd1 _03907_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout759_X net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11289__C1 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11980_ _06182_ net283 net405 net1688 vssd1 vssd1 vccd1 vccd1 _00713_ sky130_fd_sc_hd__a22o_1
XANTENNA__06829__S net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09497__A2 _04086_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10931_ net959 _05656_ _05659_ net956 vssd1 vssd1 vccd1 vccd1 _05660_ sky130_fd_sc_hd__o22a_1
XFILLER_0_19_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10862_ _05569_ _05586_ _05587_ _05592_ vssd1 vssd1 vccd1 vccd1 _05594_ sky130_fd_sc_hd__or4_1
X_13650_ clknet_leaf_38_clk _00881_ net1189 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[638\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1883 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12601_ net1480 net996 net982 final_design.data_from_mem\[19\] vssd1 vssd1 vccd1
+ vccd1 _01294_ sky130_fd_sc_hd__a22o_1
XFILLER_0_71_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12253__A1 net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13581_ clknet_leaf_53_clk _00812_ net1185 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[569\]
+ sky130_fd_sc_hd__dfrtp_1
X_10793_ net76 net1044 vssd1 vssd1 vccd1 vccd1 _05528_ sky130_fd_sc_hd__and2_1
XANTENNA__11470__S net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11323__X _06017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12532_ _06195_ net349 net323 net1991 vssd1 vssd1 vccd1 vccd1 _01236_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_26_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12463_ net1795 net177 net336 vssd1 vssd1 vccd1 vccd1 _01170_ sky130_fd_sc_hd__mux2_1
XANTENNA__08304__S0 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14202_ net1260 vssd1 vssd1 vccd1 vccd1 gpio_oeb[14] sky130_fd_sc_hd__buf_2
XFILLER_0_69_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11414_ net2178 net239 net311 vssd1 vssd1 vccd1 vccd1 _00311_ sky130_fd_sc_hd__mux2_1
XANTENNA__12556__A2 net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12394_ net1835 net179 net270 vssd1 vssd1 vccd1 vccd1 _01105_ sky130_fd_sc_hd__mux2_1
XANTENNA__13536__CLK clknet_leaf_11_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14133_ clknet_leaf_18_clk final_design.vga.h_next_count\[2\] net1114 vssd1 vssd1
+ vccd1 vccd1 final_design.VGA_data_control.h_count\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_65_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13195__RESET_B net1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11345_ _01691_ net641 _06035_ net643 net656 vssd1 vssd1 vccd1 vccd1 _06036_ sky130_fd_sc_hd__a221o_1
XFILLER_0_39_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07395__S net913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07983__A2 _02929_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14064_ clknet_leaf_15_clk _00026_ net1091 vssd1 vssd1 vccd1 vccd1 final_design.uart.BAUD_counter\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_11276_ net738 _03927_ vssd1 vssd1 vccd1 vccd1 _05975_ sky130_fd_sc_hd__nand2_1
XFILLER_0_43_1843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10319__B2 final_design.data_from_mem\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13015_ clknet_leaf_5_clk _00246_ net1081 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_10227_ _05104_ _05105_ vssd1 vssd1 vccd1 vccd1 _00037_ sky130_fd_sc_hd__nor2_1
XANTENNA__13686__CLK clknet_leaf_61_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10158_ net1048 final_design.VGA_data_control.h_count\[5\] _05050_ vssd1 vssd1 vccd1
+ vccd1 _05054_ sky130_fd_sc_hd__and3_1
Xhold3 net116 vssd1 vssd1 vccd1 vccd1 net1345 sky130_fd_sc_hd__dlygate4sd3_1
X_10089_ final_design.vga.v_current_state\[1\] final_design.vga.v_current_state\[0\]
+ vssd1 vssd1 vccd1 vccd1 _05005_ sky130_fd_sc_hd__nor2_1
XFILLER_0_55_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_11_clk_A clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07424__A net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13917_ clknet_leaf_1_clk _01148_ net1078 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[905\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_77_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_911 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13848_ clknet_leaf_64_clk _01079_ net1076 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[836\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12244__A1 net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13066__CLK clknet_leaf_60_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_26_clk_A clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13779_ clknet_leaf_39_clk _01010_ net1207 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[767\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09645__C1 net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1792 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_76_2807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12547__A2 net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold403 final_design.cpu.reg_window\[159\] vssd1 vssd1 vccd1 vccd1 net1745 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold414 final_design.cpu.reg_window\[596\] vssd1 vssd1 vccd1 vccd1 net1756 sky130_fd_sc_hd__dlygate4sd3_1
Xhold425 final_design.cpu.reg_window\[858\] vssd1 vssd1 vccd1 vccd1 net1767 sky130_fd_sc_hd__dlygate4sd3_1
Xhold436 final_design.cpu.reg_window\[760\] vssd1 vssd1 vccd1 vccd1 net1778 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12903__CLK clknet_leaf_61_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1066 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold447 final_design.cpu.reg_window\[45\] vssd1 vssd1 vccd1 vccd1 net1789 sky130_fd_sc_hd__dlygate4sd3_1
Xhold458 net155 vssd1 vssd1 vccd1 vccd1 net1800 sky130_fd_sc_hd__dlygate4sd3_1
Xhold469 final_design.cpu.reg_window\[779\] vssd1 vssd1 vccd1 vccd1 net1811 sky130_fd_sc_hd__dlygate4sd3_1
X_09941_ _04719_ _04859_ vssd1 vssd1 vccd1 vccd1 _04860_ sky130_fd_sc_hd__nand2_1
XANTENNA_clkload24_A clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout905 net910 vssd1 vssd1 vccd1 vccd1 net905 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_22_1927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout916 net917 vssd1 vssd1 vccd1 vccd1 net916 sky130_fd_sc_hd__buf_2
Xfanout927 net953 vssd1 vssd1 vccd1 vccd1 net927 sky130_fd_sc_hd__buf_2
XFILLER_0_0_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09872_ _03522_ _04087_ net440 _03520_ _04790_ vssd1 vssd1 vccd1 vccd1 _04791_ sky130_fd_sc_hd__a221o_1
Xfanout938 net940 vssd1 vssd1 vccd1 vccd1 net938 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12180__B1 _06270_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout949 net950 vssd1 vssd1 vccd1 vccd1 net949 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_77_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08823_ _03660_ _03773_ _03661_ vssd1 vssd1 vccd1 vccd1 _03774_ sky130_fd_sc_hd__o21a_1
Xhold1103 final_design.cpu.reg_window\[482\] vssd1 vssd1 vccd1 vccd1 net2445 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1114 final_design.cpu.reg_window\[43\] vssd1 vssd1 vccd1 vccd1 net2456 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1125 final_design.cpu.reg_window\[115\] vssd1 vssd1 vccd1 vccd1 net2467 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout287_A _06228_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1136 final_design.cpu.reg_window\[872\] vssd1 vssd1 vccd1 vccd1 net2478 sky130_fd_sc_hd__dlygate4sd3_1
X_08754_ _03703_ _03704_ vssd1 vssd1 vccd1 vccd1 _03705_ sky130_fd_sc_hd__nand2b_1
Xhold1147 final_design.cpu.reg_window\[636\] vssd1 vssd1 vccd1 vccd1 net2489 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1158 final_design.cpu.reg_window\[639\] vssd1 vssd1 vccd1 vccd1 net2500 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1169 final_design.cpu.reg_window\[284\] vssd1 vssd1 vccd1 vccd1 net2511 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_59_1861 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07705_ final_design.cpu.reg_window\[603\] final_design.cpu.reg_window\[635\] net861
+ vssd1 vssd1 vccd1 vccd1 _02656_ sky130_fd_sc_hd__mux2_1
XANTENNA__11286__A2 net235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08685_ _03486_ _03487_ _03520_ _03521_ vssd1 vssd1 vccd1 vccd1 _03636_ sky130_fd_sc_hd__o22a_1
XFILLER_0_68_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout454_A net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13409__CLK clknet_leaf_48_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1196_A net1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07636_ final_design.cpu.reg_window\[156\] final_design.cpu.reg_window\[188\] net860
+ vssd1 vssd1 vccd1 vccd1 _02587_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_0_166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_0_188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12386__S net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12235__A1 net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07567_ final_design.cpu.reg_window\[479\] final_design.cpu.reg_window\[511\] net859
+ vssd1 vssd1 vccd1 vccd1 _02518_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout242_X net242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout621_A _02507_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout719_A net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09306_ net472 net463 net527 vssd1 vssd1 vccd1 vccd1 _04225_ sky130_fd_sc_hd__a21oi_1
X_06518_ _01466_ _01467_ vssd1 vssd1 vccd1 vccd1 _01469_ sky130_fd_sc_hd__nor2_1
XFILLER_0_76_796 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08165__A net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07498_ _02067_ _02101_ _02446_ _02065_ _02033_ vssd1 vssd1 vccd1 vccd1 _02449_ sky130_fd_sc_hd__o311a_1
XANTENNA__13559__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09237_ _04141_ _04155_ vssd1 vssd1 vccd1 vccd1 _04156_ sky130_fd_sc_hd__or2_1
X_06449_ final_design.VGA_data_control.v_count\[7\] final_design.VGA_data_control.v_count\[8\]
+ vssd1 vssd1 vccd1 vccd1 _01403_ sky130_fd_sc_hd__nand2_1
X_12801__32 clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 net1342 sky130_fd_sc_hd__inv_2
XFILLER_0_63_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout507_X net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12538__A2 net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09168_ _03631_ net659 vssd1 vssd1 vccd1 vccd1 _04087_ sky130_fd_sc_hd__nor2_4
XTAP_TAPCELL_ROW_40_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11746__A0 net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_40_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08119_ _03067_ _03069_ vssd1 vssd1 vccd1 vccd1 _03070_ sky130_fd_sc_hd__nor2_1
X_09099_ final_design.CPU_instr_adr\[3\] net1018 vssd1 vssd1 vccd1 vccd1 _04022_ sky130_fd_sc_hd__xor2_1
XANTENNA__11957__C net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08612__B net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11130_ _05842_ _05843_ vssd1 vssd1 vccd1 vccd1 _05845_ sky130_fd_sc_hd__nor2_4
Xhold970 final_design.cpu.reg_window\[287\] vssd1 vssd1 vccd1 vccd1 net2312 sky130_fd_sc_hd__dlygate4sd3_1
Xhold981 final_design.cpu.reg_window\[341\] vssd1 vssd1 vccd1 vccd1 net2323 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout876_X net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11061_ _05763_ _05765_ _05779_ _05782_ vssd1 vssd1 vccd1 vccd1 _05784_ sky130_fd_sc_hd__o211a_1
Xhold992 final_design.cpu.reg_window\[54\] vssd1 vssd1 vccd1 vccd1 net2334 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10012_ net470 _04930_ vssd1 vssd1 vccd1 vccd1 _04931_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_34_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08914__B2 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11465__S net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input15_A DAT_I[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13089__CLK clknet_leaf_47_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11963_ _06165_ net282 net405 net1827 vssd1 vssd1 vccd1 vccd1 _00696_ sky130_fd_sc_hd__a22o_1
XFILLER_0_73_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13702_ clknet_leaf_51_clk _00933_ net1172 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[690\]
+ sky130_fd_sc_hd__dfrtp_1
X_10914_ net50 _05642_ vssd1 vssd1 vccd1 vccd1 _05644_ sky130_fd_sc_hd__nor2_1
X_11894_ net219 net1997 net272 vssd1 vssd1 vccd1 vccd1 _00636_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_15_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10845_ _05566_ _05575_ _05577_ net46 vssd1 vssd1 vccd1 vccd1 _05578_ sky130_fd_sc_hd__a31oi_2
XTAP_TAPCELL_ROW_15_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13633_ clknet_leaf_46_clk _00864_ net1203 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[621\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_15_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14206__1264 vssd1 vssd1 vccd1 vccd1 _14206__1264/HI net1264 sky130_fd_sc_hd__conb_1
XFILLER_0_55_936 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10776_ _05510_ _05511_ _05486_ vssd1 vssd1 vccd1 vccd1 _05512_ sky130_fd_sc_hd__o21bai_1
X_13564_ clknet_leaf_3_clk _00795_ net1067 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[552\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11985__B1 net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09642__A2 _04559_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12515_ _06177_ net351 net329 net1770 vssd1 vssd1 vccd1 vccd1 _01220_ sky130_fd_sc_hd__a22o_1
XANTENNA__07653__A1 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13495_ clknet_leaf_6_clk _00726_ net1130 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[483\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12926__CLK clknet_leaf_49_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12529__A2 net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12446_ net1874 net207 net334 vssd1 vssd1 vccd1 vccd1 _01153_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07405__B2 net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12377_ net1574 net210 net271 vssd1 vssd1 vccd1 vccd1 _01088_ sky130_fd_sc_hd__mux2_1
XANTENNA__09618__B net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08602__B1 _03524_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14116_ clknet_leaf_15_clk _01313_ net1095 vssd1 vssd1 vccd1 vccd1 final_design.reqhand.data_from_UART\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_11328_ final_design.data_from_mem\[22\] net235 net233 vssd1 vssd1 vccd1 vccd1 _06021_
+ sky130_fd_sc_hd__a21o_2
XANTENNA__10960__A1 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10960__B2 net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14047_ clknet_leaf_16_clk _00008_ net1094 vssd1 vssd1 vccd1 vccd1 final_design.uart.BAUD_counter\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_11259_ final_design.data_from_mem\[14\] _05914_ _05917_ vssd1 vssd1 vccd1 vccd1
+ _05960_ sky130_fd_sc_hd__a21o_1
XFILLER_0_24_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11883__B _06116_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12331__Y _06277_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08118__C1 net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08470_ net529 net495 vssd1 vssd1 vccd1 vccd1 _03421_ sky130_fd_sc_hd__or2_2
XFILLER_0_82_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07421_ final_design.cpu.reg_window\[193\] final_design.cpu.reg_window\[225\] net916
+ vssd1 vssd1 vccd1 vccd1 _02372_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13701__CLK clknet_leaf_49_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12217__A1 net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08516__S0 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12768__A2 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07352_ final_design.cpu.reg_window\[451\] final_design.cpu.reg_window\[483\] net908
+ vssd1 vssd1 vccd1 vccd1 _02303_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11976__B1 net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07283_ final_design.cpu.reg_window\[518\] final_design.cpu.reg_window\[550\] net904
+ vssd1 vssd1 vccd1 vccd1 _02234_ sky130_fd_sc_hd__mux2_1
XANTENNA__13851__CLK clknet_leaf_65_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09022_ _02067_ _02447_ _03953_ vssd1 vssd1 vccd1 vccd1 _03954_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_31_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11728__B1 net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09397__A1 net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold200 final_design.VGA_data_control.ready_data\[20\] vssd1 vssd1 vccd1 vccd1 net1542
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold211 final_design.cpu.reg_window\[847\] vssd1 vssd1 vccd1 vccd1 net1553 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout202_A _05996_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold222 final_design.cpu.reg_window\[528\] vssd1 vssd1 vccd1 vccd1 net1564 sky130_fd_sc_hd__dlygate4sd3_1
Xhold233 final_design.cpu.reg_window\[209\] vssd1 vssd1 vccd1 vccd1 net1575 sky130_fd_sc_hd__dlygate4sd3_1
Xhold244 final_design.cpu.reg_window\[463\] vssd1 vssd1 vccd1 vccd1 net1586 sky130_fd_sc_hd__dlygate4sd3_1
Xhold255 final_design.cpu.reg_window\[726\] vssd1 vssd1 vccd1 vccd1 net1597 sky130_fd_sc_hd__dlygate4sd3_1
Xhold266 final_design.cpu.reg_window\[900\] vssd1 vssd1 vccd1 vccd1 net1608 sky130_fd_sc_hd__dlygate4sd3_1
Xhold277 final_design.cpu.reg_window\[132\] vssd1 vssd1 vccd1 vccd1 net1619 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_1871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold288 final_design.cpu.reg_window\[234\] vssd1 vssd1 vccd1 vccd1 net1630 sky130_fd_sc_hd__dlygate4sd3_1
Xhold299 final_design.cpu.reg_window\[467\] vssd1 vssd1 vccd1 vccd1 net1641 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout702 _01752_ vssd1 vssd1 vccd1 vccd1 net702 sky130_fd_sc_hd__buf_4
XFILLER_0_22_1713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09924_ net263 _04837_ _04841_ _04842_ vssd1 vssd1 vccd1 vccd1 _04843_ sky130_fd_sc_hd__and4_1
Xfanout713 net714 vssd1 vssd1 vccd1 vccd1 net713 sky130_fd_sc_hd__clkbuf_4
Xfanout724 _01688_ vssd1 vssd1 vccd1 vccd1 net724 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_0_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout735 net736 vssd1 vssd1 vccd1 vccd1 net735 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07763__S net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1209_A net1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout746 _01438_ vssd1 vssd1 vccd1 vccd1 net746 sky130_fd_sc_hd__clkbuf_4
XANTENNA_input7_A DAT_I[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09855_ _03627_ _04266_ vssd1 vssd1 vccd1 vccd1 _04774_ sky130_fd_sc_hd__nand2_1
Xfanout757 net759 vssd1 vssd1 vccd1 vccd1 net757 sky130_fd_sc_hd__buf_2
XANTENNA__11900__A0 net206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout768 net771 vssd1 vssd1 vccd1 vccd1 net768 sky130_fd_sc_hd__buf_4
XANTENNA_fanout571_A _05868_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout779 _01422_ vssd1 vssd1 vccd1 vccd1 net779 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout669_A net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08806_ _03754_ _03756_ vssd1 vssd1 vccd1 vccd1 _03757_ sky130_fd_sc_hd__nor2_1
XANTENNA__13231__CLK clknet_leaf_43_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10042__X _04961_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06998_ final_design.cpu.reg_window\[15\] final_design.cpu.reg_window\[47\] net888
+ vssd1 vssd1 vccd1 vccd1 _01949_ sky130_fd_sc_hd__mux2_1
X_09786_ _03391_ _04149_ _04150_ vssd1 vssd1 vccd1 vccd1 _04705_ sky130_fd_sc_hd__o21ai_1
X_08737_ final_design.CPU_instr_adr\[11\] _02097_ vssd1 vssd1 vccd1 vccd1 _03688_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_55_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_65_clk clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_65_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout836_A net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_4_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08668_ _01463_ net740 _03618_ _01486_ vssd1 vssd1 vccd1 vccd1 _03619_ sky130_fd_sc_hd__a31o_1
XANTENNA__13381__CLK clknet_leaf_52_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09872__A2 _04087_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07619_ net877 _02569_ _02558_ _02557_ vssd1 vssd1 vccd1 vccd1 _02570_ sky130_fd_sc_hd__o2bb2a_2
X_08599_ net874 _03542_ _03548_ _03535_ _03536_ vssd1 vssd1 vccd1 vccd1 _03550_ sky130_fd_sc_hd__a32o_4
XANTENNA__12949__CLK clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10630_ _05368_ _05369_ _05349_ vssd1 vssd1 vccd1 vccd1 _05373_ sky130_fd_sc_hd__a21o_1
XFILLER_0_14_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_27_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_1875 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_722 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09085__B1 net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11967__B1 net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10561_ net1005 _05304_ _05307_ vssd1 vssd1 vccd1 vccd1 _05308_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_42_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12300_ net1636 net227 net365 vssd1 vssd1 vccd1 vccd1 _01014_ sky130_fd_sc_hd__mux2_1
XANTENNA__07938__S net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13280_ clknet_leaf_10_clk _00511_ net1101 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[268\]
+ sky130_fd_sc_hd__dfrtp_1
X_10492_ net964 _05241_ vssd1 vssd1 vccd1 vccd1 _05242_ sky130_fd_sc_hd__nand2_1
XFILLER_0_23_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08623__A _02185_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12231_ _06161_ net500 net373 net1774 vssd1 vssd1 vccd1 vccd1 _00948_ sky130_fd_sc_hd__a22o_1
XFILLER_0_62_1504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11195__A1 _04723_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09483__S1 net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12162_ _06117_ _06260_ vssd1 vssd1 vccd1 vccd1 _06269_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_9_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11113_ final_design.uart.bits_received\[0\] final_design.uart.bits_received\[1\]
+ vssd1 vssd1 vccd1 vccd1 _05832_ sky130_fd_sc_hd__nand2_1
X_12093_ net579 _06090_ net511 net394 net2243 vssd1 vssd1 vccd1 vccd1 _00818_ sky130_fd_sc_hd__a32o_1
XFILLER_0_25_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12144__A0 net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11044_ final_design.CPU_instr_adr\[28\] net1001 _05767_ net1042 net963 vssd1 vssd1
+ vccd1 vccd1 _05768_ sky130_fd_sc_hd__o221a_1
XFILLER_0_36_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09173__B net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12447__A1 net206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13724__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_1622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12995_ net1326 _00226_ net1194 vssd1 vssd1 vccd1 vccd1 final_design.CPU_instr_adr\[15\]
+ sky130_fd_sc_hd__dfrtp_4
Xclkbuf_leaf_56_clk clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_56_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_59_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07549__S1 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11946_ _06147_ net283 net409 net2079 vssd1 vssd1 vccd1 vccd1 _00681_ sky130_fd_sc_hd__a22o_1
XFILLER_0_52_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11877_ _06111_ net291 net520 net2049 vssd1 vssd1 vccd1 vccd1 _00621_ sky130_fd_sc_hd__a22o_1
XANTENNA__13874__CLK clknet_leaf_44_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13616_ clknet_leaf_36_clk _00847_ net1237 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[604\]
+ sky130_fd_sc_hd__dfrtp_1
X_10828_ _05559_ _05561_ vssd1 vssd1 vccd1 vccd1 _05562_ sky130_fd_sc_hd__or2_1
XFILLER_0_28_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08009__S net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13547_ clknet_leaf_52_clk _00778_ net1182 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[535\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_1773 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10759_ _05483_ _05493_ _05495_ net42 vssd1 vssd1 vccd1 vccd1 _05496_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_55_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13104__CLK clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13478_ clknet_leaf_51_clk _00709_ net1169 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[466\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12792__23 clknet_leaf_27_clk vssd1 vssd1 vccd1 vccd1 net1333 sky130_fd_sc_hd__inv_2
X_12429_ final_design.cpu.reg_window\[895\] net341 vssd1 vssd1 vccd1 vccd1 _06281_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_65_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_983 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09474__S1 net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07970_ final_design.cpu.reg_window\[785\] final_design.cpu.reg_window\[817\] net845
+ vssd1 vssd1 vccd1 vccd1 _02921_ sky130_fd_sc_hd__mux2_1
XANTENNA__13254__CLK clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06921_ final_design.cpu.reg_window\[914\] final_design.cpu.reg_window\[946\] net924
+ vssd1 vssd1 vccd1 vccd1 _01872_ sky130_fd_sc_hd__mux2_1
X_09640_ _04486_ _04489_ net479 vssd1 vssd1 vccd1 vccd1 _04559_ sky130_fd_sc_hd__mux2_2
X_06852_ final_design.cpu.reg_window\[852\] final_design.cpu.reg_window\[884\] net950
+ vssd1 vssd1 vccd1 vccd1 _01803_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09651__X _04570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09571_ net472 _04489_ vssd1 vssd1 vccd1 vccd1 _04490_ sky130_fd_sc_hd__nand2_1
X_06783_ final_design.cpu.reg_window\[214\] final_design.cpu.reg_window\[246\] net919
+ vssd1 vssd1 vccd1 vccd1 _01734_ sky130_fd_sc_hd__mux2_1
XANTENNA__10022__B _04940_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_47_clk clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_47_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__11833__S net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08522_ final_design.cpu.reg_window\[898\] final_design.cpu.reg_window\[930\] net832
+ vssd1 vssd1 vccd1 vccd1 _03473_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09854__A2 _04406_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08453_ final_design.cpu.reg_window\[836\] final_design.cpu.reg_window\[868\] net819
+ vssd1 vssd1 vccd1 vccd1 _03404_ sky130_fd_sc_hd__mux2_1
X_07404_ _02349_ _02354_ net752 vssd1 vssd1 vccd1 vccd1 _02355_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08384_ final_design.cpu.reg_window\[6\] final_design.cpu.reg_window\[38\] net820
+ vssd1 vssd1 vccd1 vccd1 _03335_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11949__B1 net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07335_ final_design.cpu.reg_window\[900\] final_design.cpu.reg_window\[932\] net900
+ vssd1 vssd1 vccd1 vccd1 _02286_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12610__B2 final_design.data_from_mem\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1061_A net1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout417_A net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1159_A net1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07758__S net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07266_ final_design.cpu.reg_window\[262\] final_design.cpu.reg_window\[294\] net912
+ vssd1 vssd1 vccd1 vccd1 _02217_ sky130_fd_sc_hd__mux2_1
XANTENNA__11788__B net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09005_ final_design.CPU_instr_adr\[14\] _03790_ vssd1 vssd1 vccd1 vccd1 _03939_
+ sky130_fd_sc_hd__nor2_1
X_07197_ net749 _02147_ vssd1 vssd1 vccd1 vccd1 _02148_ sky130_fd_sc_hd__or2_1
XANTENNA__11177__A1 final_design.data_from_mem\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout786_A net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout510 net511 vssd1 vssd1 vccd1 vccd1 net510 sky130_fd_sc_hd__clkbuf_4
Xfanout521 net522 vssd1 vssd1 vccd1 vccd1 net521 sky130_fd_sc_hd__clkbuf_8
Xfanout532 _02239_ vssd1 vssd1 vccd1 vccd1 net532 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_50_1906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09907_ _04072_ _04824_ _04810_ net728 vssd1 vssd1 vccd1 vccd1 _04826_ sky130_fd_sc_hd__o211a_1
XFILLER_0_61_1592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14205__1263 vssd1 vssd1 vccd1 vccd1 _14205__1263/HI net1263 sky130_fd_sc_hd__conb_1
XANTENNA__13747__CLK clknet_leaf_39_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12677__B2 final_design.data_from_mem\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout554 _06238_ vssd1 vssd1 vccd1 vccd1 net554 sky130_fd_sc_hd__buf_2
XANTENNA_fanout574_X net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout565 net571 vssd1 vssd1 vccd1 vccd1 net565 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_50_1928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout576 _05868_ vssd1 vssd1 vccd1 vccd1 net576 sky130_fd_sc_hd__buf_2
X_09838_ net490 _04435_ _04756_ vssd1 vssd1 vccd1 vccd1 _04757_ sky130_fd_sc_hd__a21o_1
Xfanout587 _05868_ vssd1 vssd1 vccd1 vccd1 net587 sky130_fd_sc_hd__buf_2
Xfanout598 net601 vssd1 vssd1 vccd1 vccd1 net598 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_77_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09769_ _03588_ net443 net439 _03587_ vssd1 vssd1 vccd1 vccd1 _04688_ sky130_fd_sc_hd__o22a_1
XFILLER_0_77_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_38_clk clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_38_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout839_X net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11743__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11800_ net2475 net413 _06236_ net430 vssd1 vssd1 vccd1 vccd1 _00553_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_1_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09721__B net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13897__CLK clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_48_1846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11731_ net178 net628 vssd1 vssd1 vccd1 vccd1 _06224_ sky130_fd_sc_hd__and2_1
XANTENNA__11652__A2 net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13127__CLK clknet_leaf_62_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11662_ net435 net586 _06188_ net300 net1901 vssd1 vssd1 vccd1 vccd1 _00463_ sky130_fd_sc_hd__a32o_1
XFILLER_0_14_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13401_ clknet_leaf_56_clk _00632_ net1146 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[389\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_64_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10613_ final_design.CPU_instr_adr\[8\] _03988_ net1058 vssd1 vssd1 vccd1 vccd1 _05357_
+ sky130_fd_sc_hd__mux2_1
X_11593_ net585 net424 _06152_ net304 net1836 vssd1 vssd1 vccd1 vccd1 _00430_ sky130_fd_sc_hd__a32o_1
XANTENNA__12601__B2 final_design.data_from_mem\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11331__X _06024_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input82_A memory_size[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10544_ net94 final_design.VGA_adr\[2\] _05289_ vssd1 vssd1 vccd1 vccd1 _05291_ sky130_fd_sc_hd__and3_1
XANTENNA__07703__S1 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13332_ clknet_leaf_8_clk _00563_ net1151 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[320\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_68_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10475_ net79 net958 net955 final_design.CPU_instr_adr\[1\] vssd1 vssd1 vccd1 vccd1
+ _05226_ sky130_fd_sc_hd__o22a_1
XANTENNA__13277__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13263_ clknet_leaf_43_clk _00494_ net1218 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[251\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09168__B net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11168__A1 final_design.data_from_mem\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08072__B net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12214_ net574 _06142_ net509 net379 net1902 vssd1 vssd1 vccd1 vccd1 _00932_ sky130_fd_sc_hd__a32o_1
X_13194_ clknet_leaf_61_clk _00425_ net1136 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[182\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_output169_A net169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12145_ net205 net2290 net384 vssd1 vssd1 vccd1 vccd1 _00866_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12076_ net2304 net392 net498 _05966_ vssd1 vssd1 vccd1 vccd1 _00801_ sky130_fd_sc_hd__a22o_1
XFILLER_0_60_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11027_ net1003 _05750_ _05751_ net1033 net1376 vssd1 vssd1 vccd1 vccd1 _00200_ sky130_fd_sc_hd__a32o_1
XFILLER_0_75_1717 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_29_clk clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_29_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__09190__Y _04109_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12978_ clknet_leaf_19_clk _00003_ net1156 vssd1 vssd1 vccd1 vccd1 wb_manage.curr_state\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_73_1463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08195__S1 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11929_ _06131_ net280 net408 net2002 vssd1 vssd1 vccd1 vccd1 _00665_ sky130_fd_sc_hd__a22o_1
XFILLER_0_73_1496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_2382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_2393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10851__B1 net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_2246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14052__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_2257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_17 _06228_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_2268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12199__A3 net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_28 _06257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07120_ final_design.cpu.reg_window\[395\] final_design.cpu.reg_window\[427\] net915
+ vssd1 vssd1 vccd1 vccd1 _02071_ sky130_fd_sc_hd__mux2_1
X_07051_ _01996_ _02000_ vssd1 vssd1 vccd1 vccd1 _02002_ sky130_fd_sc_hd__xnor2_2
XTAP_TAPCELL_ROW_11_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput102 net102 vssd1 vssd1 vccd1 vccd1 ADR_O[10] sky130_fd_sc_hd__clkbuf_4
XANTENNA__12356__B1 net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09793__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_2175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput113 net113 vssd1 vssd1 vccd1 vccd1 ADR_O[20] sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_58_2186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput124 net124 vssd1 vssd1 vccd1 vccd1 ADR_O[30] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_23_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_2197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_2039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput135 net135 vssd1 vssd1 vccd1 vccd1 DAT_O[10] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10017__B net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput146 net146 vssd1 vssd1 vccd1 vccd1 DAT_O[20] sky130_fd_sc_hd__clkbuf_4
XANTENNA__11828__S net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput157 net157 vssd1 vssd1 vccd1 vccd1 DAT_O[30] sky130_fd_sc_hd__buf_2
Xoutput168 net168 vssd1 vssd1 vccd1 vccd1 SEL_O[2] sky130_fd_sc_hd__buf_2
XANTENNA__06586__A1 final_design.data_from_mem\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10382__A2 net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08710__B _01599_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06511__A final_design.data_from_mem\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07953_ _01910_ net613 vssd1 vssd1 vccd1 vccd1 _02904_ sky130_fd_sc_hd__nor2_1
XANTENNA__12659__B2 final_design.data_from_mem\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06904_ net548 _01854_ vssd1 vssd1 vccd1 vccd1 _01855_ sky130_fd_sc_hd__and2_1
X_07884_ net605 _02830_ _02805_ _01815_ vssd1 vssd1 vccd1 vccd1 _02835_ sky130_fd_sc_hd__o211a_1
XANTENNA__11331__A1 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09381__X _04300_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09623_ _04536_ _04537_ _04538_ _04534_ vssd1 vssd1 vccd1 vccd1 _04542_ sky130_fd_sc_hd__a31o_1
X_06835_ final_design.reqhand.instruction\[21\] net969 vssd1 vssd1 vccd1 vccd1 _01786_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_78_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11882__A2 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06766_ net886 _01710_ _01716_ _01703_ _01704_ vssd1 vssd1 vccd1 vccd1 _01717_ sky130_fd_sc_hd__a32oi_4
X_09554_ net448 _04472_ _04470_ vssd1 vssd1 vccd1 vccd1 _04473_ sky130_fd_sc_hd__o21ai_1
XANTENNA__09288__B1 _03524_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11095__B1 net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08505_ net595 _03450_ _03452_ _02326_ vssd1 vssd1 vccd1 vccd1 _03456_ sky130_fd_sc_hd__o211ai_1
X_06697_ final_design.cpu.reg_window\[921\] final_design.cpu.reg_window\[953\] net933
+ vssd1 vssd1 vccd1 vccd1 _01648_ sky130_fd_sc_hd__mux2_1
X_09485_ _02502_ net458 _04203_ net462 vssd1 vssd1 vccd1 vccd1 _04404_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout534_A _02184_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08436_ net610 _03384_ _03385_ net530 vssd1 vssd1 vccd1 vccd1 _03387_ sky130_fd_sc_hd__a211oi_1
XANTENNA__11799__A net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08367_ final_design.cpu.reg_window\[519\] final_design.cpu.reg_window\[551\] net806
+ vssd1 vssd1 vccd1 vccd1 _03318_ sky130_fd_sc_hd__mux2_1
XANTENNA__12394__S net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10907__S net1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout701_A _01752_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout322_X net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11398__A1 net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12595__B1 net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1255 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07318_ net531 _02267_ vssd1 vssd1 vccd1 vccd1 _02269_ sky130_fd_sc_hd__nand2_1
XFILLER_0_11_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08298_ _03245_ _03246_ _03247_ _03248_ net674 net696 vssd1 vssd1 vccd1 vccd1 _03249_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__07697__S0 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09460__B1 _04378_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07249_ final_design.cpu.reg_window\[839\] final_design.cpu.reg_window\[871\] net900
+ vssd1 vssd1 vccd1 vccd1 _02200_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12347__B1 net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10260_ final_design.uart.BAUD_counter\[22\] _05124_ net797 vssd1 vssd1 vccd1 vccd1
+ _05126_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07449__S0 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout691_X net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11738__S net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout789_X net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10191_ net1052 _01392_ _05080_ vssd1 vssd1 vccd1 vccd1 _00039_ sky130_fd_sc_hd__o21a_1
XFILLER_0_24_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_1075 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10373__A2 net1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout956_X net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout340 net341 vssd1 vssd1 vccd1 vccd1 net340 sky130_fd_sc_hd__clkbuf_8
Xfanout351 net359 vssd1 vssd1 vccd1 vccd1 net351 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09515__A1 net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout362 net363 vssd1 vssd1 vccd1 vccd1 net362 sky130_fd_sc_hd__clkbuf_8
Xfanout373 _06272_ vssd1 vssd1 vccd1 vccd1 net373 sky130_fd_sc_hd__buf_4
X_13950_ clknet_leaf_13_clk _01181_ net1099 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[938\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout384 net385 vssd1 vssd1 vccd1 vccd1 net384 sky130_fd_sc_hd__clkbuf_8
Xfanout395 _06263_ vssd1 vssd1 vccd1 vccd1 net395 sky130_fd_sc_hd__buf_4
X_12901_ clknet_leaf_25_clk _00139_ net1155 vssd1 vssd1 vccd1 vccd1 net167 sky130_fd_sc_hd__dfrtp_2
XANTENNA__11873__A2 net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13881_ clknet_leaf_55_clk _01112_ net1178 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[869\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11473__S net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12832_ net1353 vssd1 vssd1 vccd1 vccd1 _00273_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__14075__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12763_ _06339_ _06392_ vssd1 vssd1 vccd1 vccd1 _06399_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_33_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10833__B1 _04990_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11714_ net435 net586 _06215_ net296 net2061 vssd1 vssd1 vccd1 vccd1 _00488_ sky130_fd_sc_hd__a32o_1
X_12694_ _01369_ final_design.VGA_data_control.v_count\[6\] _06334_ vssd1 vssd1 vccd1
+ vccd1 _06335_ sky130_fd_sc_hd__a21o_1
XANTENNA__06501__A1 net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11645_ net197 net632 vssd1 vssd1 vccd1 vccd1 _06180_ sky130_fd_sc_hd__and2_1
XFILLER_0_25_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_1721 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12586__B1 net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09179__A _02502_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput15 DAT_I[21] vssd1 vssd1 vccd1 vccd1 net15 sky130_fd_sc_hd__clkbuf_1
Xinput26 DAT_I[31] vssd1 vssd1 vccd1 vccd1 net26 sky130_fd_sc_hd__clkbuf_1
X_11576_ net199 net635 vssd1 vssd1 vccd1 vccd1 _06144_ sky130_fd_sc_hd__and2_1
XANTENNA_clkbuf_leaf_5_clk_X clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08083__A _01815_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput37 mem_adr_start[10] vssd1 vssd1 vccd1 vccd1 net37 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_1765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput48 mem_adr_start[20] vssd1 vssd1 vccd1 vccd1 net48 sky130_fd_sc_hd__clkbuf_1
Xinput59 mem_adr_start[30] vssd1 vssd1 vccd1 vccd1 net59 sky130_fd_sc_hd__clkbuf_1
X_13315_ clknet_leaf_1_clk _00546_ net1072 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[303\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10527_ _05273_ _05274_ vssd1 vssd1 vccd1 vccd1 _05275_ sky130_fd_sc_hd__nor2_1
XANTENNA__06804__A2 _01498_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12338__B1 net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13246_ clknet_leaf_13_clk _00477_ net1099 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[234\]
+ sky130_fd_sc_hd__dfrtp_1
X_10458_ _02570_ net592 vssd1 vssd1 vccd1 vccd1 _05213_ sky130_fd_sc_hd__nor2_1
XANTENNA__11010__B1 _04990_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_2651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13177_ clknet_leaf_59_clk _00408_ net1142 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[165\]
+ sky130_fd_sc_hd__dfrtp_1
X_10389_ net801 net1002 _05175_ net1029 net2551 vssd1 vssd1 vccd1 vccd1 _00138_ sky130_fd_sc_hd__a32o_1
XANTENNA__10364__A2 net1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_2673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11561__A1 net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12128_ final_design.cpu.reg_window\[608\] net385 vssd1 vssd1 vccd1 vccd1 _06267_
+ sky130_fd_sc_hd__and2_1
XANTENNA__08022__S net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08309__A2 _03257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_13 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12059_ _05840_ _05841_ vssd1 vssd1 vccd1 vccd1 _06262_ sky130_fd_sc_hd__nand2_2
XFILLER_0_79_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12510__B1 net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07612__S0 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11864__A2 net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06620_ _01567_ _01570_ vssd1 vssd1 vccd1 vccd1 _01571_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_66_2444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_2308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11077__B1 _04990_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_2319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06551_ final_design.data_from_mem\[31\] net970 _01500_ vssd1 vssd1 vccd1 vccd1 _01502_
+ sky130_fd_sc_hd__o21ai_4
XANTENNA__11616__A2 net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1244 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13442__CLK clknet_leaf_11_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09270_ net78 _04188_ vssd1 vssd1 vccd1 vccd1 _04189_ sky130_fd_sc_hd__or2_2
X_06482_ final_design.cpu.reg_window\[222\] final_design.cpu.reg_window\[254\] net933
+ vssd1 vssd1 vccd1 vccd1 _01433_ sky130_fd_sc_hd__mux2_1
X_08221_ final_design.cpu.reg_window\[395\] final_design.cpu.reg_window\[427\] net835
+ vssd1 vssd1 vccd1 vccd1 _03172_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_1318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14204__1262 vssd1 vssd1 vccd1 vccd1 _14204__1262/HI net1262 sky130_fd_sc_hd__conb_1
XANTENNA__08705__B _01507_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08152_ _03067_ _03069_ _03099_ _03100_ vssd1 vssd1 vccd1 vccd1 _03103_ sky130_fd_sc_hd__o22a_1
XANTENNA__07048__A2 net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09442__B1 _04046_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06506__A final_design.data_from_mem\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13592__CLK clknet_leaf_65_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07103_ final_design.cpu.reg_window\[588\] final_design.cpu.reg_window\[620\] net893
+ vssd1 vssd1 vccd1 vccd1 _02054_ sky130_fd_sc_hd__mux2_1
XANTENNA__11131__B net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08083_ _01815_ _02832_ vssd1 vssd1 vccd1 vccd1 _03034_ sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_9_clk clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_9_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__09239__D _04157_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07034_ final_design.cpu.reg_window\[974\] final_design.cpu.reg_window\[1006\] net897
+ vssd1 vssd1 vccd1 vccd1 _01985_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11001__B1 _05239_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10355__A2 net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08985_ _01942_ _02455_ vssd1 vssd1 vccd1 vccd1 _03921_ sky130_fd_sc_hd__xor2_1
XANTENNA_fanout484_A net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07936_ net715 _02886_ vssd1 vssd1 vccd1 vccd1 _02887_ sky130_fd_sc_hd__nor2_1
XANTENNA__12530__X _06285_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14098__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07771__S net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12501__B1 net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12389__S net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout272_X net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07867_ final_design.cpu.reg_window\[852\] final_design.cpu.reg_window\[884\] net868
+ vssd1 vssd1 vccd1 vccd1 _02818_ sky130_fd_sc_hd__mux2_1
XANTENNA__11855__A2 net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout651_A net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout749_A net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07343__Y _02294_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09606_ _04222_ _04524_ _04218_ vssd1 vssd1 vccd1 vccd1 _04525_ sky130_fd_sc_hd__a21o_1
XFILLER_0_3_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06818_ final_design.cpu.reg_window\[405\] final_design.cpu.reg_window\[437\] net938
+ vssd1 vssd1 vccd1 vccd1 _01769_ sky130_fd_sc_hd__mux2_1
X_07798_ _02745_ _02746_ _02747_ _02748_ net684 net703 vssd1 vssd1 vccd1 vccd1 _02749_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_35_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08159__S1 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09537_ net260 _03589_ _02935_ _02963_ vssd1 vssd1 vccd1 vccd1 _04456_ sky130_fd_sc_hd__o211ai_1
X_06749_ final_design.cpu.reg_window\[215\] final_design.cpu.reg_window\[247\] net929
+ vssd1 vssd1 vccd1 vccd1 _01700_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout916_A net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout537_X net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09468_ _04193_ _04386_ vssd1 vssd1 vccd1 vccd1 _04387_ sky130_fd_sc_hd__and2_1
XANTENNA__09525__A1_N _04116_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08419_ _03366_ _03367_ _03368_ _03369_ net680 net700 vssd1 vssd1 vccd1 vccd1 _03370_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__13935__CLK clknet_leaf_42_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout704_X net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09399_ _02574_ net439 _04314_ _04317_ vssd1 vssd1 vccd1 vccd1 _04318_ sky130_fd_sc_hd__o211a_1
XFILLER_0_69_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_1039 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11430_ net1751 net198 net312 vssd1 vssd1 vccd1 vccd1 _00327_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06416__A net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1885 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11361_ _01630_ net642 _06049_ net644 vssd1 vssd1 vccd1 vccd1 _06050_ sky130_fd_sc_hd__a22o_1
XFILLER_0_46_1104 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06798__A1 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1749 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10312_ net1042 _01395_ vssd1 vssd1 vccd1 vccd1 _05165_ sky130_fd_sc_hd__or2_1
X_13100_ clknet_leaf_46_clk _00331_ net1214 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[88\]
+ sky130_fd_sc_hd__dfrtp_1
X_14080_ clknet_leaf_24_clk _01277_ net1161 vssd1 vssd1 vccd1 vccd1 final_design.reqhand.instruction\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_11292_ net650 net203 vssd1 vssd1 vccd1 vccd1 _05990_ sky130_fd_sc_hd__and2_1
X_10243_ _05114_ _05115_ vssd1 vssd1 vccd1 vccd1 _00012_ sky130_fd_sc_hd__nor2_1
X_13031_ clknet_leaf_62_clk _00262_ net1123 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09446__B _04223_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08095__S0 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11543__A1 net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input45_A mem_adr_start[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10174_ final_design.uart.bits_received\[0\] final_design.uart.bits_received\[3\]
+ vssd1 vssd1 vccd1 vccd1 _05064_ sky130_fd_sc_hd__nand2_1
XANTENNA__13315__CLK clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1102 net1105 vssd1 vssd1 vccd1 vccd1 net1102 sky130_fd_sc_hd__buf_2
Xfanout1113 net1115 vssd1 vssd1 vccd1 vccd1 net1113 sky130_fd_sc_hd__clkbuf_4
Xfanout1124 net1127 vssd1 vssd1 vccd1 vccd1 net1124 sky130_fd_sc_hd__buf_2
Xfanout1135 net1167 vssd1 vssd1 vccd1 vccd1 net1135 sky130_fd_sc_hd__clkbuf_2
Xfanout1146 net1148 vssd1 vssd1 vccd1 vccd1 net1146 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_76_1801 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1157 net1162 vssd1 vssd1 vccd1 vccd1 net1157 sky130_fd_sc_hd__clkbuf_4
Xfanout1168 net1176 vssd1 vssd1 vccd1 vccd1 net1168 sky130_fd_sc_hd__clkbuf_4
Xfanout1179 net1180 vssd1 vssd1 vccd1 vccd1 net1179 sky130_fd_sc_hd__clkbuf_4
Xfanout181 _06074_ vssd1 vssd1 vccd1 vccd1 net181 sky130_fd_sc_hd__clkbuf_2
Xfanout192 _06031_ vssd1 vssd1 vccd1 vccd1 net192 sky130_fd_sc_hd__buf_2
X_13933_ clknet_leaf_53_clk _01164_ net1186 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[921\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_1845 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12299__S net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11846__A2 net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13465__CLK clknet_leaf_56_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_1889 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13864_ clknet_leaf_41_clk _01095_ net1225 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[852\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12815_ net1348 vssd1 vssd1 vccd1 vccd1 _00256_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_80_2920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13795_ clknet_leaf_1_clk _01026_ net1072 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[783\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_80_2931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12746_ _05058_ _06359_ _06366_ _06376_ vssd1 vssd1 vccd1 vccd1 _06385_ sky130_fd_sc_hd__nor4_1
XTAP_TAPCELL_ROW_80_2953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12965__RESET_B net1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07710__A net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07290__A_N _02239_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12677_ final_design.VGA_data_control.ready_data\[26\] net1019 net974 final_design.data_from_mem\[26\]
+ vssd1 vssd1 vccd1 vccd1 _06326_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_13_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12559__B1 net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11628_ net429 net568 _06171_ net299 net1612 vssd1 vssd1 vccd1 vccd1 _00446_ sky130_fd_sc_hd__a32o_1
XANTENNA__12023__A2 net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_78_2860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08322__S1 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11231__B1 net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_2871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11559_ net425 net560 _06135_ net302 net1825 vssd1 vssd1 vccd1 vccd1 _00413_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_78_2882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_2724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10585__A2 _04903_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold607 final_design.cpu.reg_window\[536\] vssd1 vssd1 vccd1 vccd1 net1949 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_55_2101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_2735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold618 final_design.cpu.reg_window\[152\] vssd1 vssd1 vccd1 vccd1 net1960 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold629 final_design.cpu.reg_window\[586\] vssd1 vssd1 vccd1 vccd1 net1971 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_81_1551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_1502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13229_ clknet_leaf_48_clk _00460_ net1202 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[217\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10135__X _05039_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08770_ _03708_ _03720_ _03706_ vssd1 vssd1 vccd1 vccd1 _03721_ sky130_fd_sc_hd__a21o_1
XANTENNA__13808__CLK clknet_leaf_34_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_2517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_2528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_1877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07721_ _02670_ _02671_ vssd1 vssd1 vccd1 vccd1 _02672_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_68_2539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09360__C1 net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07652_ _01570_ net616 vssd1 vssd1 vccd1 vccd1 _02603_ sky130_fd_sc_hd__nor2_1
XFILLER_0_79_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07016__B1_N _01821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06603_ final_design.cpu.reg_window\[860\] final_design.cpu.reg_window\[892\] net951
+ vssd1 vssd1 vccd1 vccd1 _01554_ sky130_fd_sc_hd__mux2_1
XANTENNA__13958__CLK clknet_leaf_51_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07583_ final_design.cpu.reg_window\[863\] final_design.cpu.reg_window\[895\] net859
+ vssd1 vssd1 vccd1 vccd1 _02534_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11841__S net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09322_ net476 _04240_ _04236_ vssd1 vssd1 vccd1 vccd1 _04241_ sky130_fd_sc_hd__a21o_1
XFILLER_0_47_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06534_ _01474_ _01481_ _01482_ vssd1 vssd1 vccd1 vccd1 _01485_ sky130_fd_sc_hd__or3_2
XFILLER_0_76_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11470__A0 net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07620__A _01539_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06465_ net1039 net994 net991 vssd1 vssd1 vccd1 vccd1 _01416_ sky130_fd_sc_hd__or3_1
X_09253_ _02574_ _02606_ _04171_ _02575_ vssd1 vssd1 vccd1 vccd1 _04172_ sky130_fd_sc_hd__a31o_1
XFILLER_0_47_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08204_ final_design.cpu.reg_window\[654\] final_design.cpu.reg_window\[686\] net816
+ vssd1 vssd1 vccd1 vccd1 _03155_ sky130_fd_sc_hd__mux2_1
X_09184_ net614 _03550_ _01536_ _02423_ vssd1 vssd1 vccd1 vccd1 _04103_ sky130_fd_sc_hd__a211o_1
XANTENNA__12014__A2 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09415__B1 _04116_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08135_ final_design.cpu.reg_window\[525\] final_design.cpu.reg_window\[557\] net855
+ vssd1 vssd1 vccd1 vccd1 _03086_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1141_A net1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11773__B2 net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1239_A net1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08066_ final_design.cpu.reg_window\[658\] final_design.cpu.reg_window\[690\] net845
+ vssd1 vssd1 vccd1 vccd1 _03017_ sky130_fd_sc_hd__mux2_1
XANTENNA__11796__B _05869_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07619__X _02570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13338__CLK clknet_leaf_58_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08451__A net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07017_ _01967_ vssd1 vssd1 vccd1 vccd1 _01968_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout699_A net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09813__S1 net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11525__B2 net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout866_A net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13488__CLK clknet_leaf_36_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08968_ _03675_ _03750_ vssd1 vssd1 vccd1 vccd1 _03906_ sky130_fd_sc_hd__xnor2_1
X_07919_ final_design.cpu.reg_window\[342\] final_design.cpu.reg_window\[374\] net839
+ vssd1 vssd1 vccd1 vccd1 _02870_ sky130_fd_sc_hd__mux2_1
X_08899_ net256 _03844_ net1015 vssd1 vssd1 vccd1 vccd1 _03845_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09497__A3 _04411_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10930_ final_design.CPU_instr_adr\[23\] _03870_ net1059 vssd1 vssd1 vccd1 vccd1
+ _05659_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07006__S net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10861_ _05569_ _05586_ _05587_ _05592_ vssd1 vssd1 vccd1 vccd1 _05593_ sky130_fd_sc_hd__o31a_1
XANTENNA_fanout821_X net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11751__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout919_X net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11604__X _06159_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12600_ net1409 net996 net982 final_design.data_from_mem\[18\] vssd1 vssd1 vccd1
+ vccd1 _01293_ sky130_fd_sc_hd__a22o_1
XFILLER_0_13_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13580_ clknet_leaf_47_clk _00811_ net1204 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[568\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_36_1895 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10792_ _04474_ net253 vssd1 vssd1 vccd1 vccd1 _05527_ sky130_fd_sc_hd__nor2_1
XFILLER_0_32_1737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11461__A0 net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12531_ net671 net626 _06268_ net322 net2497 vssd1 vssd1 vccd1 vccd1 _01235_ sky130_fd_sc_hd__a32o_1
XFILLER_0_53_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14113__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08209__A1 net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12005__A2 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12462_ net2062 net179 net336 vssd1 vssd1 vccd1 vccd1 _01169_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14201_ net1259 vssd1 vssd1 vccd1 vccd1 gpio_oeb[13] sky130_fd_sc_hd__buf_2
XANTENNA__08304__S1 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11413_ net1734 net226 net310 vssd1 vssd1 vccd1 vccd1 _00310_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11213__B1 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12393_ net2211 net181 net270 vssd1 vssd1 vccd1 vccd1 _01104_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07676__S net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14132_ clknet_leaf_17_clk final_design.vga.h_next_count\[1\] net1114 vssd1 vssd1
+ vccd1 vccd1 final_design.VGA_data_control.h_count\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_1_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11344_ final_design.data_from_mem\[24\] net235 net233 vssd1 vssd1 vccd1 vccd1 _06035_
+ sky130_fd_sc_hd__a21o_2
XFILLER_0_50_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11198__S net251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14063_ clknet_leaf_15_clk _00025_ net1091 vssd1 vssd1 vccd1 vccd1 final_design.uart.BAUD_counter\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_11275_ net660 _03923_ net733 vssd1 vssd1 vccd1 vccd1 _05974_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_24_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10319__A2 net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11516__A1 net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13014_ clknet_leaf_60_clk _00245_ net1136 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_10226_ final_design.uart.BAUD_counter\[9\] _05103_ net799 vssd1 vssd1 vccd1 vccd1
+ _05105_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_20_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10157_ net1048 _05050_ _05053_ vssd1 vssd1 vccd1 vccd1 final_design.vga.h_next_count\[4\]
+ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_7_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14203__1261 vssd1 vssd1 vccd1 vccd1 _14203__1261/HI net1261 sky130_fd_sc_hd__conb_1
Xhold4 final_design.cpu.reg_window\[11\] vssd1 vssd1 vccd1 vccd1 net1346 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09192__A _03617_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12855__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10088_ _04997_ _05003_ vssd1 vssd1 vccd1 vccd1 _05004_ sky130_fd_sc_hd__nor2_1
XFILLER_0_76_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11227__A net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13916_ clknet_leaf_4_clk _01147_ net1079 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[904\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12492__A2 net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_1528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13847_ clknet_leaf_58_clk _01078_ net1129 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[835\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_945 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13778_ clknet_leaf_39_clk _01009_ net1207 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[766\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09645__B1 _04556_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12729_ _06364_ _06369_ vssd1 vssd1 vccd1 vccd1 _06370_ sky130_fd_sc_hd__nor2_1
XANTENNA__07656__C1 _01566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09919__X _04838_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_2808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11204__B1 net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07586__S net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold404 final_design.cpu.reg_window\[795\] vssd1 vssd1 vccd1 vccd1 net1746 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06490__S net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_856 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09367__A net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold415 final_design.cpu.reg_window\[986\] vssd1 vssd1 vccd1 vccd1 net1757 sky130_fd_sc_hd__dlygate4sd3_1
Xhold426 final_design.cpu.reg_window\[844\] vssd1 vssd1 vccd1 vccd1 net1768 sky130_fd_sc_hd__dlygate4sd3_1
Xhold437 final_design.cpu.reg_window\[841\] vssd1 vssd1 vccd1 vccd1 net1779 sky130_fd_sc_hd__dlygate4sd3_1
Xhold448 final_design.cpu.reg_window\[597\] vssd1 vssd1 vccd1 vccd1 net1790 sky130_fd_sc_hd__dlygate4sd3_1
Xhold459 final_design.cpu.reg_window\[240\] vssd1 vssd1 vccd1 vccd1 net1801 sky130_fd_sc_hd__dlygate4sd3_1
X_09940_ _03391_ _03563_ _04718_ _04046_ vssd1 vssd1 vccd1 vccd1 _04859_ sky130_fd_sc_hd__o31a_1
XFILLER_0_42_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11507__A1 net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout906 net910 vssd1 vssd1 vccd1 vccd1 net906 sky130_fd_sc_hd__clkbuf_4
X_09871_ _03521_ net441 vssd1 vssd1 vccd1 vccd1 _04790_ sky130_fd_sc_hd__nor2_1
Xfanout917 net953 vssd1 vssd1 vccd1 vccd1 net917 sky130_fd_sc_hd__buf_2
Xfanout928 net932 vssd1 vssd1 vccd1 vccd1 net928 sky130_fd_sc_hd__clkbuf_4
XANTENNA_clkload17_A clknet_leaf_17_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout939 net940 vssd1 vssd1 vccd1 vccd1 net939 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11836__S net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08822_ _03663_ _03772_ _03662_ vssd1 vssd1 vccd1 vccd1 _03773_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_29_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1104 final_design.cpu.reg_window\[129\] vssd1 vssd1 vccd1 vccd1 net2446 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10191__B1 _05080_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1115 final_design.cpu.reg_window\[396\] vssd1 vssd1 vccd1 vccd1 net2457 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1126 final_design.cpu.reg_window\[423\] vssd1 vssd1 vccd1 vccd1 net2468 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1137 final_design.cpu.reg_window\[619\] vssd1 vssd1 vccd1 vccd1 net2479 sky130_fd_sc_hd__dlygate4sd3_1
X_08753_ net666 _01659_ final_design.CPU_instr_adr\[5\] vssd1 vssd1 vccd1 vccd1 _03704_
+ sky130_fd_sc_hd__a21o_1
Xhold1148 final_design.cpu.reg_window\[293\] vssd1 vssd1 vccd1 vccd1 net2490 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13780__CLK clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout182_A _06067_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1159 final_design.cpu.reg_window\[486\] vssd1 vssd1 vccd1 vccd1 net2501 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07704_ net719 _02654_ vssd1 vssd1 vccd1 vccd1 _02655_ sky130_fd_sc_hd__nor2_1
XFILLER_0_59_1873 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08684_ _03617_ net594 vssd1 vssd1 vccd1 vccd1 _03635_ sky130_fd_sc_hd__nand2b_2
XANTENNA__12483__A2 net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07635_ final_design.cpu.reg_window\[220\] final_design.cpu.reg_window\[252\] net860
+ vssd1 vssd1 vccd1 vccd1 _02586_ sky130_fd_sc_hd__mux2_1
XANTENNA__10684__A_N net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14136__CLK clknet_leaf_17_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout447_A net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07566_ final_design.cpu.reg_window\[287\] final_design.cpu.reg_window\[319\] net859
+ vssd1 vssd1 vccd1 vccd1 _02517_ sky130_fd_sc_hd__mux2_1
XANTENNA__09636__B1 _04116_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09305_ _02503_ net477 vssd1 vssd1 vccd1 vccd1 _04224_ sky130_fd_sc_hd__nand2_1
X_06517_ _01466_ _01467_ vssd1 vssd1 vccd1 vccd1 _01468_ sky130_fd_sc_hd__or2_4
XFILLER_0_35_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout235_X net235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07497_ _02067_ _02447_ _02065_ vssd1 vssd1 vccd1 vccd1 _02448_ sky130_fd_sc_hd__o21a_1
XFILLER_0_5_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11994__B2 net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09236_ _03261_ _03291_ _03259_ vssd1 vssd1 vccd1 vccd1 _04155_ sky130_fd_sc_hd__a21oi_1
X_06448_ _01397_ _01400_ vssd1 vssd1 vccd1 vccd1 _01402_ sky130_fd_sc_hd__nand2_1
XANTENNA_clkbuf_leaf_30_clk_X clknet_leaf_30_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_17_Right_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13160__CLK clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1833 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout402_X net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09167_ _04054_ net319 vssd1 vssd1 vccd1 vccd1 _04086_ sky130_fd_sc_hd__nand2_2
XANTENNA__08298__S0 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11600__A net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08118_ net599 _03065_ _03041_ net539 vssd1 vssd1 vccd1 vccd1 _03069_ sky130_fd_sc_hd__o211a_1
XFILLER_0_66_1877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_3_0_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09098_ _02432_ _04019_ _04020_ net619 vssd1 vssd1 vccd1 vccd1 _04021_ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_45_clk_X clknet_leaf_45_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08049_ final_design.cpu.reg_window\[402\] final_design.cpu.reg_window\[434\] net844
+ vssd1 vssd1 vccd1 vccd1 _03000_ sky130_fd_sc_hd__mux2_1
Xhold960 final_design.cpu.reg_window\[118\] vssd1 vssd1 vccd1 vccd1 net2302 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold971 final_design.cpu.reg_window\[302\] vssd1 vssd1 vccd1 vccd1 net2313 sky130_fd_sc_hd__dlygate4sd3_1
X_11060_ _05779_ _05782_ _05763_ _05765_ vssd1 vssd1 vccd1 vccd1 _05783_ sky130_fd_sc_hd__a211oi_1
Xhold982 final_design.cpu.reg_window\[405\] vssd1 vssd1 vccd1 vccd1 net2324 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12878__CLK clknet_leaf_17_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold993 final_design.cpu.reg_window\[259\] vssd1 vssd1 vccd1 vccd1 net2335 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout771_X net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12171__A1 net244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10011_ net460 _03641_ _04237_ _04929_ vssd1 vssd1 vccd1 vccd1 _04930_ sky130_fd_sc_hd__a31o_1
XANTENNA__08375__B1 _02211_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11746__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_34_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_26_Right_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_34_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11962_ _06164_ net280 net405 net1726 vssd1 vssd1 vccd1 vccd1 _00695_ sky130_fd_sc_hd__a22o_1
XANTENNA__08222__S0 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12474__A2 net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13701_ clknet_leaf_49_clk _00932_ net1182 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[689\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_1394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10913_ net50 _05642_ vssd1 vssd1 vccd1 vccd1 _05643_ sky130_fd_sc_hd__and2_1
XANTENNA__11682__B1 net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11893_ net221 net2199 net272 vssd1 vssd1 vccd1 vccd1 _00635_ sky130_fd_sc_hd__mux2_1
XANTENNA__11481__S net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13632_ clknet_leaf_11_clk _00863_ net1090 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[620\]
+ sky130_fd_sc_hd__dfrtp_1
X_10844_ net962 _05576_ vssd1 vssd1 vccd1 vccd1 _05577_ sky130_fd_sc_hd__nand2_1
XFILLER_0_71_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_15_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12874__Q final_design.data_from_mem\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13503__CLK clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09722__S0 net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13563_ clknet_leaf_0_clk _00794_ net1063 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[551\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10775_ net75 net1044 vssd1 vssd1 vccd1 vccd1 _05511_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_35_Right_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12514_ _06176_ net348 net329 net1737 vssd1 vssd1 vccd1 vccd1 _01219_ sky130_fd_sc_hd__a22o_1
X_13494_ clknet_leaf_59_clk _00725_ net1138 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[482\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07653__A2 _02602_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12445_ net2436 net210 net336 vssd1 vssd1 vccd1 vccd1 _01152_ sky130_fd_sc_hd__mux2_1
XANTENNA__13653__CLK clknet_leaf_58_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08803__B _01722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1917 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12376_ net1768 net213 net268 vssd1 vssd1 vccd1 vccd1 _01087_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14115_ clknet_leaf_14_clk _01312_ net1110 vssd1 vssd1 vccd1 vccd1 final_design.reqhand.data_from_UART\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11327_ net737 _03878_ _06019_ vssd1 vssd1 vccd1 vccd1 _06020_ sky130_fd_sc_hd__a21oi_1
X_14046_ clknet_leaf_16_clk _00007_ net1092 vssd1 vssd1 vccd1 vccd1 final_design.uart.BAUD_counter\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14009__CLK clknet_leaf_56_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11258_ net434 net578 _05959_ net316 net1789 vssd1 vssd1 vccd1 vccd1 _00288_ sky130_fd_sc_hd__a32o_1
XFILLER_0_5_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_44_Right_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10209_ final_design.uart.BAUD_counter\[3\] _05093_ vssd1 vssd1 vccd1 vccd1 _05094_
+ sky130_fd_sc_hd__and2_1
X_11189_ net430 net569 _05898_ net315 net1667 vssd1 vssd1 vccd1 vccd1 _00280_ sky130_fd_sc_hd__a32o_1
XANTENNA__13033__CLK clknet_leaf_40_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14159__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12465__A2 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1833 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07420_ final_design.cpu.reg_window\[1\] final_design.cpu.reg_window\[33\] net916
+ vssd1 vssd1 vccd1 vccd1 _02371_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_1877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13183__CLK clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_53_Right_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08516__S1 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07351_ final_design.cpu.reg_window\[259\] final_design.cpu.reg_window\[291\] net915
+ vssd1 vssd1 vccd1 vccd1 _02302_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09094__A1 net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07282_ final_design.cpu.reg_window\[582\] final_design.cpu.reg_window\[614\] net902
+ vssd1 vssd1 vccd1 vccd1 _02233_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09021_ _02067_ _02447_ net623 vssd1 vssd1 vccd1 vccd1 _03953_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_54_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11728__A1 net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold201 final_design.cpu.reg_window\[969\] vssd1 vssd1 vccd1 vccd1 net1543 sky130_fd_sc_hd__dlygate4sd3_1
Xhold212 final_design.cpu.reg_window\[462\] vssd1 vssd1 vccd1 vccd1 net1554 sky130_fd_sc_hd__dlygate4sd3_1
Xhold223 final_design.reqhand.instruction\[1\] vssd1 vssd1 vccd1 vccd1 net1565 sky130_fd_sc_hd__dlygate4sd3_1
Xhold234 final_design.cpu.reg_window\[50\] vssd1 vssd1 vccd1 vccd1 net1576 sky130_fd_sc_hd__dlygate4sd3_1
Xhold245 final_design.cpu.reg_window\[474\] vssd1 vssd1 vccd1 vccd1 net1587 sky130_fd_sc_hd__dlygate4sd3_1
Xhold256 final_design.cpu.reg_window\[684\] vssd1 vssd1 vccd1 vccd1 net1598 sky130_fd_sc_hd__dlygate4sd3_1
Xhold267 final_design.cpu.reg_window\[758\] vssd1 vssd1 vccd1 vccd1 net1609 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_62_Right_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold278 final_design.cpu.reg_window\[478\] vssd1 vssd1 vccd1 vccd1 net1620 sky130_fd_sc_hd__dlygate4sd3_1
X_09923_ _04109_ _04398_ _04838_ _04222_ _04833_ vssd1 vssd1 vccd1 vccd1 _04842_ sky130_fd_sc_hd__o221a_1
Xfanout703 net706 vssd1 vssd1 vccd1 vccd1 net703 sky130_fd_sc_hd__clkbuf_4
Xhold289 final_design.cpu.reg_window\[686\] vssd1 vssd1 vccd1 vccd1 net1631 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06801__X _01752_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout714 net715 vssd1 vssd1 vccd1 vccd1 net714 sky130_fd_sc_hd__buf_4
XANTENNA_fanout397_A _06261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout725 net726 vssd1 vssd1 vccd1 vccd1 net725 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_0_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout736 _01490_ vssd1 vssd1 vccd1 vccd1 net736 sky130_fd_sc_hd__clkbuf_4
X_09854_ net480 _04406_ _04691_ net492 vssd1 vssd1 vccd1 vccd1 _04773_ sky130_fd_sc_hd__a211o_1
Xfanout747 _01438_ vssd1 vssd1 vccd1 vccd1 net747 sky130_fd_sc_hd__clkbuf_8
XANTENNA__09544__B _04094_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout758 net759 vssd1 vssd1 vccd1 vccd1 net758 sky130_fd_sc_hd__clkbuf_2
Xfanout769 net771 vssd1 vssd1 vccd1 vccd1 net769 sky130_fd_sc_hd__buf_4
XANTENNA_fanout1104_A net1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09036__S net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08805_ final_design.CPU_instr_adr\[23\] _01722_ vssd1 vssd1 vccd1 vccd1 _03756_
+ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_52_1981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09785_ net96 _04179_ vssd1 vssd1 vccd1 vccd1 _04704_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_52_1992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06997_ final_design.cpu.reg_window\[79\] final_design.cpu.reg_window\[111\] net888
+ vssd1 vssd1 vccd1 vccd1 _01948_ sky130_fd_sc_hd__mux2_1
X_08736_ _01365_ _02064_ vssd1 vssd1 vccd1 vccd1 _03687_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09857__B1 net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10467__A1 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13526__CLK clknet_leaf_61_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10467__B2 net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11664__B1 net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout731_A net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08667_ _01998_ _02061_ vssd1 vssd1 vccd1 vccd1 _03618_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout352_X net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_71_Right_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11154__X _05868_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout829_A _01818_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07618_ _02563_ _02568_ net719 vssd1 vssd1 vccd1 vccd1 _02569_ sky130_fd_sc_hd__mux2_1
XANTENNA__12208__A2 _06136_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08598_ net875 _03542_ _03548_ _03535_ _03536_ vssd1 vssd1 vccd1 vccd1 _03549_ sky130_fd_sc_hd__a32oi_4
XTAP_TAPCELL_ROW_27_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07549_ _02496_ _02497_ _02498_ _02499_ net774 net783 vssd1 vssd1 vccd1 vccd1 _02500_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_46_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13676__CLK clknet_leaf_45_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1887 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_23_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12129__C net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10560_ _05283_ _05303_ vssd1 vssd1 vccd1 vccd1 _05307_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_42_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14202__1260 vssd1 vssd1 vccd1 vccd1 _14202__1260/HI net1260 sky130_fd_sc_hd__conb_1
X_09219_ _03132_ _03162_ vssd1 vssd1 vccd1 vccd1 _04138_ sky130_fd_sc_hd__and2b_1
X_10491_ net960 _05237_ _05238_ _04042_ vssd1 vssd1 vccd1 vccd1 _05241_ sky130_fd_sc_hd__a22o_1
XANTENNA__09388__A2 _02325_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12230_ net230 net2505 net372 vssd1 vssd1 vccd1 vccd1 _00947_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_10_clk_A clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06438__1 clknet_leaf_26_clk vssd1 vssd1 vccd1 vccd1 net1311 sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_80_Right_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11195__A2 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12161_ net176 net2500 net386 vssd1 vssd1 vccd1 vccd1 _00882_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11112_ _05831_ _05830_ final_design.uart.bits_received\[0\] vssd1 vssd1 vccd1 vccd1
+ _00205_ sky130_fd_sc_hd__mux2_1
XANTENNA__09735__A net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12092_ net578 _06082_ net510 net394 net1837 vssd1 vssd1 vccd1 vccd1 _00817_ sky130_fd_sc_hd__a32o_1
Xhold790 final_design.cpu.reg_window\[39\] vssd1 vssd1 vccd1 vccd1 net2132 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11476__S net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13056__CLK clknet_leaf_11_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_25_clk_A clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11043_ _05765_ _05766_ vssd1 vssd1 vccd1 vccd1 _05767_ sky130_fd_sc_hd__nor2_1
XFILLER_0_60_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12869__Q final_design.data_from_mem\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12994_ net1325 _00225_ net1194 vssd1 vssd1 vccd1 vccd1 final_design.CPU_instr_adr\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_8_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_1765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11945_ _06146_ net289 net411 net2433 vssd1 vssd1 vccd1 vccd1 _00680_ sky130_fd_sc_hd__a22o_1
XFILLER_0_52_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12100__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11876_ net2527 net519 _06245_ net434 vssd1 vssd1 vccd1 vccd1 _00620_ sky130_fd_sc_hd__a22o_1
XFILLER_0_54_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13615_ clknet_leaf_44_clk _00846_ net1208 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[603\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11407__B1 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10827_ net45 _05558_ vssd1 vssd1 vccd1 vccd1 _05561_ sky130_fd_sc_hd__nor2_1
XANTENNA__12080__B1 net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13546_ clknet_leaf_60_clk _00777_ net1141 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[534\]
+ sky130_fd_sc_hd__dfrtp_1
X_10758_ net962 _05494_ vssd1 vssd1 vccd1 vccd1 _05495_ sky130_fd_sc_hd__nand2_1
XANTENNA__13597__RESET_B net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13477_ clknet_leaf_49_clk _00708_ net1182 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[465\]
+ sky130_fd_sc_hd__dfrtp_1
X_10689_ _05427_ _05428_ vssd1 vssd1 vccd1 vccd1 _05429_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12428_ _06115_ net353 net340 net1930 vssd1 vssd1 vccd1 vccd1 _01137_ sky130_fd_sc_hd__a22o_1
XANTENNA__12383__A1 _06003_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_995 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12623__X _06298_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12359_ net2535 net362 net357 _06068_ vssd1 vssd1 vccd1 vccd1 _01071_ sky130_fd_sc_hd__a22o_1
XFILLER_0_77_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07717__X _02668_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14029_ clknet_leaf_48_clk _01260_ net1200 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[1017\]
+ sky130_fd_sc_hd__dfrtp_1
X_06920_ final_design.cpu.reg_window\[978\] final_design.cpu.reg_window\[1010\] net925
+ vssd1 vssd1 vccd1 vccd1 _01871_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_1501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13549__CLK clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11894__A0 net219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06851_ net761 _01801_ vssd1 vssd1 vccd1 vccd1 _01802_ sky130_fd_sc_hd__nor2_1
XANTENNA__09551__A2 _04046_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06996__S0 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09570_ _01626_ _01657_ net552 _01717_ net453 net462 vssd1 vssd1 vccd1 vccd1 _04489_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_56_1810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06782_ final_design.cpu.reg_window\[22\] final_design.cpu.reg_window\[54\] net918
+ vssd1 vssd1 vccd1 vccd1 _01733_ sky130_fd_sc_hd__mux2_1
X_08521_ final_design.cpu.reg_window\[962\] final_design.cpu.reg_window\[994\] net833
+ vssd1 vssd1 vccd1 vccd1 _03472_ sky130_fd_sc_hd__mux2_1
XANTENNA__10449__B2 net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11646__B1 net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08708__B _01570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13699__CLK clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08452_ net709 _03396_ net722 vssd1 vssd1 vccd1 vccd1 _03403_ sky130_fd_sc_hd__o21a_1
XFILLER_0_9_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07403_ _02350_ _02351_ _02352_ _02353_ net769 net782 vssd1 vssd1 vccd1 vccd1 _02354_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_4_1527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11134__B net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08383_ final_design.cpu.reg_window\[70\] final_design.cpu.reg_window\[102\] net823
+ vssd1 vssd1 vccd1 vccd1 _03334_ sky130_fd_sc_hd__mux2_1
X_07334_ final_design.cpu.reg_window\[964\] final_design.cpu.reg_window\[996\] net905
+ vssd1 vssd1 vccd1 vccd1 _02285_ sky130_fd_sc_hd__mux2_1
XANTENNA__12071__B1 net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07173__S0 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07265_ final_design.cpu.reg_window\[326\] final_design.cpu.reg_window\[358\] net912
+ vssd1 vssd1 vccd1 vccd1 _02216_ sky130_fd_sc_hd__mux2_1
XANTENNA__11788__C net207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout312_A net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1054_A net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09004_ _03683_ _03737_ vssd1 vssd1 vccd1 vccd1 _03938_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_28_1901 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07196_ _02143_ _02144_ _02145_ _02146_ net764 net785 vssd1 vssd1 vccd1 vccd1 _02147_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__11177__A2 net251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12374__A1 net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13079__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08042__A2 _02991_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07774__S net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout500 net501 vssd1 vssd1 vccd1 vccd1 net500 sky130_fd_sc_hd__buf_4
XANTENNA__12126__A1 net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout681_A net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout511 net515 vssd1 vssd1 vccd1 vccd1 net511 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout779_A _01422_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout522 net524 vssd1 vssd1 vccd1 vccd1 net522 sky130_fd_sc_hd__buf_4
X_09906_ _04072_ _04824_ _04810_ vssd1 vssd1 vccd1 vccd1 _04825_ sky130_fd_sc_hd__o21ai_2
Xfanout533 _02211_ vssd1 vssd1 vccd1 vccd1 net533 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_50_1907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout544 _01937_ vssd1 vssd1 vccd1 vccd1 net544 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_50_1918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout555 _05869_ vssd1 vssd1 vccd1 vccd1 net555 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_50_1929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout566 net567 vssd1 vssd1 vccd1 vccd1 net566 sky130_fd_sc_hd__buf_2
Xfanout577 net587 vssd1 vssd1 vccd1 vccd1 net577 sky130_fd_sc_hd__clkbuf_4
X_09837_ net481 _04755_ _04341_ vssd1 vssd1 vccd1 vccd1 _04756_ sky130_fd_sc_hd__a21o_1
XANTENNA__09542__A2 _04366_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout588 net591 vssd1 vssd1 vccd1 vccd1 net588 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout946_A net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout567_X net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout599 net601 vssd1 vssd1 vccd1 vccd1 net599 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12916__CLK clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09768_ net320 _04683_ _04684_ net319 _04686_ vssd1 vssd1 vccd1 vccd1 _04687_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_1_240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08719_ _03669_ vssd1 vssd1 vccd1 vccd1 _03670_ sky130_fd_sc_hd__inv_2
XFILLER_0_35_1905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_1_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09699_ net544 net542 net541 net540 net454 net464 vssd1 vssd1 vccd1 vccd1 _04618_
+ sky130_fd_sc_hd__mux4_2
XTAP_TAPCELL_ROW_29_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11730_ net436 net584 _06223_ net296 net2156 vssd1 vssd1 vccd1 vccd1 _00496_ sky130_fd_sc_hd__a32o_1
XFILLER_0_7_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07014__S net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11661_ net182 net632 vssd1 vssd1 vccd1 vccd1 _06188_ sky130_fd_sc_hd__and2_1
X_13400_ clknet_leaf_63_clk _00631_ net1121 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[388\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_64_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10612_ _05354_ _05355_ vssd1 vssd1 vccd1 vccd1 _05356_ sky130_fd_sc_hd__nand2_1
XANTENNA__12062__A0 net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11592_ net184 net637 vssd1 vssd1 vccd1 vccd1 _06152_ sky130_fd_sc_hd__and2_1
XFILLER_0_25_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13331_ clknet_leaf_40_clk _00562_ net1211 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[319\]
+ sky130_fd_sc_hd__dfrtp_1
X_10543_ net94 final_design.VGA_adr\[2\] _05289_ vssd1 vssd1 vccd1 vccd1 _05290_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_49_1157 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input75_A memory_size[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13262_ clknet_leaf_45_clk _00493_ net1213 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[250\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10474_ net801 _05224_ vssd1 vssd1 vccd1 vccd1 _05225_ sky130_fd_sc_hd__or2_1
X_12213_ net573 _06141_ net508 net379 net1570 vssd1 vssd1 vccd1 vccd1 _00931_ sky130_fd_sc_hd__a32o_1
X_13193_ clknet_leaf_36_clk _00424_ net1228 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[181\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10376__B1 net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12144_ net208 net2420 net384 vssd1 vssd1 vccd1 vccd1 _00865_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12117__A1 net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12075_ net577 _05959_ net511 net394 net1610 vssd1 vssd1 vccd1 vccd1 _00800_ sky130_fd_sc_hd__a32o_1
XANTENNA__10404__A _03450_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_2590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input30_X net30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11026_ _05729_ _05733_ _05749_ vssd1 vssd1 vccd1 vccd1 _05751_ sky130_fd_sc_hd__o21ai_1
XANTENNA__06978__S0 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13841__CLK clknet_leaf_34_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11628__B1 net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12977_ clknet_leaf_21_clk _00002_ net1160 vssd1 vssd1 vccd1 vccd1 final_design.reqhand.current_client\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_11928_ _06130_ net283 net409 net2113 vssd1 vssd1 vccd1 vccd1 _00664_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_64_2383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13991__CLK clknet_leaf_63_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_2394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_25_Left_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11859_ net2431 net517 _06241_ net427 vssd1 vssd1 vccd1 vccd1 _00607_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_60_2247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_2258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_18 _06228_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_2269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06616__X _01567_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_29 _06257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07155__S0 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13529_ clknet_leaf_54_clk _00760_ net1177 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[517\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13221__CLK clknet_leaf_49_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07050_ _01996_ _02000_ vssd1 vssd1 vccd1 vccd1 _02001_ sky130_fd_sc_hd__nand2_1
XFILLER_0_42_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12356__B2 _06046_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput103 net103 vssd1 vssd1 vccd1 vccd1 ADR_O[11] sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_58_2176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput114 net114 vssd1 vssd1 vccd1 vccd1 ADR_O[21] sky130_fd_sc_hd__clkbuf_4
XANTENNA__09221__A1 _02126_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_2187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput125 net125 vssd1 vssd1 vccd1 vccd1 ADR_O[31] sky130_fd_sc_hd__clkbuf_4
XANTENNA__10367__B1 net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_2198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput136 net136 vssd1 vssd1 vccd1 vccd1 DAT_O[11] sky130_fd_sc_hd__clkbuf_4
Xoutput147 net147 vssd1 vssd1 vccd1 vccd1 DAT_O[21] sky130_fd_sc_hd__buf_2
XFILLER_0_10_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput158 net158 vssd1 vssd1 vccd1 vccd1 DAT_O[31] sky130_fd_sc_hd__clkbuf_4
Xoutput169 net169 vssd1 vssd1 vccd1 vccd1 SEL_O[3] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_34_Left_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12939__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07952_ _02838_ _02901_ vssd1 vssd1 vccd1 vccd1 _02903_ sky130_fd_sc_hd__nand2_1
XANTENNA__07619__A1_N net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09662__X _04581_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06903_ _01853_ vssd1 vssd1 vccd1 vccd1 _01854_ sky130_fd_sc_hd__inv_2
XANTENNA__11867__B1 net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07883_ net549 _02832_ vssd1 vssd1 vccd1 vccd1 _02834_ sky130_fd_sc_hd__nand2b_2
X_09622_ _02868_ net446 net442 _02866_ _04535_ vssd1 vssd1 vccd1 vccd1 _04541_ sky130_fd_sc_hd__o221ai_2
X_06834_ net886 _01777_ _01783_ _01765_ _01771_ vssd1 vssd1 vccd1 vccd1 _01785_ sky130_fd_sc_hd__a32o_1
XFILLER_0_37_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11882__A3 net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07623__A _01536_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09553_ _02935_ _04471_ vssd1 vssd1 vccd1 vccd1 _04472_ sky130_fd_sc_hd__xnor2_1
X_06765_ net763 _01715_ vssd1 vssd1 vccd1 vccd1 _01716_ sky130_fd_sc_hd__or2_1
XFILLER_0_77_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout262_A net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08504_ _02325_ net490 vssd1 vssd1 vccd1 vccd1 _03455_ sky130_fd_sc_hd__nor2_1
X_09484_ _04401_ _04402_ net477 vssd1 vssd1 vccd1 vccd1 _04403_ sky130_fd_sc_hd__mux2_1
XANTENNA__12292__B1 net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06696_ final_design.cpu.reg_window\[985\] final_design.cpu.reg_window\[1017\] net933
+ vssd1 vssd1 vccd1 vccd1 _01647_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_43_Left_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09693__D1 _04045_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08435_ net597 _03384_ _03360_ vssd1 vssd1 vccd1 vccd1 _03386_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_59_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1171_A net1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout527_A _02502_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07769__S net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08366_ final_design.cpu.reg_window\[583\] final_design.cpu.reg_window\[615\] net806
+ vssd1 vssd1 vccd1 vccd1 _03317_ sky130_fd_sc_hd__mux2_1
XANTENNA__11799__B _05869_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11398__A2 net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12972__Q final_design.CPU_instr_adr\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12595__B2 final_design.data_from_mem\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07317_ net531 _02267_ vssd1 vssd1 vccd1 vccd1 _02268_ sky130_fd_sc_hd__nor2_1
XFILLER_0_11_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08297_ final_design.cpu.reg_window\[649\] final_design.cpu.reg_window\[681\] net807
+ vssd1 vssd1 vccd1 vccd1 _03248_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout315_X net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09460__A1 net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07697__S1 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09460__B2 _04117_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1057_X net1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10070__A2 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07248_ net749 _02198_ net745 vssd1 vssd1 vccd1 vccd1 _02199_ sky130_fd_sc_hd__o21a_1
XANTENNA__13714__CLK clknet_leaf_38_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout896_A net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09748__C1 _04097_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10358__B1 net1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_52_Left_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07449__S1 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12263__X _06274_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07179_ _02127_ _02128_ vssd1 vssd1 vccd1 vccd1 _02130_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_24_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10190_ _05066_ _05079_ vssd1 vssd1 vccd1 vccd1 _05080_ sky130_fd_sc_hd__nand2_4
XANTENNA_fanout684_X net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_1098 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13864__CLK clknet_leaf_41_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout330 net331 vssd1 vssd1 vccd1 vccd1 net330 sky130_fd_sc_hd__buf_4
Xfanout341 _06279_ vssd1 vssd1 vccd1 vccd1 net341 sky130_fd_sc_hd__buf_4
Xfanout352 net359 vssd1 vssd1 vccd1 vccd1 net352 sky130_fd_sc_hd__buf_2
XANTENNA__09515__A2 net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout851_X net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout363 _06276_ vssd1 vssd1 vccd1 vccd1 net363 sky130_fd_sc_hd__clkbuf_8
Xfanout374 net375 vssd1 vssd1 vccd1 vccd1 net374 sky130_fd_sc_hd__buf_4
Xfanout385 _06266_ vssd1 vssd1 vccd1 vccd1 net385 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11754__S net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout396 net397 vssd1 vssd1 vccd1 vccd1 net396 sky130_fd_sc_hd__clkbuf_8
X_12900_ clknet_leaf_25_clk _00138_ net1154 vssd1 vssd1 vccd1 vccd1 net166 sky130_fd_sc_hd__dfrtp_2
X_13880_ clknet_leaf_63_clk _01111_ net1076 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[868\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12831_ net1377 vssd1 vssd1 vccd1 vccd1 _00272_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_61_Left_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12762_ _06397_ vssd1 vssd1 vccd1 vccd1 _06398_ sky130_fd_sc_hd__inv_2
XANTENNA__12283__B1 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11713_ net590 net196 net628 vssd1 vssd1 vccd1 vccd1 _06215_ sky130_fd_sc_hd__and3_1
X_12693_ final_design.VGA_data_control.v_count\[6\] _01403_ vssd1 vssd1 vccd1 vccd1
+ _06334_ sky130_fd_sc_hd__nor2_1
XANTENNA__13244__CLK clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07679__S net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11644_ net428 net567 _06179_ net299 net2121 vssd1 vssd1 vccd1 vccd1 _00454_ sky130_fd_sc_hd__a32o_1
XANTENNA__12882__Q final_design.data_from_mem\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12586__B2 final_design.data_from_mem\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput16 DAT_I[22] vssd1 vssd1 vccd1 vccd1 net16 sky130_fd_sc_hd__clkbuf_1
X_11575_ net573 net424 _06143_ net305 net1698 vssd1 vssd1 vccd1 vccd1 _00421_ sky130_fd_sc_hd__a32o_1
Xinput27 DAT_I[3] vssd1 vssd1 vccd1 vccd1 net27 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_80_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput38 mem_adr_start[11] vssd1 vssd1 vccd1 vccd1 net38 sky130_fd_sc_hd__buf_1
X_13314_ clknet_leaf_4_clk _00545_ net1083 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[302\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput49 mem_adr_start[21] vssd1 vssd1 vccd1 vccd1 net49 sky130_fd_sc_hd__buf_1
X_10526_ _05270_ _05271_ _05272_ vssd1 vssd1 vccd1 vccd1 _05274_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_1777 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13394__CLK clknet_leaf_39_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_70_Left_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12338__B2 _05911_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13245_ clknet_leaf_2_clk _00476_ net1065 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[233\]
+ sky130_fd_sc_hd__dfrtp_1
X_10457_ net2353 net1033 _05212_ net248 vssd1 vssd1 vccd1 vccd1 _00169_ sky130_fd_sc_hd__a22o_1
XANTENNA__08370__Y _03321_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_72_2652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13176_ clknet_leaf_65_clk _00407_ net1073 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[164\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_72_2663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10388_ _03648_ _04991_ _04987_ vssd1 vssd1 vccd1 vccd1 _05175_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_72_2674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11561__A2 net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12127_ _06094_ net506 vssd1 vssd1 vccd1 vccd1 _06266_ sky130_fd_sc_hd__nand2_2
XANTENNA__11849__B1 net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12058_ net2348 net176 net398 vssd1 vssd1 vccd1 vccd1 _00786_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11009_ _05733_ _05734_ net1433 net1033 vssd1 vssd1 vccd1 vccd1 _00199_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__07612__S1 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_2445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_66_2467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_2309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12274__B1 net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06550_ final_design.reqhand.instruction\[31\] final_design.data_from_mem\[31\] net973
+ vssd1 vssd1 vccd1 vccd1 _01501_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10824__A1 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10824__B2 net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06481_ final_design.cpu.reg_window\[30\] final_design.cpu.reg_window\[62\] net936
+ vssd1 vssd1 vccd1 vccd1 _01432_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08220_ final_design.cpu.reg_window\[459\] final_design.cpu.reg_window\[491\] net835
+ vssd1 vssd1 vccd1 vccd1 _03171_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13737__CLK clknet_leaf_36_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08151_ _03099_ _03100_ vssd1 vssd1 vccd1 vccd1 _03102_ sky130_fd_sc_hd__or2_1
XANTENNA__08245__A2 _03192_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07102_ final_design.cpu.reg_window\[652\] final_design.cpu.reg_window\[684\] net893
+ vssd1 vssd1 vccd1 vccd1 _02053_ sky130_fd_sc_hd__mux2_1
X_08082_ _02965_ _02996_ _03028_ _03032_ vssd1 vssd1 vccd1 vccd1 _03033_ sky130_fd_sc_hd__o31ai_2
XFILLER_0_71_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08650__C1 _01597_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11839__S net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07033_ final_design.cpu.reg_window\[782\] final_design.cpu.reg_window\[814\] net906
+ vssd1 vssd1 vccd1 vccd1 _01984_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13887__CLK clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_1238 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08984_ final_design.CPU_instr_adr\[17\] net1016 _03916_ _03920_ vssd1 vssd1 vccd1
+ vccd1 _00228_ sky130_fd_sc_hd__a22o_1
XANTENNA__13117__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07935_ _02882_ _02883_ _02884_ _02885_ net680 net700 vssd1 vssd1 vccd1 vccd1 _02886_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_23_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07866_ net720 _02816_ vssd1 vssd1 vccd1 vccd1 _02817_ sky130_fd_sc_hd__nor2_1
XFILLER_0_58_1746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09044__S net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09605_ _04446_ _04523_ _04228_ vssd1 vssd1 vccd1 vccd1 _04524_ sky130_fd_sc_hd__o21ai_1
X_06817_ final_design.cpu.reg_window\[469\] final_design.cpu.reg_window\[501\] net939
+ vssd1 vssd1 vccd1 vccd1 _01768_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout644_A net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07797_ final_design.cpu.reg_window\[153\] final_design.cpu.reg_window\[185\] net855
+ vssd1 vssd1 vccd1 vccd1 _02748_ sky130_fd_sc_hd__mux2_1
XANTENNA__13629__RESET_B net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13267__CLK clknet_leaf_40_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout265_X net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09536_ _04454_ vssd1 vssd1 vccd1 vccd1 _04455_ sky130_fd_sc_hd__inv_2
XANTENNA__12265__B1 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06748_ final_design.cpu.reg_window\[23\] final_design.cpu.reg_window\[55\] net929
+ vssd1 vssd1 vccd1 vccd1 _01699_ sky130_fd_sc_hd__mux2_1
XANTENNA__08469__C1 _02294_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09467_ net85 _04192_ vssd1 vssd1 vccd1 vccd1 _04386_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_1290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14186__A net169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout432_X net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout811_A net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06679_ net741 _01497_ net665 _01629_ vssd1 vssd1 vccd1 vccd1 _01630_ sky130_fd_sc_hd__a211o_4
XANTENNA__12280__A3 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout909_A net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11162__X _05875_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12017__B1 net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08418_ final_design.cpu.reg_window\[133\] final_design.cpu.reg_window\[165\] net841
+ vssd1 vssd1 vccd1 vccd1 _03369_ sky130_fd_sc_hd__mux2_1
XANTENNA__11603__A net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09398_ net479 _04302_ _04316_ _04109_ vssd1 vssd1 vccd1 vccd1 _04317_ sky130_fd_sc_hd__a211o_1
XANTENNA__12775__6_A clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10028__C1 net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12418__B net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08349_ final_design.cpu.reg_window\[455\] final_design.cpu.reg_window\[487\] net811
+ vssd1 vssd1 vccd1 vccd1 _03300_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11240__A1 final_design.data_from_mem\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11360_ final_design.data_from_mem\[26\] net235 net233 vssd1 vssd1 vccd1 vccd1 _06049_
+ sky130_fd_sc_hd__a21o_2
XFILLER_0_69_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout899_X net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10311_ _04999_ _05040_ _05164_ vssd1 vssd1 vccd1 vccd1 final_design.pixel_data sky130_fd_sc_hd__and3_2
XANTENNA__11749__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11791__A2 net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10653__S net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11291_ _04473_ net658 _05843_ _05988_ vssd1 vssd1 vccd1 vccd1 _05989_ sky130_fd_sc_hd__a211oi_4
X_13030_ clknet_leaf_50_clk _00261_ net1168 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_10242_ final_design.uart.BAUD_counter\[15\] _05113_ net798 vssd1 vssd1 vccd1 vccd1
+ _05115_ sky130_fd_sc_hd__o21ai_1
XPHY_EDGE_ROW_5_Left_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08123__S net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08095__S1 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11543__A2 net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07747__B2 net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10173_ _05017_ _05061_ vssd1 vssd1 vccd1 vccd1 final_design.vga.h_next_state\[1\]
+ sky130_fd_sc_hd__nor2_1
Xfanout1103 net1105 vssd1 vssd1 vccd1 vccd1 net1103 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_28_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1114 net1115 vssd1 vssd1 vccd1 vccd1 net1114 sky130_fd_sc_hd__clkbuf_4
Xfanout1125 net1127 vssd1 vssd1 vccd1 vccd1 net1125 sky130_fd_sc_hd__clkbuf_4
XANTENNA__14042__CLK clknet_leaf_15_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1136 net1137 vssd1 vssd1 vccd1 vccd1 net1136 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09743__A net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input38_A mem_adr_start[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1147 net1148 vssd1 vssd1 vccd1 vccd1 net1147 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_41_1783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1158 net1159 vssd1 vssd1 vccd1 vccd1 net1158 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11484__S net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1169 net1176 vssd1 vssd1 vccd1 vccd1 net1169 sky130_fd_sc_hd__clkbuf_2
Xfanout182 _06067_ vssd1 vssd1 vccd1 vccd1 net182 sky130_fd_sc_hd__clkbuf_2
X_13932_ clknet_leaf_46_clk _01163_ net1217 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[920\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout193 _06031_ vssd1 vssd1 vccd1 vccd1 net193 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_76_1857 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12877__Q final_design.data_from_mem\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13863_ clknet_leaf_59_clk _01094_ net1126 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[851\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12814_ net1415 vssd1 vssd1 vccd1 vccd1 _00255_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__12256__B1 net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13794_ clknet_leaf_4_clk _01025_ net1084 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[782\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_80_2921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12745_ _06359_ _06379_ vssd1 vssd1 vccd1 vccd1 _06384_ sky130_fd_sc_hd__nand2_1
XANTENNA__12271__A3 net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06486__A1 final_design.data_from_mem\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12008__B1 net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12676_ _06325_ net1495 net978 vssd1 vssd1 vccd1 vccd1 _01340_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11627_ net215 net631 vssd1 vssd1 vccd1 vccd1 _06171_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_13_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_2861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11558_ net216 net634 vssd1 vssd1 vccd1 vccd1 _06135_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_78_2872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12934__RESET_B net1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_2883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08273__A1_N net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_2725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10585__A3 net247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11782__A2 net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold608 final_design.cpu.reg_window\[270\] vssd1 vssd1 vccd1 vccd1 net1950 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_55_2102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10509_ _05256_ _05257_ vssd1 vssd1 vccd1 vccd1 _05258_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_74_2736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold619 final_design.cpu.reg_window\[567\] vssd1 vssd1 vccd1 vccd1 net1961 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11489_ net184 net2218 net308 vssd1 vssd1 vccd1 vccd1 _00366_ sky130_fd_sc_hd__mux2_1
X_13228_ clknet_leaf_46_clk _00459_ net1214 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[216\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13159_ clknet_leaf_62_clk _00390_ net1123 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[147\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_68_2518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07720_ net615 _02668_ _02669_ _01596_ vssd1 vssd1 vccd1 vccd1 _02671_ sky130_fd_sc_hd__a211oi_2
XTAP_TAPCELL_ROW_68_2529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11298__A1 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12495__B1 net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1889 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07651_ net878 _02583_ _02589_ _02595_ _02601_ vssd1 vssd1 vccd1 vccd1 _02602_ sky130_fd_sc_hd__o32a_2
X_06602_ net754 _01552_ net747 vssd1 vssd1 vccd1 vccd1 _01553_ sky130_fd_sc_hd__o21a_1
X_07582_ net720 _02532_ vssd1 vssd1 vccd1 vccd1 _02533_ sky130_fd_sc_hd__nor2_1
XFILLER_0_34_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09321_ net460 _04237_ _04238_ _04239_ vssd1 vssd1 vccd1 vccd1 _04240_ sky130_fd_sc_hd__a31o_1
XFILLER_0_76_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06533_ _01474_ _01481_ _01482_ vssd1 vssd1 vccd1 vccd1 _01484_ sky130_fd_sc_hd__nor3_2
XFILLER_0_34_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09663__A1 net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12262__A3 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08716__B _01660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09252_ _04167_ _04170_ _02609_ vssd1 vssd1 vccd1 vccd1 _04171_ sky130_fd_sc_hd__a21o_1
X_06464_ net1041 net993 net990 vssd1 vssd1 vccd1 vccd1 _01415_ sky130_fd_sc_hd__and3_2
XFILLER_0_44_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08203_ final_design.cpu.reg_window\[718\] final_design.cpu.reg_window\[750\] net816
+ vssd1 vssd1 vccd1 vccd1 _03154_ sky130_fd_sc_hd__mux2_1
X_09183_ net614 net525 _03523_ _01567_ vssd1 vssd1 vccd1 vccd1 _04102_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout225_A _05897_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08134_ final_design.cpu.reg_window\[589\] final_design.cpu.reg_window\[621\] net855
+ vssd1 vssd1 vccd1 vccd1 _03085_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1436 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11773__A2 net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10473__S net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08065_ final_design.cpu.reg_window\[722\] final_design.cpu.reg_window\[754\] net845
+ vssd1 vssd1 vccd1 vccd1 _03016_ sky130_fd_sc_hd__mux2_1
XANTENNA__11796__C net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07348__A _02294_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07016_ net927 _01852_ _01821_ vssd1 vssd1 vccd1 vccd1 _01967_ sky130_fd_sc_hd__a21bo_1
XANTENNA__14065__CLK clknet_leaf_15_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11525__A2 _06120_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout594_A _03627_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08967_ _01884_ _02457_ vssd1 vssd1 vccd1 vccd1 _03905_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout761_A net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout382_X net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout859_A net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07918_ _01755_ net613 vssd1 vssd1 vccd1 vccd1 _02869_ sky130_fd_sc_hd__or2_1
XANTENNA__12486__B1 net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08898_ _03799_ _03843_ vssd1 vssd1 vccd1 vccd1 _03844_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_32_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_4_clk_X clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07849_ net606 _02797_ _02773_ net550 vssd1 vssd1 vccd1 vccd1 _02800_ sky130_fd_sc_hd__o211a_1
XANTENNA__13902__CLK clknet_leaf_43_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout647_X net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10860_ _05591_ vssd1 vssd1 vccd1 vccd1 _05592_ sky130_fd_sc_hd__inv_2
XANTENNA__12238__B1 net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09519_ net492 _04437_ vssd1 vssd1 vccd1 vccd1 _04438_ sky130_fd_sc_hd__and2_1
X_10791_ _05525_ _05526_ net1425 net1032 vssd1 vssd1 vccd1 vccd1 _00189_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_78_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12253__A3 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12530_ net673 _06193_ _06260_ vssd1 vssd1 vccd1 vccd1 _06285_ sky130_fd_sc_hd__or3_4
XANTENNA__06468__A1 final_design.data_from_mem\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12461_ net2215 net181 net336 vssd1 vssd1 vccd1 vccd1 _01168_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_23_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14200_ net1258 vssd1 vssd1 vccd1 vccd1 gpio_oeb[12] sky130_fd_sc_hd__buf_2
XFILLER_0_1_1861 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11412_ net1678 net242 net311 vssd1 vssd1 vccd1 vccd1 _00309_ sky130_fd_sc_hd__mux2_1
XANTENNA__12410__B1 net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12392_ net2168 net183 net270 vssd1 vssd1 vccd1 vccd1 _01103_ sky130_fd_sc_hd__mux2_1
X_14131_ clknet_leaf_18_clk final_design.vga.h_next_count\[0\] net1114 vssd1 vssd1
+ vccd1 vccd1 final_design.VGA_data_control.h_count\[0\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__11479__S net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11343_ net737 _03859_ _06033_ vssd1 vssd1 vccd1 vccd1 _06034_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_82_1861 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14062_ clknet_leaf_16_clk _00024_ net1091 vssd1 vssd1 vccd1 vccd1 final_design.uart.BAUD_counter\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_11274_ net426 net556 _05973_ net314 net1797 vssd1 vssd1 vccd1 vccd1 _00290_ sky130_fd_sc_hd__a32o_1
XFILLER_0_39_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13013_ clknet_leaf_56_clk _00244_ net1145 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_10225_ final_design.uart.BAUD_counter\[9\] _05103_ vssd1 vssd1 vccd1 vccd1 _05104_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_24_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10156_ net1048 _05050_ _05045_ vssd1 vssd1 vccd1 vccd1 _05053_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_7_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold5 final_design.cpu.reg_window\[14\] vssd1 vssd1 vccd1 vccd1 net1347 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12103__S net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12477__B1 net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09192__B _03649_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10087_ _04999_ _05002_ vssd1 vssd1 vccd1 vccd1 _05003_ sky130_fd_sc_hd__or2_1
XANTENNA__10412__A _03321_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13915_ clknet_leaf_65_clk _01146_ net1070 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[903\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13582__CLK clknet_leaf_45_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload3_A clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13846_ clknet_leaf_59_clk _01077_ net1125 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[834\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13777_ clknet_leaf_34_clk _01008_ net1242 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[765\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10989_ _01360_ _03844_ net1059 vssd1 vssd1 vccd1 vccd1 _05715_ sky130_fd_sc_hd__mux2_1
XANTENNA__12244__A3 net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12728_ _06363_ _06361_ final_design.VGA_data_control.v_count\[1\] vssd1 vssd1 vccd1
+ vccd1 _06369_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12659_ final_design.VGA_data_control.ready_data\[17\] net1020 net975 final_design.data_from_mem\[17\]
+ vssd1 vssd1 vccd1 vccd1 _06317_ sky130_fd_sc_hd__a22o_1
XFILLER_0_44_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_2809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11204__A1 net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12401__B1 net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14088__CLK clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold405 final_design.cpu.reg_window\[754\] vssd1 vssd1 vccd1 vccd1 net1747 sky130_fd_sc_hd__dlygate4sd3_1
Xhold416 final_design.cpu.reg_window\[150\] vssd1 vssd1 vccd1 vccd1 net1758 sky130_fd_sc_hd__dlygate4sd3_1
Xhold427 final_design.cpu.reg_window\[659\] vssd1 vssd1 vccd1 vccd1 net1769 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold438 final_design.cpu.reg_window\[751\] vssd1 vssd1 vccd1 vccd1 net1780 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07168__A net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold449 final_design.cpu.reg_window\[154\] vssd1 vssd1 vccd1 vccd1 net1791 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_46_1480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_1322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09870_ _03520_ _03521_ _03554_ _03555_ _04046_ vssd1 vssd1 vccd1 vccd1 _04789_ sky130_fd_sc_hd__o311a_1
Xfanout907 net910 vssd1 vssd1 vccd1 vccd1 net907 sky130_fd_sc_hd__clkbuf_2
Xfanout918 net919 vssd1 vssd1 vccd1 vccd1 net918 sky130_fd_sc_hd__clkbuf_4
Xfanout929 net932 vssd1 vssd1 vccd1 vccd1 net929 sky130_fd_sc_hd__clkbuf_4
X_08821_ _03666_ _03771_ _03667_ vssd1 vssd1 vccd1 vccd1 _03772_ sky130_fd_sc_hd__a21o_1
XANTENNA__12180__A2 net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10191__A1 net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13925__CLK clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1105 final_design.cpu.reg_window\[629\] vssd1 vssd1 vccd1 vccd1 net2447 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07592__C1 net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1116 final_design.cpu.reg_window\[101\] vssd1 vssd1 vccd1 vccd1 net2458 sky130_fd_sc_hd__dlygate4sd3_1
X_08752_ final_design.CPU_instr_adr\[5\] net666 _01659_ vssd1 vssd1 vccd1 vccd1 _03703_
+ sky130_fd_sc_hd__and3_1
Xhold1127 final_design.cpu.reg_window\[533\] vssd1 vssd1 vccd1 vccd1 net2469 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12468__B1 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1138 final_design.cpu.reg_window\[299\] vssd1 vssd1 vccd1 vccd1 net2480 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1149 final_design.cpu.reg_window\[811\] vssd1 vssd1 vccd1 vccd1 net2491 sky130_fd_sc_hd__dlygate4sd3_1
X_07703_ _02650_ _02651_ _02652_ _02653_ net688 net704 vssd1 vssd1 vccd1 vccd1 _02654_
+ sky130_fd_sc_hd__mux4_1
X_08683_ _03632_ _03633_ _02510_ vssd1 vssd1 vccd1 vccd1 _03634_ sky130_fd_sc_hd__a21o_1
XFILLER_0_59_1885 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07634_ final_design.cpu.reg_window\[28\] final_design.cpu.reg_window\[60\] net866
+ vssd1 vssd1 vccd1 vccd1 _02585_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07565_ final_design.cpu.reg_window\[351\] final_design.cpu.reg_window\[383\] net859
+ vssd1 vssd1 vccd1 vccd1 _02516_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout342_A net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12235__A3 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1084_A net1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09304_ net595 _03514_ _03516_ _02503_ vssd1 vssd1 vccd1 vccd1 _04223_ sky130_fd_sc_hd__o211a_2
X_06516_ net1039 net994 net991 final_design.reqhand.instruction\[3\] vssd1 vssd1 vccd1
+ vccd1 _01467_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_17_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07496_ _02101_ _02446_ vssd1 vssd1 vccd1 vccd1 _02447_ sky130_fd_sc_hd__or2_1
XANTENNA__13305__CLK clknet_leaf_56_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07111__A2 net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11994__A2 net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09235_ _03326_ _03357_ _03324_ vssd1 vssd1 vccd1 vccd1 _04154_ sky130_fd_sc_hd__a21oi_2
X_06447_ _01397_ _01400_ vssd1 vssd1 vccd1 vccd1 _01401_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_20_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout228_X net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout607_A _02514_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1801 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1157 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12777__8 clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 net1318 sky130_fd_sc_hd__inv_2
XANTENNA__07777__S net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09166_ net495 net481 vssd1 vssd1 vccd1 vccd1 _04085_ sky130_fd_sc_hd__nand2_1
XFILLER_0_50_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08298__S1 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_1845 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08117_ net611 _03065_ _03066_ _02058_ vssd1 vssd1 vccd1 vccd1 _03068_ sky130_fd_sc_hd__a211o_1
XFILLER_0_9_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11600__B net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13455__CLK clknet_leaf_42_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09097_ _03711_ _03719_ vssd1 vssd1 vccd1 vccd1 _04020_ sky130_fd_sc_hd__xor2_1
XFILLER_0_66_1889 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08048_ final_design.cpu.reg_window\[466\] final_design.cpu.reg_window\[498\] net844
+ vssd1 vssd1 vccd1 vccd1 _02999_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold950 final_design.cpu.reg_window\[358\] vssd1 vssd1 vccd1 vccd1 net2292 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout976_A _06299_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold961 final_design.cpu.reg_window\[195\] vssd1 vssd1 vccd1 vccd1 net2303 sky130_fd_sc_hd__dlygate4sd3_1
Xhold972 final_design.cpu.reg_window\[757\] vssd1 vssd1 vccd1 vccd1 net2314 sky130_fd_sc_hd__dlygate4sd3_1
Xhold983 final_design.cpu.reg_window\[509\] vssd1 vssd1 vccd1 vccd1 net2325 sky130_fd_sc_hd__dlygate4sd3_1
Xhold994 final_design.reqhand.instruction\[20\] vssd1 vssd1 vccd1 vccd1 net2336 sky130_fd_sc_hd__dlygate4sd3_1
X_10010_ _02326_ net452 _04238_ net465 vssd1 vssd1 vccd1 vccd1 _04929_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_38_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout764_X net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09999_ net451 _04907_ _04916_ net727 vssd1 vssd1 vccd1 vccd1 _04918_ sky130_fd_sc_hd__a211o_2
XANTENNA__06710__A _01658_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09324__A0 _04234_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1805 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11961_ _06163_ net281 net404 net1661 vssd1 vssd1 vccd1 vccd1 _00694_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout931_X net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08222__S1 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11762__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10912_ net669 _05627_ _05638_ net962 _05641_ vssd1 vssd1 vccd1 vccd1 _05642_ sky130_fd_sc_hd__o221a_1
X_13700_ clknet_leaf_54_clk _00931_ net1179 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[688\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_1849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07812__Y _02763_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11682__A1 net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11892_ net244 net2158 net272 vssd1 vssd1 vccd1 vccd1 _00634_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06709__X _01660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13631_ clknet_leaf_10_clk _00862_ net1102 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[619\]
+ sky130_fd_sc_hd__dfrtp_1
X_10843_ final_design.CPU_instr_adr\[19\] net1000 _05572_ net1055 vssd1 vssd1 vccd1
+ vccd1 _05576_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_15_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09627__A1 _04046_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12226__A3 net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13562_ clknet_leaf_1_clk _00793_ net1075 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[550\]
+ sky130_fd_sc_hd__dfrtp_1
X_10774_ net75 net1044 vssd1 vssd1 vccd1 vccd1 _05510_ sky130_fd_sc_hd__and2_1
XANTENNA__09722__S1 net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07733__S0 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12513_ _06175_ net342 net326 net1614 vssd1 vssd1 vccd1 vccd1 _01218_ sky130_fd_sc_hd__a22o_1
XANTENNA__11985__A2 net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_234 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13493_ clknet_leaf_56_clk _00724_ net1144 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[481\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12444_ net1708 net213 net334 vssd1 vssd1 vccd1 vccd1 _01151_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12890__Q final_design.data_from_mem\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12375_ net2512 net214 net268 vssd1 vssd1 vccd1 vccd1 _01086_ sky130_fd_sc_hd__mux2_1
XANTENNA__08602__A2 _03550_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14114_ clknet_leaf_14_clk _01311_ net1107 vssd1 vssd1 vccd1 vccd1 final_design.reqhand.data_from_UART\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_11326_ net661 _03874_ net733 vssd1 vssd1 vccd1 vccd1 _06019_ sky130_fd_sc_hd__o21a_1
XFILLER_0_61_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13948__CLK clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14045_ clknet_leaf_16_clk _00037_ net1092 vssd1 vssd1 vccd1 vccd1 final_design.uart.BAUD_counter\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_11257_ net649 net209 vssd1 vssd1 vccd1 vccd1 _05959_ sky130_fd_sc_hd__and2_1
XFILLER_0_66_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10208_ _05093_ net800 _05092_ vssd1 vssd1 vccd1 vccd1 _00028_ sky130_fd_sc_hd__and3b_1
XPHY_EDGE_ROW_8_Left_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06620__A _01567_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11188_ net648 net224 vssd1 vssd1 vccd1 vccd1 _05898_ sky130_fd_sc_hd__and2_1
XANTENNA__11238__A net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10139_ final_design.vga.h_current_state\[0\] final_design.VGA_data_control.h_count\[8\]
+ final_design.VGA_data_control.h_count\[9\] final_design.vga.h_current_state\[1\]
+ vssd1 vssd1 vccd1 vccd1 _05041_ sky130_fd_sc_hd__or4b_1
XANTENNA__08118__A1 net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11672__S net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06619__X _01570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13328__CLK clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1845 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11244__Y _05947_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13829_ clknet_leaf_51_clk _01060_ net1173 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[817\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_4_1709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1880 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12217__A3 net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1889 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07350_ final_design.cpu.reg_window\[323\] final_design.cpu.reg_window\[355\] net912
+ vssd1 vssd1 vccd1 vccd1 _02301_ sky130_fd_sc_hd__mux2_1
XANTENNA__11976__A2 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07281_ _02228_ _02229_ _02230_ _02231_ net767 net787 vssd1 vssd1 vccd1 vccd1 _02232_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__13478__CLK clknet_leaf_51_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09020_ net2524 net1017 _03948_ _03952_ vssd1 vssd1 vccd1 vccd1 _00224_ sky130_fd_sc_hd__a22o_1
XFILLER_0_32_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11189__B1 net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11728__A2 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold202 final_design.VGA_data_control.ready_data\[10\] vssd1 vssd1 vccd1 vccd1 net1544
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_1406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold213 final_design.VGA_data_control.data_to_VGA\[4\] vssd1 vssd1 vccd1 vccd1 net1555
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold224 final_design.cpu.reg_window\[176\] vssd1 vssd1 vccd1 vccd1 net1566 sky130_fd_sc_hd__dlygate4sd3_1
Xhold235 final_design.cpu.reg_window\[971\] vssd1 vssd1 vccd1 vccd1 net1577 sky130_fd_sc_hd__dlygate4sd3_1
Xhold246 final_design.cpu.reg_window\[71\] vssd1 vssd1 vccd1 vccd1 net1588 sky130_fd_sc_hd__dlygate4sd3_1
Xhold257 final_design.cpu.reg_window\[57\] vssd1 vssd1 vccd1 vccd1 net1599 sky130_fd_sc_hd__dlygate4sd3_1
Xhold268 final_design.cpu.reg_window\[557\] vssd1 vssd1 vccd1 vccd1 net1610 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold279 final_design.cpu.reg_window\[589\] vssd1 vssd1 vccd1 vccd1 net1621 sky130_fd_sc_hd__dlygate4sd3_1
X_09922_ _04341_ _04840_ vssd1 vssd1 vccd1 vccd1 _04841_ sky130_fd_sc_hd__or2_1
Xfanout704 net706 vssd1 vssd1 vccd1 vccd1 net704 sky130_fd_sc_hd__buf_4
Xfanout715 _01721_ vssd1 vssd1 vccd1 vccd1 net715 sky130_fd_sc_hd__clkbuf_4
Xfanout726 _01493_ vssd1 vssd1 vccd1 vccd1 net726 sky130_fd_sc_hd__clkbuf_4
Xfanout737 net738 vssd1 vssd1 vccd1 vccd1 net737 sky130_fd_sc_hd__buf_2
X_09853_ _04741_ _04771_ net450 vssd1 vssd1 vccd1 vccd1 _04772_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07626__A _01570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08221__S net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout748 _01438_ vssd1 vssd1 vccd1 vccd1 net748 sky130_fd_sc_hd__buf_2
XANTENNA__11361__B1 _06049_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout759 net760 vssd1 vssd1 vccd1 vccd1 net759 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout292_A net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14103__CLK clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08804_ final_design.CPU_instr_adr\[23\] _01722_ vssd1 vssd1 vccd1 vccd1 _03755_
+ sky130_fd_sc_hd__or2_1
X_09784_ _04657_ _04678_ _04679_ _04702_ vssd1 vssd1 vccd1 vccd1 _04703_ sky130_fd_sc_hd__and4_1
XANTENNA__13055__RESET_B net1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06996_ _01943_ _01944_ _01945_ _01946_ net766 net785 vssd1 vssd1 vccd1 vccd1 _01947_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_52_1982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09306__B1 net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08735_ final_design.CPU_instr_adr\[13\] _02030_ vssd1 vssd1 vccd1 vccd1 _03686_
+ sky130_fd_sc_hd__or2_1
XANTENNA__09841__A _04072_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout557_A net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08666_ _01487_ _03615_ _03616_ _02094_ vssd1 vssd1 vccd1 vccd1 _03617_ sky130_fd_sc_hd__o22a_4
XANTENNA__11664__A1 net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07617_ _02564_ _02565_ _02566_ _02567_ net688 net705 vssd1 vssd1 vccd1 vccd1 _02568_
+ sky130_fd_sc_hd__mux4_1
X_08597_ net717 _03547_ vssd1 vssd1 vccd1 vccd1 _03548_ sky130_fd_sc_hd__or2_1
XANTENNA__12208__A3 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout345_X net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07548_ final_design.cpu.reg_window\[543\] final_design.cpu.reg_window\[575\] net937
+ vssd1 vssd1 vccd1 vccd1 _02499_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_46_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12613__B1 net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09085__A2 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07715__S0 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11967__A2 net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_42_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07479_ _02364_ _02429_ vssd1 vssd1 vccd1 vccd1 _02430_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout512_X net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09218_ _03068_ _03099_ _03100_ vssd1 vssd1 vccd1 vccd1 _04137_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_17_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_1590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10490_ net1053 _05237_ net1001 net1018 vssd1 vssd1 vccd1 vccd1 _05240_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__12845__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06705__A net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07300__S net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_930 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09149_ _04056_ _04067_ vssd1 vssd1 vccd1 vccd1 _04068_ sky130_fd_sc_hd__or2_1
XFILLER_0_32_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12160_ net178 net2395 net386 vssd1 vssd1 vccd1 vccd1 _00881_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_9_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout881_X net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11757__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11111_ _05830_ net1052 vssd1 vssd1 vccd1 vccd1 _05831_ sky130_fd_sc_hd__and2b_1
X_12091_ net584 _06075_ net512 net394 net2023 vssd1 vssd1 vccd1 vccd1 _00816_ sky130_fd_sc_hd__a32o_1
Xhold780 final_design.cpu.reg_window\[556\] vssd1 vssd1 vccd1 vccd1 net2122 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_6_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold791 final_design.cpu.reg_window\[503\] vssd1 vssd1 vccd1 vccd1 net2133 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09545__B1 net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11042_ _05760_ _05764_ vssd1 vssd1 vccd1 vccd1 _05766_ sky130_fd_sc_hd__and2b_1
XANTENNA__11352__B1 net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input20_A DAT_I[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12993_ net1324 _00224_ net1194 vssd1 vssd1 vccd1 vccd1 final_design.CPU_instr_adr\[13\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_77_1793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06586__S net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11944_ _06145_ net292 net410 net2080 vssd1 vssd1 vccd1 vccd1 _00679_ sky130_fd_sc_hd__a22o_1
XANTENNA__12885__Q final_design.data_from_mem\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_1900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11875_ net188 net554 vssd1 vssd1 vccd1 vccd1 _06245_ sky130_fd_sc_hd__and2_1
X_10826_ _05559_ vssd1 vssd1 vccd1 vccd1 _05560_ sky130_fd_sc_hd__inv_2
X_13614_ clknet_leaf_44_clk _00845_ net1208 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[602\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11407__A1 net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13620__CLK clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11958__A2 net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10757_ final_design.CPU_instr_adr\[15\] net1000 _05490_ net1055 vssd1 vssd1 vccd1
+ vccd1 _05494_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__12080__A1 net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13545_ clknet_leaf_37_clk _00776_ net1228 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[533\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09198__A net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06834__A1 net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13476_ clknet_leaf_54_clk _00707_ net1179 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[464\]
+ sky130_fd_sc_hd__dfrtp_1
X_10688_ net70 final_design.VGA_adr\[9\] _05426_ vssd1 vssd1 vccd1 vccd1 _05428_ sky130_fd_sc_hd__or3_1
XFILLER_0_36_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13770__CLK clknet_leaf_60_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12427_ _06114_ net357 net340 net2472 vssd1 vssd1 vccd1 vccd1 _01136_ sky130_fd_sc_hd__a22o_1
XANTENNA__10918__B1 net1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08131__S0 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12358_ net2241 net363 net356 _06061_ vssd1 vssd1 vccd1 vccd1 _01070_ sky130_fd_sc_hd__a22o_1
XANTENNA__09926__A _04124_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11591__B1 net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11309_ net2542 net315 net422 _06004_ vssd1 vssd1 vccd1 vccd1 _00294_ sky130_fd_sc_hd__a22o_1
XANTENNA__14126__CLK clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12289_ net578 _06219_ net510 net370 net1857 vssd1 vssd1 vccd1 vccd1 _01004_ sky130_fd_sc_hd__a32o_1
XFILLER_0_77_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14028_ clknet_leaf_46_clk _01259_ net1214 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[1016\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06850_ _01797_ _01798_ _01799_ _01800_ net777 net794 vssd1 vssd1 vccd1 vccd1 _01801_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__13150__CLK clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06996__S1 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire525_A _03549_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06781_ final_design.cpu.reg_window\[86\] final_design.cpu.reg_window\[118\] net918
+ vssd1 vssd1 vccd1 vccd1 _01732_ sky130_fd_sc_hd__mux2_1
X_08520_ final_design.cpu.reg_window\[770\] final_design.cpu.reg_window\[802\] net833
+ vssd1 vssd1 vccd1 vccd1 _03471_ sky130_fd_sc_hd__mux2_1
XANTENNA__10449__A2 net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11646__A1 net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06496__S net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_19_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08451_ net717 _03401_ vssd1 vssd1 vccd1 vccd1 _03402_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_19_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_44_clk_X clknet_leaf_44_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07402_ final_design.cpu.reg_window\[514\] final_design.cpu.reg_window\[546\] net913
+ vssd1 vssd1 vccd1 vccd1 _02353_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08382_ _03329_ _03330_ _03331_ _03332_ net679 net692 vssd1 vssd1 vccd1 vccd1 _03333_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__12868__CLK clknet_leaf_25_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07333_ final_design.cpu.reg_window\[772\] final_design.cpu.reg_window\[804\] net900
+ vssd1 vssd1 vccd1 vccd1 _02284_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11949__A2 net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07078__A1 final_design.data_from_mem\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07173__S1 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10737__A1_N net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07264_ _02213_ _02214_ vssd1 vssd1 vccd1 vccd1 _02215_ sky130_fd_sc_hd__and2b_1
XFILLER_0_61_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_59_clk_X clknet_leaf_59_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12246__B net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07120__S net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09003_ _02002_ _02450_ vssd1 vssd1 vccd1 vccd1 _03937_ sky130_fd_sc_hd__and2_1
X_12783__14 clknet_leaf_28_clk vssd1 vssd1 vccd1 vccd1 net1324 sky130_fd_sc_hd__inv_2
XFILLER_0_14_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07195_ final_design.cpu.reg_window\[905\] final_design.cpu.reg_window\[937\] net891
+ vssd1 vssd1 vccd1 vccd1 _02146_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_1913 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout305_A _06125_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1047_A final_design.VGA_adr\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_1501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1214_A net1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout501 _06264_ vssd1 vssd1 vccd1 vccd1 net501 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_35_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09905_ _04819_ _04821_ _04823_ _04820_ vssd1 vssd1 vccd1 vccd1 _04824_ sky130_fd_sc_hd__or4b_1
Xfanout512 net513 vssd1 vssd1 vccd1 vccd1 net512 sky130_fd_sc_hd__clkbuf_4
Xfanout523 net524 vssd1 vssd1 vccd1 vccd1 net523 sky130_fd_sc_hd__buf_8
Xfanout534 _02184_ vssd1 vssd1 vccd1 vccd1 net534 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_50_1908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout674_A net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout545 _01908_ vssd1 vssd1 vccd1 vccd1 net545 sky130_fd_sc_hd__buf_2
XANTENNA_fanout295_X net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout556 net562 vssd1 vssd1 vccd1 vccd1 net556 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_50_1919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout567 net568 vssd1 vssd1 vccd1 vccd1 net567 sky130_fd_sc_hd__buf_2
X_09836_ _04606_ _04711_ net471 vssd1 vssd1 vccd1 vccd1 _04755_ sky130_fd_sc_hd__mux2_1
Xfanout578 net587 vssd1 vssd1 vccd1 vccd1 net578 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout1002_X net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout589 net590 vssd1 vssd1 vccd1 vccd1 net589 sky130_fd_sc_hd__buf_2
X_06979_ net756 _01929_ vssd1 vssd1 vccd1 vccd1 _01930_ sky130_fd_sc_hd__or2_2
XANTENNA_fanout841_A net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09767_ net490 _04685_ net318 vssd1 vssd1 vccd1 vccd1 _04686_ sky130_fd_sc_hd__o21a_1
XFILLER_0_38_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout939_A net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08189__S0 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08718_ final_design.CPU_instr_adr\[20\] _01823_ vssd1 vssd1 vccd1 vccd1 _03669_
+ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_1_241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13643__CLK clknet_leaf_52_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_1_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09698_ _03100_ net440 net441 _03099_ vssd1 vssd1 vccd1 vccd1 _04617_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_29_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1917 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_1837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08649_ _02769_ _03597_ _03598_ vssd1 vssd1 vccd1 vccd1 _03600_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_48_1848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout727_X net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11660_ net582 net423 _06187_ net300 net1538 vssd1 vssd1 vccd1 vccd1 _00462_ sky130_fd_sc_hd__a32o_1
XFILLER_0_33_1652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10611_ _05334_ _05337_ _05353_ vssd1 vssd1 vccd1 vccd1 _05355_ sky130_fd_sc_hd__or3_1
XANTENNA__13793__CLK clknet_leaf_47_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11591_ net581 net423 _06151_ net305 net1627 vssd1 vssd1 vccd1 vccd1 _00429_ sky130_fd_sc_hd__a32o_1
XANTENNA__06706__Y _01657_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13330_ clknet_leaf_38_clk _00561_ net1189 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[318\]
+ sky130_fd_sc_hd__dfrtp_1
X_10542_ net95 final_design.VGA_adr\[3\] vssd1 vssd1 vccd1 vccd1 _05289_ sky130_fd_sc_hd__xor2_1
XANTENNA__11270__C1 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13261_ clknet_leaf_48_clk _00492_ net1200 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[249\]
+ sky130_fd_sc_hd__dfrtp_1
X_10473_ final_design.CPU_instr_adr\[1\] net79 net1053 vssd1 vssd1 vccd1 vccd1 _05224_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__13023__CLK clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14149__CLK clknet_leaf_15_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12212_ net558 _06140_ net502 net376 net2106 vssd1 vssd1 vccd1 vccd1 _00930_ sky130_fd_sc_hd__a32o_1
X_13192_ clknet_leaf_35_clk _00423_ net1237 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[180\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input68_A memory_size[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10376__B2 final_design.data_from_mem\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11573__B1 net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11487__S net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12143_ net210 net2404 net386 vssd1 vssd1 vccd1 vccd1 _00864_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13173__CLK clknet_leaf_57_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12074_ net559 _05952_ net503 net392 net2122 vssd1 vssd1 vccd1 vccd1 _00799_ sky130_fd_sc_hd__a32o_1
XFILLER_0_47_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10404__B _05181_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11325__B1 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11025_ _05729_ _05733_ _05749_ vssd1 vssd1 vccd1 vccd1 _05750_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_70_2580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_70_2591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11876__B2 net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06978__S1 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08809__B _01788_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11628__A1 net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12111__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12976_ clknet_leaf_20_clk _00001_ net1160 vssd1 vssd1 vccd1 vccd1 final_design.reqhand.current_client\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_59_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11927_ net2556 net408 _06253_ net427 vssd1 vssd1 vccd1 vccd1 _00663_ sky130_fd_sc_hd__a22o_1
XFILLER_0_75_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_64_2384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11858_ net213 net553 vssd1 vssd1 vccd1 vccd1 _06241_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_64_2395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_2248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_2259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10809_ _05522_ _05540_ vssd1 vssd1 vccd1 vccd1 _05544_ sky130_fd_sc_hd__and2_1
XANTENNA_19 _06228_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12053__A1 net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11789_ net2313 net412 _06233_ net427 vssd1 vssd1 vccd1 vccd1 _00545_ sky130_fd_sc_hd__a22o_1
XANTENNA__07155__S1 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13528_ clknet_leaf_65_clk _00759_ net1070 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[516\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11800__B2 net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13459_ clknet_leaf_40_clk _00690_ net1211 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[447\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_11_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_11_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07875__S net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12356__A2 net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput104 net104 vssd1 vssd1 vccd1 vccd1 ADR_O[12] sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_58_2177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput115 net115 vssd1 vssd1 vccd1 vccd1 ADR_O[22] sky130_fd_sc_hd__clkbuf_4
XANTENNA__13516__CLK clknet_leaf_46_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_58_2188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput126 net126 vssd1 vssd1 vccd1 vccd1 ADR_O[3] sky130_fd_sc_hd__clkbuf_4
XANTENNA__10367__B2 final_design.data_from_mem\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_2199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput137 net137 vssd1 vssd1 vccd1 vccd1 DAT_O[12] sky130_fd_sc_hd__buf_2
Xoutput148 net148 vssd1 vssd1 vccd1 vccd1 DAT_O[22] sky130_fd_sc_hd__buf_2
Xoutput159 net159 vssd1 vssd1 vccd1 vccd1 DAT_O[3] sky130_fd_sc_hd__buf_2
XANTENNA__07783__A2 _02731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07951_ _02838_ _02901_ vssd1 vssd1 vccd1 vccd1 _02902_ sky130_fd_sc_hd__and2_1
XFILLER_0_23_1854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06902_ net747 net664 _01821_ vssd1 vssd1 vccd1 vccd1 _01853_ sky130_fd_sc_hd__o21ai_4
XANTENNA__13666__CLK clknet_leaf_11_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07882_ net616 _02830_ _02831_ net549 vssd1 vssd1 vccd1 vccd1 _02833_ sky130_fd_sc_hd__a211oi_1
X_09621_ _04342_ _04539_ vssd1 vssd1 vccd1 vccd1 _04540_ sky130_fd_sc_hd__and2b_1
X_06833_ net884 _01777_ _01783_ _01765_ _01771_ vssd1 vssd1 vccd1 vccd1 _01784_ sky130_fd_sc_hd__a32oi_4
XFILLER_0_78_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09552_ _03590_ _04143_ _04157_ _03587_ vssd1 vssd1 vccd1 vccd1 _04471_ sky130_fd_sc_hd__o31a_1
X_06764_ _01711_ _01712_ _01713_ _01714_ net772 net784 vssd1 vssd1 vccd1 vccd1 _01715_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__09288__A2 _03550_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08503_ net608 _03450_ _03451_ vssd1 vssd1 vccd1 vccd1 _03454_ sky130_fd_sc_hd__a21o_1
XFILLER_0_37_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09483_ net544 net542 net541 net540 net459 net469 vssd1 vssd1 vccd1 vccd1 _04402_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_17_1647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06695_ final_design.cpu.reg_window\[793\] final_design.cpu.reg_window\[825\] net931
+ vssd1 vssd1 vccd1 vccd1 _01646_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09693__C1 _03649_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout255_A net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08434_ _02267_ net597 vssd1 vssd1 vccd1 vccd1 _03385_ sky130_fd_sc_hd__and2_1
XFILLER_0_19_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1347 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08365_ final_design.cpu.reg_window\[647\] final_design.cpu.reg_window\[679\] net809
+ vssd1 vssd1 vccd1 vccd1 _03316_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_24_clk_A clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13046__CLK clknet_leaf_61_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11799__C _06024_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout422_A _05877_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1164_A net1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07316_ net666 _01659_ vssd1 vssd1 vccd1 vccd1 _02267_ sky130_fd_sc_hd__nand2_1
XANTENNA__12595__A2 net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08296_ final_design.cpu.reg_window\[713\] final_design.cpu.reg_window\[745\] net808
+ vssd1 vssd1 vccd1 vccd1 _03247_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_1071 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09460__A2 _04373_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07247_ _02194_ _02195_ _02196_ _02197_ net766 net785 vssd1 vssd1 vccd1 vccd1 _02198_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_5_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout308_X net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12347__A2 net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09748__B1 net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13196__CLK clknet_leaf_45_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_39_clk_A clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06542__X _01493_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07178_ _02127_ _02128_ vssd1 vssd1 vccd1 vccd1 _02129_ sky130_fd_sc_hd__nand2_1
XFILLER_0_63_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10358__A1 net31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout791_A net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11555__B1 net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout889_A net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout320 _04073_ vssd1 vssd1 vccd1 vccd1 net320 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout677_X net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11307__B1 net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout331 _06283_ vssd1 vssd1 vccd1 vccd1 net331 sky130_fd_sc_hd__buf_4
Xfanout342 net343 vssd1 vssd1 vccd1 vccd1 net342 sky130_fd_sc_hd__clkbuf_4
Xfanout353 net359 vssd1 vssd1 vccd1 vccd1 net353 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09515__A3 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout364 net365 vssd1 vssd1 vccd1 vccd1 net364 sky130_fd_sc_hd__buf_4
Xfanout375 _06272_ vssd1 vssd1 vccd1 vccd1 net375 sky130_fd_sc_hd__buf_4
Xfanout386 net387 vssd1 vssd1 vccd1 vccd1 net386 sky130_fd_sc_hd__clkbuf_8
Xfanout397 _06261_ vssd1 vssd1 vccd1 vccd1 net397 sky130_fd_sc_hd__buf_4
X_09819_ _03294_ _03569_ vssd1 vssd1 vccd1 vccd1 _04738_ sky130_fd_sc_hd__nand2_1
X_12830_ net1395 vssd1 vssd1 vccd1 vccd1 _00271_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_74_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12761_ _06339_ _06391_ vssd1 vssd1 vccd1 vccd1 _06397_ sky130_fd_sc_hd__or2_1
XANTENNA__12283__A1 net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08487__B1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11712_ net435 net585 _06214_ net296 net1629 vssd1 vssd1 vccd1 vccd1 _00487_ sky130_fd_sc_hd__a32o_1
X_12692_ _05008_ net954 _05059_ net796 final_design.VGA_adr\[1\] vssd1 vssd1 vccd1
+ vccd1 _01348_ sky130_fd_sc_hd__a32o_1
XANTENNA__10833__A2 net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08645__A _02772_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11643_ net200 net631 vssd1 vssd1 vccd1 vccd1 _06179_ sky130_fd_sc_hd__and2_1
XANTENNA__12035__A1 net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10046__B1 _04421_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08334__S0 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09987__B1 _04905_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12586__A2 net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11574_ net201 net635 vssd1 vssd1 vccd1 vccd1 _06143_ sky130_fd_sc_hd__and2_1
XFILLER_0_80_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13539__CLK clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09179__C net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput17 DAT_I[23] vssd1 vssd1 vccd1 vccd1 net17 sky130_fd_sc_hd__clkbuf_1
Xinput28 DAT_I[4] vssd1 vssd1 vccd1 vccd1 net28 sky130_fd_sc_hd__clkbuf_1
Xinput39 mem_adr_start[12] vssd1 vssd1 vccd1 vccd1 net39 sky130_fd_sc_hd__clkbuf_1
X_10525_ _05270_ _05271_ _05272_ vssd1 vssd1 vccd1 vccd1 _05273_ sky130_fd_sc_hd__and3_1
X_13313_ clknet_leaf_49_clk _00544_ net1186 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[301\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_1789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12338__A2 net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13244_ clknet_leaf_3_clk _00475_ net1066 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[232\]
+ sky130_fd_sc_hd__dfrtp_1
X_10456_ _02602_ net593 vssd1 vssd1 vccd1 vccd1 _05212_ sky130_fd_sc_hd__nor2_1
XFILLER_0_66_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11010__A2 net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13175_ clknet_leaf_5_clk _00406_ net1082 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[163\]
+ sky130_fd_sc_hd__dfrtp_1
X_10387_ net1389 net1028 _05174_ vssd1 vssd1 vccd1 vccd1 _00137_ sky130_fd_sc_hd__a21bo_1
XANTENNA__13689__CLK clknet_leaf_57_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10415__A _03287_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12106__S net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_72_2653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_2030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12126_ net1917 net176 net390 vssd1 vssd1 vccd1 vccd1 _00850_ sky130_fd_sc_hd__mux2_1
XANTENNA__11561__A3 _06136_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1188 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06973__B1 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12057_ net1881 net178 net398 vssd1 vssd1 vccd1 vccd1 _00785_ sky130_fd_sc_hd__mux2_1
X_11008_ _05711_ _05731_ _05732_ net1005 vssd1 vssd1 vccd1 vccd1 _05734_ sky130_fd_sc_hd__a31o_1
XANTENNA__12510__A2 net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07073__S0 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1901 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_2446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11077__A2 net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12274__A1 net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12959_ clknet_leaf_32_clk _00197_ net1233 vssd1 vssd1 vccd1 vccd1 net117 sky130_fd_sc_hd__dfrtp_1
XANTENNA__13069__CLK clknet_leaf_44_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06480_ final_design.cpu.reg_window\[94\] final_design.cpu.reg_window\[126\] net936
+ vssd1 vssd1 vccd1 vccd1 _01431_ sky130_fd_sc_hd__mux2_1
XANTENNA__08555__A net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09978__B1 _04046_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08150_ _03099_ _03100_ vssd1 vssd1 vccd1 vccd1 _03101_ sky130_fd_sc_hd__nor2_1
X_07101_ final_design.cpu.reg_window\[716\] final_design.cpu.reg_window\[748\] net894
+ vssd1 vssd1 vccd1 vccd1 _02052_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08081_ net547 _02996_ _03024_ _02993_ _01850_ vssd1 vssd1 vccd1 vccd1 _03032_ sky130_fd_sc_hd__o32a_1
XANTENNA__12906__CLK clknet_leaf_61_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07032_ final_design.cpu.reg_window\[846\] final_design.cpu.reg_window\[878\] net906
+ vssd1 vssd1 vccd1 vccd1 _01983_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07205__A1 net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08983_ net258 _03918_ net1016 vssd1 vssd1 vccd1 vccd1 _03920_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_47_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07934_ final_design.cpu.reg_window\[918\] final_design.cpu.reg_window\[950\] net841
+ vssd1 vssd1 vccd1 vccd1 _02885_ sky130_fd_sc_hd__mux2_1
XANTENNA__09833__B net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12501__A2 net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07865_ _02812_ _02813_ _02814_ _02815_ net687 net705 vssd1 vssd1 vccd1 vccd1 _02816_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__10512__B2 net1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_1124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout372_A net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09604_ net486 _04437_ vssd1 vssd1 vccd1 vccd1 _04523_ sky130_fd_sc_hd__nand2_1
XANTENNA__08181__A2 net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06816_ final_design.cpu.reg_window\[277\] final_design.cpu.reg_window\[309\] net938
+ vssd1 vssd1 vccd1 vccd1 _01767_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07796_ final_design.cpu.reg_window\[217\] final_design.cpu.reg_window\[249\] net855
+ vssd1 vssd1 vccd1 vccd1 _02747_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09535_ _04188_ _04453_ vssd1 vssd1 vccd1 vccd1 _04454_ sky130_fd_sc_hd__and2_1
XANTENNA__12265__A1 net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06747_ final_design.cpu.reg_window\[87\] final_design.cpu.reg_window\[119\] net929
+ vssd1 vssd1 vccd1 vccd1 _01698_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout258_X net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout637_A _06123_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09466_ _04382_ _04383_ net729 _04381_ vssd1 vssd1 vccd1 vccd1 _04385_ sky130_fd_sc_hd__o211a_1
XFILLER_0_52_1346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06678_ net744 _01628_ vssd1 vssd1 vccd1 vccd1 _01629_ sky130_fd_sc_hd__and2_1
XFILLER_0_59_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08417_ final_design.cpu.reg_window\[197\] final_design.cpu.reg_window\[229\] net838
+ vssd1 vssd1 vccd1 vccd1 _03368_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09397_ net463 _04080_ _04315_ net473 vssd1 vssd1 vccd1 vccd1 _04316_ sky130_fd_sc_hd__o211a_1
XANTENNA__12783__14_A clknet_leaf_28_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout425_X net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1167_X net1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08184__B net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08348_ final_design.cpu.reg_window\[263\] final_design.cpu.reg_window\[295\] net811
+ vssd1 vssd1 vccd1 vccd1 _03299_ sky130_fd_sc_hd__mux2_1
XANTENNA__09969__B1 net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11776__B1 net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1707 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08279_ _03229_ vssd1 vssd1 vccd1 vccd1 _03230_ sky130_fd_sc_hd__inv_2
X_10310_ final_design.VGA_data_control.h_count\[4\] final_design.VGA_data_control.h_count\[5\]
+ _05153_ _05163_ vssd1 vssd1 vccd1 vccd1 _05164_ sky130_fd_sc_hd__a31o_1
XANTENNA__13831__CLK clknet_leaf_59_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11290_ net643 _05984_ _05987_ vssd1 vssd1 vccd1 vccd1 _05988_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout794_X net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10241_ final_design.uart.BAUD_counter\[15\] _05113_ vssd1 vssd1 vccd1 vccd1 _05114_
+ sky130_fd_sc_hd__and2_1
XANTENNA__10553__A1_N net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10172_ _05061_ _05063_ final_design.h_out vssd1 vssd1 vccd1 vccd1 final_design.vga.h_next_state\[0\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_63_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout961_X net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13981__CLK clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1104 net1105 vssd1 vssd1 vccd1 vccd1 net1104 sky130_fd_sc_hd__clkbuf_2
XANTENNA__11765__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1115 net1116 vssd1 vssd1 vccd1 vccd1 net1115 sky130_fd_sc_hd__clkbuf_2
Xfanout1126 net1127 vssd1 vssd1 vccd1 vccd1 net1126 sky130_fd_sc_hd__clkbuf_2
Xfanout1137 net1139 vssd1 vssd1 vccd1 vccd1 net1137 sky130_fd_sc_hd__clkbuf_4
Xfanout1148 net1149 vssd1 vssd1 vccd1 vccd1 net1148 sky130_fd_sc_hd__clkbuf_2
Xfanout1159 net1162 vssd1 vssd1 vccd1 vccd1 net1159 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07544__A net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13931_ clknet_leaf_53_clk _01162_ net1185 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[919\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout183 _06067_ vssd1 vssd1 vccd1 vccd1 net183 sky130_fd_sc_hd__clkbuf_2
Xfanout194 net195 vssd1 vssd1 vccd1 vccd1 net194 sky130_fd_sc_hd__buf_2
XANTENNA__11700__B1 net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13862_ clknet_leaf_52_clk _01093_ net1175 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[850\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_44_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12256__A1 net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12813_ net1346 vssd1 vssd1 vccd1 vccd1 _00254_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_69_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13793_ clknet_leaf_47_clk _01024_ net1203 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[781\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_74_1582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_2922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12744_ _05059_ _06373_ net954 vssd1 vssd1 vccd1 vccd1 _06383_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_80_2944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13361__CLK clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12893__Q final_design.data_from_mem\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12675_ final_design.VGA_data_control.ready_data\[25\] net1019 net974 final_design.data_from_mem\[25\]
+ vssd1 vssd1 vccd1 vccd1 _06325_ sky130_fd_sc_hd__a22o_1
XFILLER_0_38_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_1891 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12929__CLK clknet_leaf_47_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12559__A2 net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11626_ net425 net560 _06170_ net298 net1469 vssd1 vssd1 vccd1 vccd1 _00445_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_13_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11231__A2 net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11557_ net556 net420 _06134_ net302 net1617 vssd1 vssd1 vccd1 vccd1 _00412_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_78_2862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_2873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_2884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_2726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10508_ final_design.CPU_instr_adr\[2\] net1057 final_design.CPU_instr_adr\[3\] vssd1
+ vssd1 vccd1 vccd1 _05257_ sky130_fd_sc_hd__a21oi_1
Xhold609 final_design.cpu.reg_window\[891\] vssd1 vssd1 vccd1 vccd1 net1951 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_55_2103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_2737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11488_ net185 _06093_ vssd1 vssd1 vccd1 vccd1 _06112_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_74_2748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10439_ net1457 net1027 _05203_ net245 vssd1 vssd1 vccd1 vccd1 _00160_ sky130_fd_sc_hd__a22o_1
X_13227_ clknet_leaf_53_clk _00458_ net1187 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[215\]
+ sky130_fd_sc_hd__dfrtp_1
X_13158_ clknet_leaf_50_clk _00389_ net1168 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[146\]
+ sky130_fd_sc_hd__dfrtp_1
X_12109_ net1680 net208 net388 vssd1 vssd1 vccd1 vccd1 _00833_ sky130_fd_sc_hd__mux2_1
X_13089_ clknet_leaf_47_clk _00320_ net1198 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[77\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08148__C1 net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_2519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11298__A2 _05994_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07650_ net719 _02600_ net877 vssd1 vssd1 vccd1 vccd1 _02601_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_36_1319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06601_ _01548_ _01549_ _01550_ _01551_ net776 net794 vssd1 vssd1 vccd1 vccd1 _01552_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__12247__A1 net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13704__CLK clknet_leaf_40_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07581_ _02528_ _02529_ _02530_ _02531_ net685 net706 vssd1 vssd1 vccd1 vccd1 _02532_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_57_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09320_ net460 _03639_ vssd1 vssd1 vccd1 vccd1 _04239_ sky130_fd_sc_hd__nor2_1
X_06532_ _01478_ _01479_ _01457_ _01459_ vssd1 vssd1 vccd1 vccd1 _01483_ sky130_fd_sc_hd__a211o_1
XFILLER_0_38_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09663__A2 _04581_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09251_ _02673_ _02705_ _04168_ _04169_ vssd1 vssd1 vccd1 vccd1 _04170_ sky130_fd_sc_hd__o31a_1
X_06463_ _01405_ _01412_ _00211_ vssd1 vssd1 vccd1 vccd1 _01414_ sky130_fd_sc_hd__a21o_2
X_08202_ net707 _03152_ vssd1 vssd1 vccd1 vccd1 _03153_ sky130_fd_sc_hd__nor2_1
XANTENNA__13854__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09182_ _04097_ _04099_ vssd1 vssd1 vccd1 vccd1 _04101_ sky130_fd_sc_hd__nor2_1
XANTENNA__13009__RESET_B net1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11758__A0 net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08133_ net713 _03077_ net723 vssd1 vssd1 vccd1 vccd1 _03084_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_50_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10754__S net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12094__X _06265_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09820__C1 net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout218_A net219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08064_ _03011_ _03012_ _03013_ _03014_ net682 net702 vssd1 vssd1 vccd1 vccd1 _03015_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__08224__S net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10981__A1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07015_ _01953_ _01954_ _01965_ net881 vssd1 vssd1 vccd1 vccd1 _01966_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_25_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1127_A net1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout587_A _05868_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13234__CLK clknet_leaf_39_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08966_ net2513 net1038 _03904_ vssd1 vssd1 vccd1 vccd1 _00230_ sky130_fd_sc_hd__o21a_1
X_07917_ _02866_ _02867_ vssd1 vssd1 vccd1 vccd1 _02868_ sky130_fd_sc_hd__or2_2
X_08897_ final_design.CPU_instr_adr\[26\] _03798_ vssd1 vssd1 vccd1 vccd1 _03843_
+ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout375_X net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout754_A net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08179__B net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07848_ net606 _02797_ _02773_ vssd1 vssd1 vccd1 vccd1 _02799_ sky130_fd_sc_hd__o21a_1
XANTENNA__07651__X _02602_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13384__CLK clknet_leaf_41_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout921_A net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout542_X net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07779_ _02724_ _02729_ net711 vssd1 vssd1 vccd1 vccd1 _02730_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09518_ _04204_ _04336_ net472 vssd1 vssd1 vccd1 vccd1 _04437_ sky130_fd_sc_hd__mux2_1
X_10790_ _05508_ _05524_ net1005 vssd1 vssd1 vccd1 vccd1 _05526_ sky130_fd_sc_hd__a21o_1
XANTENNA__12429__B net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11997__B1 net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09449_ _04296_ _04364_ net473 vssd1 vssd1 vccd1 vccd1 _04368_ sky130_fd_sc_hd__mux2_2
X_12460_ net2214 net183 net336 vssd1 vssd1 vccd1 vccd1 _01167_ sky130_fd_sc_hd__mux2_1
XANTENNA__11749__A0 net209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08923__A net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11411_ net2157 net228 net311 vssd1 vssd1 vccd1 vccd1 _00308_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_1873 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12391_ net1675 net185 net270 vssd1 vssd1 vccd1 vccd1 _01102_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14130_ clknet_leaf_20_clk final_design.vga.v_next_state\[1\] net1159 vssd1 vssd1
+ vccd1 vccd1 final_design.vga.v_current_state\[1\] sky130_fd_sc_hd__dfrtp_1
X_11342_ net663 _03857_ net737 vssd1 vssd1 vccd1 vccd1 _06033_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_34_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08134__S net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14061_ clknet_leaf_15_clk _00023_ net1091 vssd1 vssd1 vccd1 vccd1 final_design.uart.BAUD_counter\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_11273_ net646 net205 vssd1 vssd1 vccd1 vccd1 _05973_ sky130_fd_sc_hd__and2_1
XFILLER_0_82_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input50_A mem_adr_start[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10224_ _05103_ net800 _05102_ vssd1 vssd1 vccd1 vccd1 _00036_ sky130_fd_sc_hd__and3b_1
X_13012_ clknet_leaf_12_clk _00243_ net1090 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11495__S net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10155_ _05045_ _05051_ _05052_ vssd1 vssd1 vccd1 vccd1 final_design.vga.h_next_count\[3\]
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_7_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12888__Q final_design.data_from_mem\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10086_ _01369_ _01397_ _01398_ _05001_ vssd1 vssd1 vccd1 vccd1 _05002_ sky130_fd_sc_hd__and4_1
Xhold6 final_design.cpu.reg_window\[13\] vssd1 vssd1 vccd1 vccd1 net1348 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13727__CLK clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10412__B _05181_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13914_ clknet_leaf_63_clk _01145_ net1122 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[902\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13845_ clknet_leaf_57_clk _01076_ net1145 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[833\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_71_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08528__S0 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13877__CLK clknet_leaf_56_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13776_ clknet_leaf_34_clk _01007_ net1236 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[764\]
+ sky130_fd_sc_hd__dfrtp_1
X_10988_ _04529_ net252 vssd1 vssd1 vccd1 vccd1 _05714_ sky130_fd_sc_hd__nor2_1
XANTENNA__06618__A net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11988__B1 net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12727_ final_design.VGA_data_control.v_count\[1\] _06361_ _06363_ _06367_ vssd1
+ vssd1 vccd1 vccd1 _06368_ sky130_fd_sc_hd__a31o_1
XANTENNA__07656__A1 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12658_ _06316_ net1450 net979 vssd1 vssd1 vccd1 vccd1 _01331_ sky130_fd_sc_hd__mux2_1
XANTENNA__13107__CLK clknet_leaf_36_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07408__A1 final_design.data_from_mem\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10574__S net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11609_ net242 net631 vssd1 vssd1 vccd1 vccd1 _06162_ sky130_fd_sc_hd__and2_1
X_12589_ net1531 net997 net983 final_design.data_from_mem\[7\] vssd1 vssd1 vccd1 vccd1
+ _01282_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_10_clk clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_10_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_20_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08081__B2 _01850_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold406 final_design.cpu.reg_window\[248\] vssd1 vssd1 vccd1 vccd1 net1748 sky130_fd_sc_hd__dlygate4sd3_1
Xhold417 final_design.cpu.reg_window\[979\] vssd1 vssd1 vccd1 vccd1 net1759 sky130_fd_sc_hd__dlygate4sd3_1
Xhold428 final_design.cpu.reg_window\[977\] vssd1 vssd1 vccd1 vccd1 net1770 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold439 final_design.cpu.reg_window\[964\] vssd1 vssd1 vccd1 vccd1 net1781 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13257__CLK clknet_leaf_36_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10715__A1 net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout908 net909 vssd1 vssd1 vccd1 vccd1 net908 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10715__B2 net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout919 net922 vssd1 vssd1 vccd1 vccd1 net919 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_42_1356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08820_ _03768_ _03769_ _03668_ vssd1 vssd1 vccd1 vccd1 _03771_ sky130_fd_sc_hd__o21bai_1
Xhold1106 final_design.cpu.reg_window\[612\] vssd1 vssd1 vccd1 vccd1 net2448 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1117 final_design.cpu.reg_window\[149\] vssd1 vssd1 vccd1 vccd1 net2459 sky130_fd_sc_hd__dlygate4sd3_1
X_08751_ _03700_ _03701_ vssd1 vssd1 vccd1 vccd1 _03702_ sky130_fd_sc_hd__and2_1
Xhold1128 final_design.cpu.reg_window\[380\] vssd1 vssd1 vccd1 vccd1 net2470 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1139 final_design.cpu.reg_window\[317\] vssd1 vssd1 vccd1 vccd1 net2481 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_75_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07702_ final_design.cpu.reg_window\[155\] final_design.cpu.reg_window\[187\] net867
+ vssd1 vssd1 vccd1 vccd1 _02653_ sky130_fd_sc_hd__mux2_1
X_08682_ _03611_ _03630_ _03628_ _03612_ vssd1 vssd1 vccd1 vccd1 _03633_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__07344__A0 final_design.data_from_mem\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07633_ final_design.cpu.reg_window\[92\] final_design.cpu.reg_window\[124\] net860
+ vssd1 vssd1 vccd1 vccd1 _02584_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_0_169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07564_ _02504_ net602 vssd1 vssd1 vccd1 vccd1 _02515_ sky130_fd_sc_hd__nand2_1
XANTENNA__08219__S net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11979__B1 net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07123__S net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06515_ final_design.data_from_mem\[3\] net1041 net993 net990 vssd1 vssd1 vccd1 vccd1
+ _01466_ sky130_fd_sc_hd__and4_1
X_09303_ net594 _04219_ vssd1 vssd1 vccd1 vccd1 _04222_ sky130_fd_sc_hd__nand2_4
XTAP_TAPCELL_ROW_17_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07495_ _02130_ _02159_ _02443_ _02129_ _02099_ vssd1 vssd1 vccd1 vccd1 _02446_ sky130_fd_sc_hd__o311a_1
XFILLER_0_76_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout335_A net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06446_ final_design.VGA_data_control.v_count\[7\] final_design.VGA_data_control.v_count\[8\]
+ final_design.VGA_data_control.v_count\[5\] final_design.VGA_data_control.v_count\[6\]
+ vssd1 vssd1 vccd1 vccd1 _01400_ sky130_fd_sc_hd__or4_2
XPHY_EDGE_ROW_3_Right_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09234_ _03390_ _03423_ _04148_ _04152_ vssd1 vssd1 vccd1 vccd1 _04153_ sky130_fd_sc_hd__a31o_2
XFILLER_0_61_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06962__S net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14032__CLK clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09165_ net496 net492 vssd1 vssd1 vccd1 vccd1 _04084_ sky130_fd_sc_hd__nor2_1
XFILLER_0_66_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout502_A net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1244_A net1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08116_ net611 _03065_ _03066_ net539 vssd1 vssd1 vccd1 vccd1 _03067_ sky130_fd_sc_hd__a211oi_1
XTAP_TAPCELL_ROW_40_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_1857 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09096_ _02332_ _02431_ net622 vssd1 vssd1 vccd1 vccd1 _04019_ sky130_fd_sc_hd__o21a_1
XFILLER_0_47_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08047_ _01881_ net602 vssd1 vssd1 vccd1 vccd1 _02998_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout1032_X net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14182__CLK clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12156__A0 net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold940 final_design.cpu.reg_window\[643\] vssd1 vssd1 vccd1 vccd1 net2282 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_47_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_1570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold951 final_design.cpu.reg_window\[389\] vssd1 vssd1 vccd1 vccd1 net2293 sky130_fd_sc_hd__dlygate4sd3_1
Xhold962 final_design.cpu.reg_window\[558\] vssd1 vssd1 vccd1 vccd1 net2304 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07258__S0 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold973 final_design.cpu.reg_window\[296\] vssd1 vssd1 vccd1 vccd1 net2315 sky130_fd_sc_hd__dlygate4sd3_1
Xhold984 final_design.cpu.reg_window\[826\] vssd1 vssd1 vccd1 vccd1 net2326 sky130_fd_sc_hd__dlygate4sd3_1
Xhold995 final_design.CPU_instr_adr\[7\] vssd1 vssd1 vccd1 vccd1 net2337 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout871_A net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout969_A net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10072__X _04990_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11609__A net242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10513__A net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09998_ net451 _04907_ _04916_ vssd1 vssd1 vccd1 vccd1 _04917_ sky130_fd_sc_hd__a21o_1
XANTENNA__06710__B _01660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08949_ _01825_ _02460_ net621 vssd1 vssd1 vccd1 vccd1 _03889_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout757_X net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11960_ _06162_ net282 net405 net2010 vssd1 vssd1 vccd1 vccd1 _00693_ sky130_fd_sc_hd__a22o_1
XFILLER_0_73_1817 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07822__A _01788_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10911_ _05639_ _05640_ net963 vssd1 vssd1 vccd1 vccd1 _05641_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07430__S0 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11891_ net238 net2070 net272 vssd1 vssd1 vccd1 vccd1 _00633_ sky130_fd_sc_hd__mux2_1
X_13630_ clknet_leaf_12_clk _00861_ net1087 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[618\]
+ sky130_fd_sc_hd__dfrtp_1
X_10842_ net962 _05574_ vssd1 vssd1 vccd1 vccd1 _05575_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_15_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07033__S net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12789__20 clknet_leaf_30_clk vssd1 vssd1 vccd1 vccd1 net1330 sky130_fd_sc_hd__inv_2
X_13561_ clknet_leaf_54_clk _00792_ net1177 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[549\]
+ sky130_fd_sc_hd__dfrtp_1
X_10773_ net253 _04697_ vssd1 vssd1 vccd1 vccd1 _05509_ sky130_fd_sc_hd__and2b_1
XANTENNA__12631__B2 final_design.data_from_mem\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07733__S1 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12512_ _06174_ net344 net326 net1593 vssd1 vssd1 vccd1 vccd1 _01217_ sky130_fd_sc_hd__a22o_1
XANTENNA_input98_A memory_size[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13492_ clknet_leaf_10_clk _00723_ net1102 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[480\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_246 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12443_ net2364 net214 net334 vssd1 vssd1 vccd1 vccd1 _01150_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_1867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11198__A1 final_design.reqhand.data_from_UART\[7\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_1_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1889 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12374_ net1716 net217 net268 vssd1 vssd1 vccd1 vccd1 _01085_ sky130_fd_sc_hd__mux2_1
XANTENNA__10945__A1 _05508_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14113_ clknet_leaf_14_clk net2529 net1103 vssd1 vssd1 vccd1 vccd1 final_design.reqhand.data_from_UART\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_11325_ net434 net579 _06018_ net316 net2188 vssd1 vssd1 vccd1 vccd1 _00296_ sky130_fd_sc_hd__a32o_1
XFILLER_0_82_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14044_ clknet_leaf_16_clk _00036_ net1094 vssd1 vssd1 vccd1 vccd1 final_design.uart.BAUD_counter\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_11256_ _04631_ net658 _05843_ _05957_ vssd1 vssd1 vccd1 vccd1 _05958_ sky130_fd_sc_hd__a211oi_1
X_10207_ final_design.uart.BAUD_counter\[1\] final_design.uart.BAUD_counter\[0\] final_design.uart.BAUD_counter\[2\]
+ vssd1 vssd1 vccd1 vccd1 _05093_ sky130_fd_sc_hd__and3_1
XANTENNA__12114__S net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11187_ _04863_ net655 _05843_ _05896_ vssd1 vssd1 vccd1 vccd1 _05897_ sky130_fd_sc_hd__a211oi_2
XANTENNA__10423__A _03065_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06620__B _01570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10138_ _01389_ final_design.vga.h_current_state\[1\] _05009_ vssd1 vssd1 vccd1 vccd1
+ _05040_ sky130_fd_sc_hd__and3_1
XANTENNA__11238__B net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_59_clk clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_59_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__09315__A1 _04233_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08118__A2 _03065_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10069_ _04987_ vssd1 vssd1 vccd1 vccd1 _04988_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_1403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_1327 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13828_ clknet_leaf_51_clk _01059_ net1171 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[816\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_8_1857 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1892 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14055__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13759_ clknet_leaf_8_clk _00990_ net1154 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[747\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07280_ final_design.cpu.reg_window\[902\] final_design.cpu.reg_window\[934\] net903
+ vssd1 vssd1 vccd1 vccd1 _02231_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11701__B net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11189__A1 net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10399__A1_N net250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07179__A _02127_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_3_clk_X clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold203 final_design.cpu.reg_window\[708\] vssd1 vssd1 vccd1 vccd1 net1545 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold214 final_design.cpu.reg_window\[677\] vssd1 vssd1 vccd1 vccd1 net1556 sky130_fd_sc_hd__dlygate4sd3_1
Xhold225 final_design.cpu.reg_window\[897\] vssd1 vssd1 vccd1 vccd1 net1567 sky130_fd_sc_hd__dlygate4sd3_1
Xhold236 final_design.reqhand.instruction\[27\] vssd1 vssd1 vccd1 vccd1 net1578 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12138__A0 net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold247 final_design.cpu.reg_window\[80\] vssd1 vssd1 vccd1 vccd1 net1589 sky130_fd_sc_hd__dlygate4sd3_1
Xhold258 final_design.cpu.reg_window\[238\] vssd1 vssd1 vccd1 vccd1 net1600 sky130_fd_sc_hd__dlygate4sd3_1
Xhold269 net136 vssd1 vssd1 vccd1 vccd1 net1611 sky130_fd_sc_hd__dlygate4sd3_1
X_09921_ _04643_ _04839_ net481 vssd1 vssd1 vccd1 vccd1 _04840_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkload22_A clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout705 net706 vssd1 vssd1 vccd1 vccd1 net705 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09554__A1 net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout716 net718 vssd1 vssd1 vccd1 vccd1 net716 sky130_fd_sc_hd__clkbuf_4
Xfanout727 _01493_ vssd1 vssd1 vccd1 vccd1 net727 sky130_fd_sc_hd__clkbuf_4
X_09852_ _04153_ _04154_ _03293_ vssd1 vssd1 vccd1 vccd1 _04771_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07626__B net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout738 net739 vssd1 vssd1 vccd1 vccd1 net738 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11361__A1 _01630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout749 net751 vssd1 vssd1 vccd1 vccd1 net749 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11361__B2 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08803_ final_design.CPU_instr_adr\[23\] _01722_ vssd1 vssd1 vccd1 vccd1 _03754_
+ sky130_fd_sc_hd__nor2_1
X_09783_ _04697_ _04699_ vssd1 vssd1 vccd1 vccd1 _04702_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_52_1972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06995_ final_design.cpu.reg_window\[399\] final_design.cpu.reg_window\[431\] net891
+ vssd1 vssd1 vccd1 vccd1 _01946_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_52_1983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout285_A net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_52_1994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08734_ final_design.CPU_instr_adr\[13\] _02030_ vssd1 vssd1 vccd1 vccd1 _03685_
+ sky130_fd_sc_hd__nand2_1
XANTENNA__09857__A2 net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08665_ _01999_ _02028_ vssd1 vssd1 vccd1 vccd1 _03616_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout452_A net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1194_A net1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06529__Y _01480_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07616_ final_design.cpu.reg_window\[925\] final_design.cpu.reg_window\[957\] net870
+ vssd1 vssd1 vccd1 vccd1 _02567_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13024__RESET_B net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08596_ _03543_ _03544_ _03545_ _03546_ net678 net691 vssd1 vssd1 vccd1 vccd1 _03547_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_27_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout240_X net240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07547_ final_design.cpu.reg_window\[607\] final_design.cpu.reg_window\[639\] net937
+ vssd1 vssd1 vccd1 vccd1 _02498_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_27_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12613__B2 final_design.data_from_mem\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout338_X net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout717_A net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13422__CLK clknet_leaf_42_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10624__B1 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07715__S1 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09569__A net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07478_ _02426_ _02427_ _02395_ vssd1 vssd1 vccd1 vccd1 _02429_ sky130_fd_sc_hd__o21a_1
XANTENNA__11611__B net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09217_ _03070_ _03101_ _03134_ _03164_ vssd1 vssd1 vccd1 vccd1 _04136_ sky130_fd_sc_hd__and4_1
X_06429_ final_design.VGA_data_control.h_count\[3\] vssd1 vssd1 vccd1 vccd1 _01384_
+ sky130_fd_sc_hd__inv_2
XANTENNA_fanout505_X net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11103__S net1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09148_ _04059_ _04066_ net491 vssd1 vssd1 vccd1 vccd1 _04067_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13572__CLK clknet_leaf_54_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09079_ net2538 net1013 _04004_ vssd1 vssd1 vccd1 vccd1 _00217_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_9_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11110_ net1052 _05078_ _05088_ vssd1 vssd1 vccd1 vccd1 _05830_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_9_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07817__A _01657_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12090_ net586 _06068_ net513 net394 net2232 vssd1 vssd1 vccd1 vccd1 _00815_ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout874_X net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold770 final_design.cpu.reg_window\[781\] vssd1 vssd1 vccd1 vccd1 net2112 sky130_fd_sc_hd__dlygate4sd3_1
Xhold781 final_design.cpu.reg_window\[193\] vssd1 vssd1 vccd1 vccd1 net2123 sky130_fd_sc_hd__dlygate4sd3_1
X_11041_ _05764_ _05760_ vssd1 vssd1 vccd1 vccd1 _05765_ sky130_fd_sc_hd__and2b_1
Xhold792 final_design.cpu.reg_window\[337\] vssd1 vssd1 vccd1 vccd1 net2134 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06440__B net34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11352__A1 final_design.data_from_mem\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1761 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11104__A1 net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12992_ net1323 _00223_ net1193 vssd1 vssd1 vccd1 vccd1 final_design.CPU_instr_adr\[12\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__10897__B net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11104__B2 net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08505__C1 _02326_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14078__CLK clknet_leaf_19_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input13_A DAT_I[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11943_ _06144_ net280 net409 net1963 vssd1 vssd1 vccd1 vccd1 _00678_ sky130_fd_sc_hd__a22o_1
XANTENNA__07403__S0 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11874_ _06110_ net293 net520 net2171 vssd1 vssd1 vccd1 vccd1 _00619_ sky130_fd_sc_hd__a22o_1
X_13613_ clknet_leaf_48_clk _00844_ net1185 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[601\]
+ sky130_fd_sc_hd__dfrtp_1
X_10825_ net45 _05558_ vssd1 vssd1 vccd1 vccd1 _05559_ sky130_fd_sc_hd__and2_1
XANTENNA__11407__A2 net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12604__B2 final_design.data_from_mem\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13544_ clknet_leaf_41_clk _00775_ net1219 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[532\]
+ sky130_fd_sc_hd__dfrtp_1
X_10756_ net965 _05492_ vssd1 vssd1 vccd1 vccd1 _05493_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_1620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13915__CLK clknet_leaf_65_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13475_ clknet_leaf_1_clk _00706_ net1071 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[463\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12109__S net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10687_ net70 final_design.VGA_adr\[9\] _05426_ vssd1 vssd1 vccd1 vccd1 _05427_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_10_1653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12426_ _06113_ net357 net340 net2320 vssd1 vssd1 vccd1 vccd1 _01135_ sky130_fd_sc_hd__a22o_1
XFILLER_0_22_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08131__S1 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12357_ net2326 net363 net356 _06053_ vssd1 vssd1 vccd1 vccd1 _01069_ sky130_fd_sc_hd__a22o_1
X_11308_ net647 net564 net200 vssd1 vssd1 vccd1 vccd1 _06004_ sky130_fd_sc_hd__and3_1
X_12288_ net582 _06218_ net514 net370 net1778 vssd1 vssd1 vccd1 vccd1 _01003_ sky130_fd_sc_hd__a32o_1
XANTENNA__06631__A net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08339__A2 _03287_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14027_ clknet_leaf_53_clk _01258_ net1188 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[1015\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11249__A net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11239_ net2456 net315 _05942_ net429 vssd1 vssd1 vccd1 vccd1 _00286_ sky130_fd_sc_hd__a22o_1
XANTENNA__12540__B1 net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13535__RESET_B net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11536__X _06123_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06780_ net752 _01730_ vssd1 vssd1 vccd1 vccd1 _01731_ sky130_fd_sc_hd__nor2_1
XANTENNA__06770__A1 final_design.data_from_mem\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11646__A2 net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_828 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_19_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13445__CLK clknet_leaf_48_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08450_ _03397_ _03398_ _03399_ _03400_ net677 net698 vssd1 vssd1 vccd1 vccd1 _03401_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_19_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08246__A_N net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1889 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07401_ final_design.cpu.reg_window\[578\] final_design.cpu.reg_window\[610\] net913
+ vssd1 vssd1 vccd1 vccd1 _02352_ sky130_fd_sc_hd__mux2_1
X_08381_ final_design.cpu.reg_window\[262\] final_design.cpu.reg_window\[294\] net831
+ vssd1 vssd1 vccd1 vccd1 _03332_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07332_ final_design.cpu.reg_window\[836\] final_design.cpu.reg_window\[868\] net900
+ vssd1 vssd1 vccd1 vccd1 _02283_ sky130_fd_sc_hd__mux2_1
XANTENNA__08275__A1 net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07078__A2 net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08293__A net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06806__A net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07401__S net913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07263_ net533 _02212_ vssd1 vssd1 vccd1 vccd1 _02214_ sky130_fd_sc_hd__nand2_1
XFILLER_0_45_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06525__B _01468_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12359__B1 net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09002_ final_design.CPU_instr_adr\[15\] net1016 _03931_ _03936_ vssd1 vssd1 vccd1
+ vccd1 _00226_ sky130_fd_sc_hd__a22o_1
XFILLER_0_2_1297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07194_ final_design.cpu.reg_window\[969\] final_design.cpu.reg_window\[1001\] net891
+ vssd1 vssd1 vccd1 vccd1 _02145_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_1805 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout200_A _06003_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10385__A2 net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08232__S net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout502 net504 vssd1 vssd1 vccd1 vccd1 net502 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_35_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09904_ _04565_ _04822_ net494 vssd1 vssd1 vccd1 vccd1 _04823_ sky130_fd_sc_hd__a21oi_2
Xfanout513 net515 vssd1 vssd1 vccd1 vccd1 net513 sky130_fd_sc_hd__clkbuf_2
Xfanout524 _06119_ vssd1 vssd1 vccd1 vccd1 net524 sky130_fd_sc_hd__buf_6
XANTENNA__11334__A1 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07538__B1 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1207_A net1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout535 net536 vssd1 vssd1 vccd1 vccd1 net535 sky130_fd_sc_hd__buf_2
XANTENNA__12531__B1 net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout546 _01880_ vssd1 vssd1 vccd1 vccd1 net546 sky130_fd_sc_hd__buf_2
XANTENNA_input5_A DAT_I[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout557 net562 vssd1 vssd1 vccd1 vccd1 net557 sky130_fd_sc_hd__dlymetal6s2s_1
X_09835_ net481 _04442_ _04515_ net318 vssd1 vssd1 vccd1 vccd1 _04754_ sky130_fd_sc_hd__a211o_1
Xfanout568 net571 vssd1 vssd1 vccd1 vccd1 net568 sky130_fd_sc_hd__buf_4
Xfanout579 net580 vssd1 vssd1 vccd1 vccd1 net579 sky130_fd_sc_hd__buf_2
XANTENNA_fanout667_A _01498_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout288_X net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1901 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06687__S net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1008 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09766_ net476 _04055_ _04397_ vssd1 vssd1 vccd1 vccd1 _04685_ sky130_fd_sc_hd__or3_1
X_06978_ _01925_ _01926_ _01927_ _01928_ net773 net791 vssd1 vssd1 vccd1 vccd1 _01929_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__09063__S net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11098__B1 _04990_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08717_ _01361_ _01690_ vssd1 vssd1 vccd1 vccd1 _03668_ sky130_fd_sc_hd__nor2_1
XANTENNA__08189__S1 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11165__Y _05877_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11606__B net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09697_ net729 _04613_ _04615_ vssd1 vssd1 vccd1 vccd1 _04616_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_1_242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout834_A net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout455_X net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1197_X net1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08502__A2 _03450_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09160__C1 _01627_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08648_ _02769_ _03597_ _03598_ vssd1 vssd1 vccd1 vccd1 _03599_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_48_1849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09138__S0 net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13938__CLK clknet_leaf_44_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout622_X net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08579_ final_design.cpu.reg_window\[64\] final_design.cpu.reg_window\[96\] net814
+ vssd1 vssd1 vccd1 vccd1 _03530_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10610_ _05334_ _05337_ _05353_ vssd1 vssd1 vccd1 vccd1 _05354_ sky130_fd_sc_hd__o21ai_2
XANTENNA__09299__A _02503_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11590_ net187 net636 vssd1 vssd1 vccd1 vccd1 _06151_ sky130_fd_sc_hd__and2_1
XFILLER_0_0_1905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10541_ net95 final_design.VGA_adr\[3\] vssd1 vssd1 vccd1 vccd1 _05288_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13260_ clknet_leaf_46_clk _00491_ net1214 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[248\]
+ sky130_fd_sc_hd__dfrtp_1
X_10472_ net726 _04805_ net250 _04990_ vssd1 vssd1 vccd1 vccd1 _05223_ sky130_fd_sc_hd__o31ai_2
XFILLER_0_66_1440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12211_ net559 _06139_ net504 net376 net1631 vssd1 vssd1 vccd1 vccd1 _00929_ sky130_fd_sc_hd__a32o_1
X_13191_ clknet_leaf_62_clk _00422_ net1123 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[179\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_62_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10376__A2 net1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13318__CLK clknet_leaf_51_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12142_ net212 net2482 net384 vssd1 vssd1 vccd1 vccd1 _00863_ sky130_fd_sc_hd__mux2_1
XANTENNA__08142__S net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12073_ net2492 net393 net498 _05942_ vssd1 vssd1 vccd1 vccd1 _00798_ sky130_fd_sc_hd__a22o_1
XANTENNA__11325__A1 net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12522__B1 net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11024_ _05747_ _05748_ vssd1 vssd1 vccd1 vccd1 _05749_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_70_2581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_2592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11876__A2 net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11356__X _06046_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13468__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07553__Y _02504_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12975_ clknet_leaf_20_clk _00000_ net1160 vssd1 vssd1 vccd1 vccd1 final_design.reqhand.current_client\[0\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__11628__A2 net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12999__RESET_B net1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11926_ net555 net240 net634 vssd1 vssd1 vccd1 vccd1 _06253_ sky130_fd_sc_hd__and3_1
XFILLER_0_73_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1805 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11857_ net2554 net517 _06240_ net429 vssd1 vssd1 vccd1 vccd1 _00606_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_64_2385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_1849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_2396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12589__B1 net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10808_ _05508_ _05542_ vssd1 vssd1 vccd1 vccd1 _05543_ sky130_fd_sc_hd__or2_1
XANTENNA__09454__A0 _04300_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_2249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11788_ net647 net555 net207 vssd1 vssd1 vccd1 vccd1 _06233_ sky130_fd_sc_hd__and3_1
X_13527_ clknet_leaf_4_clk _00758_ net1083 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[515\]
+ sky130_fd_sc_hd__dfrtp_1
X_10739_ net41 _05476_ vssd1 vssd1 vccd1 vccd1 _05477_ sky130_fd_sc_hd__and2_1
XANTENNA__11800__A2 net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09496__X _04415_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13458_ clknet_leaf_38_clk _00689_ net1189 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[446\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_11_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09757__A1 net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12409_ _06241_ net499 net338 net2213 vssd1 vssd1 vccd1 vccd1 _01119_ sky130_fd_sc_hd__a22o_1
Xoutput105 net105 vssd1 vssd1 vccd1 vccd1 ADR_O[13] sky130_fd_sc_hd__clkbuf_4
X_13389_ clknet_leaf_44_clk _00620_ net1205 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[377\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_2178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput116 net116 vssd1 vssd1 vccd1 vccd1 ADR_O[23] sky130_fd_sc_hd__clkbuf_4
XANTENNA__10367__A2 net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07768__B1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_2189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput127 net127 vssd1 vssd1 vccd1 vccd1 ADR_O[4] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_11_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput138 net138 vssd1 vssd1 vccd1 vccd1 DAT_O[13] sky130_fd_sc_hd__buf_2
Xoutput149 net149 vssd1 vssd1 vccd1 vccd1 DAT_O[23] sky130_fd_sc_hd__buf_2
XFILLER_0_11_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07950_ _02866_ _02867_ _02897_ _02899_ vssd1 vssd1 vccd1 vccd1 _02901_ sky130_fd_sc_hd__o22a_1
XANTENNA__12513__B1 net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06901_ _01468_ net736 net744 vssd1 vssd1 vccd1 vccd1 _01852_ sky130_fd_sc_hd__a21o_1
XANTENNA__11867__A2 net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07881_ net605 _02830_ _02805_ vssd1 vssd1 vccd1 vccd1 _02832_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_78_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09620_ _04100_ _04491_ net486 vssd1 vssd1 vccd1 vccd1 _04539_ sky130_fd_sc_hd__mux2_1
X_06832_ net762 _01782_ vssd1 vssd1 vccd1 vccd1 _01783_ sky130_fd_sc_hd__or2_1
XANTENNA__12302__S net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12835__CLK clknet_leaf_19_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09551_ _02964_ _04046_ _04351_ _04456_ _04469_ vssd1 vssd1 vccd1 vccd1 _04470_ sky130_fd_sc_hd__a41o_1
X_06763_ final_design.cpu.reg_window\[535\] final_design.cpu.reg_window\[567\] net928
+ vssd1 vssd1 vccd1 vccd1 _01714_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_1642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08502_ net608 _03450_ _03451_ vssd1 vssd1 vccd1 vccd1 _03453_ sky130_fd_sc_hd__a21oi_2
XANTENNA__09142__C1 _02422_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06694_ final_design.cpu.reg_window\[857\] final_design.cpu.reg_window\[889\] net933
+ vssd1 vssd1 vccd1 vccd1 _01645_ sky130_fd_sc_hd__mux2_1
X_09482_ net549 net548 net546 net545 net459 net469 vssd1 vssd1 vccd1 vccd1 _04401_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_56_1697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08433_ _03371_ _03372_ _03383_ net876 vssd1 vssd1 vccd1 vccd1 _03384_ sky130_fd_sc_hd__a22oi_4
XFILLER_0_59_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout248_A net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11442__A net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08364_ final_design.cpu.reg_window\[711\] final_design.cpu.reg_window\[743\] net806
+ vssd1 vssd1 vccd1 vccd1 _03315_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07131__S net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11252__B1 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07315_ _02248_ _02254_ _02265_ net883 vssd1 vssd1 vccd1 vccd1 _02266_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_50_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08295_ final_design.cpu.reg_window\[521\] final_design.cpu.reg_window\[553\] net808
+ vssd1 vssd1 vccd1 vccd1 _03246_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout1157_A net1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07246_ final_design.cpu.reg_window\[391\] final_design.cpu.reg_window\[423\] net892
+ vssd1 vssd1 vccd1 vccd1 _02197_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07177_ _01477_ _01505_ net667 vssd1 vssd1 vccd1 vccd1 _02128_ sky130_fd_sc_hd__mux2_2
XFILLER_0_67_1793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10358__A2 net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11555__A1 net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08470__B net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07367__A net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout784_A _01419_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13610__CLK clknet_leaf_60_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout310 _06092_ vssd1 vssd1 vccd1 vccd1 net310 sky130_fd_sc_hd__clkbuf_8
XANTENNA__11307__A1 _04570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12504__B1 net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout321 _04047_ vssd1 vssd1 vccd1 vccd1 net321 sky130_fd_sc_hd__buf_4
Xfanout332 net333 vssd1 vssd1 vccd1 vccd1 net332 sky130_fd_sc_hd__buf_4
Xfanout343 net345 vssd1 vssd1 vccd1 vccd1 net343 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout951_A net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout572_X net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout354 net359 vssd1 vssd1 vccd1 vccd1 net354 sky130_fd_sc_hd__clkbuf_4
Xfanout365 net367 vssd1 vssd1 vccd1 vccd1 net365 sky130_fd_sc_hd__buf_4
Xfanout376 net377 vssd1 vssd1 vccd1 vccd1 net376 sky130_fd_sc_hd__clkbuf_8
Xfanout387 _06266_ vssd1 vssd1 vccd1 vccd1 net387 sky130_fd_sc_hd__clkbuf_8
X_09818_ _04222_ _04726_ _04731_ _04736_ vssd1 vssd1 vccd1 vccd1 _04737_ sky130_fd_sc_hd__o211a_1
Xfanout398 net399 vssd1 vssd1 vccd1 vccd1 net398 sky130_fd_sc_hd__clkbuf_8
XANTENNA__13760__CLK clknet_leaf_11_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09749_ _03195_ net444 net438 _03197_ vssd1 vssd1 vccd1 vccd1 _04668_ sky130_fd_sc_hd__o22a_1
X_12760_ _06339_ _06391_ vssd1 vssd1 vccd1 vccd1 _06396_ sky130_fd_sc_hd__nand2_1
XANTENNA__08487__A1 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11711_ net197 net628 vssd1 vssd1 vccd1 vccd1 _06214_ sky130_fd_sc_hd__and2_1
XFILLER_0_55_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12691_ _01390_ _05039_ net796 net2427 vssd1 vssd1 vccd1 vccd1 _01347_ sky130_fd_sc_hd__a22o_1
XANTENNA__08645__B _03593_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14116__CLK clknet_leaf_15_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11642_ net432 net573 _06178_ net301 net1490 vssd1 vssd1 vccd1 vccd1 _00453_ sky130_fd_sc_hd__a32o_1
XANTENNA__08137__S net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10046__A1 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10046__B2 _04423_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08334__S1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11573_ net575 net424 _06142_ net305 net1707 vssd1 vssd1 vccd1 vccd1 _00420_ sky130_fd_sc_hd__a32o_1
Xinput18 DAT_I[24] vssd1 vssd1 vccd1 vccd1 net18 sky130_fd_sc_hd__clkbuf_1
XANTENNA__07998__B1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input80_A memory_size[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13312_ clknet_leaf_10_clk _00543_ net1101 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[300\]
+ sky130_fd_sc_hd__dfrtp_1
X_10524_ _05235_ _05252_ _05251_ vssd1 vssd1 vccd1 vccd1 _05272_ sky130_fd_sc_hd__o21ai_1
Xinput29 DAT_I[5] vssd1 vssd1 vccd1 vccd1 net29 sky130_fd_sc_hd__clkbuf_2
X_13243_ clknet_leaf_0_clk _00474_ net1062 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[231\]
+ sky130_fd_sc_hd__dfrtp_1
X_10455_ net1516 net1035 _05211_ net248 vssd1 vssd1 vccd1 vccd1 _00168_ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09203__A3 _04119_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_2790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13174_ clknet_leaf_60_clk _00405_ net1138 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[162\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_46_1877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10386_ wb_manage.curr_state\[1\] net1 wb_manage.curr_state\[2\] vssd1 vssd1 vccd1
+ vccd1 _05174_ sky130_fd_sc_hd__or3b_2
XTAP_TAPCELL_ROW_53_2020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output167_A net167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10415__B _05190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_2031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_43_clk_X clknet_leaf_43_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12125_ net1953 net178 net390 vssd1 vssd1 vccd1 vccd1 _00849_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_72_2676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13290__CLK clknet_leaf_59_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06973__A1 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12858__CLK clknet_leaf_18_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12056_ net2439 net180 net398 vssd1 vssd1 vccd1 vccd1 _00784_ sky130_fd_sc_hd__mux2_1
XANTENNA__11849__A2 net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11007_ _05711_ _05732_ _05731_ vssd1 vssd1 vccd1 vccd1 _05733_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12122__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07073__S1 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_58_clk_X clknet_leaf_58_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_2447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_1913 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_2458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12958_ clknet_leaf_30_clk _00196_ net1196 vssd1 vssd1 vccd1 vccd1 net116 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_66_2469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11909_ final_design.cpu.reg_window\[407\] _05845_ vssd1 vssd1 vccd1 vccd1 _06249_
+ sky130_fd_sc_hd__or2_1
X_12889_ clknet_leaf_17_clk _00127_ net1109 vssd1 vssd1 vccd1 vccd1 final_design.data_from_mem\[23\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_16_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07100_ net750 _02050_ vssd1 vssd1 vccd1 vccd1 _02051_ sky130_fd_sc_hd__or2_1
XANTENNA__11785__B2 net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08080_ net547 _03024_ vssd1 vssd1 vccd1 vccd1 _03031_ sky130_fd_sc_hd__nor2_1
XFILLER_0_71_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07031_ net750 _01975_ net745 vssd1 vssd1 vccd1 vccd1 _01982_ sky130_fd_sc_hd__o21a_1
XFILLER_0_2_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13633__CLK clknet_leaf_46_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06803__B _01752_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1917 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08982_ _03918_ vssd1 vssd1 vccd1 vccd1 _03919_ sky130_fd_sc_hd__inv_2
X_07933_ final_design.cpu.reg_window\[982\] final_design.cpu.reg_window\[1014\] net837
+ vssd1 vssd1 vccd1 vccd1 _02884_ sky130_fd_sc_hd__mux2_1
XANTENNA__13783__CLK clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08166__B1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout198_A _06010_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12032__S net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07864_ final_design.cpu.reg_window\[148\] final_design.cpu.reg_window\[180\] net868
+ vssd1 vssd1 vccd1 vccd1 _02815_ sky130_fd_sc_hd__mux2_1
XANTENNA__10512__A2 net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09603_ _02702_ net439 _04519_ _04521_ vssd1 vssd1 vccd1 vccd1 _04522_ sky130_fd_sc_hd__o211a_1
XFILLER_0_39_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06815_ final_design.cpu.reg_window\[341\] final_design.cpu.reg_window\[373\] net938
+ vssd1 vssd1 vccd1 vccd1 _01766_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07795_ final_design.cpu.reg_window\[25\] final_design.cpu.reg_window\[57\] net856
+ vssd1 vssd1 vccd1 vccd1 _02746_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13013__CLK clknet_leaf_56_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout365_A net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14139__CLK clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09534_ net76 _04187_ net77 vssd1 vssd1 vccd1 vccd1 _04453_ sky130_fd_sc_hd__o21ai_1
X_06746_ _01693_ _01694_ _01695_ _01696_ net772 net795 vssd1 vssd1 vccd1 vccd1 _01697_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__11473__A0 net223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09465_ _04382_ _04383_ vssd1 vssd1 vccd1 vccd1 _04384_ sky130_fd_sc_hd__or2_1
X_06677_ final_design.reqhand.instruction\[26\] final_design.data_from_mem\[26\] net973
+ vssd1 vssd1 vccd1 vccd1 _01628_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout532_A _02239_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11172__A net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08416_ final_design.cpu.reg_window\[5\] final_design.cpu.reg_window\[37\] net840
+ vssd1 vssd1 vccd1 vccd1 _03367_ sky130_fd_sc_hd__mux2_1
XANTENNA__09418__A0 _01657_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12017__A2 net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13163__CLK clknet_leaf_38_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09396_ net467 _04104_ vssd1 vssd1 vccd1 vccd1 _04315_ sky130_fd_sc_hd__or2_1
XANTENNA__10028__A1 _04342_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08347_ final_design.cpu.reg_window\[327\] final_design.cpu.reg_window\[359\] net819
+ vssd1 vssd1 vccd1 vccd1 _03298_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout320_X net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout418_X net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07796__S net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08278_ _03227_ _03228_ vssd1 vssd1 vccd1 vccd1 _03229_ sky130_fd_sc_hd__nor2_2
XANTENNA__06553__X _01504_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1719 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07229_ final_design.cpu.reg_window\[968\] final_design.cpu.reg_window\[1000\] net897
+ vssd1 vssd1 vccd1 vccd1 _02180_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10240_ _05113_ net799 _05112_ vssd1 vssd1 vccd1 vccd1 _00011_ sky130_fd_sc_hd__and3b_1
XANTENNA__07827__S0 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout787_X net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10171_ final_design.vga.h_current_state\[0\] final_design.vga.h_current_state\[1\]
+ _05016_ _05062_ vssd1 vssd1 vccd1 vccd1 _05063_ sky130_fd_sc_hd__a31o_1
Xfanout1105 net1116 vssd1 vssd1 vccd1 vccd1 net1105 sky130_fd_sc_hd__buf_2
Xfanout1116 net1117 vssd1 vssd1 vccd1 vccd1 net1116 sky130_fd_sc_hd__clkbuf_2
Xfanout1127 net1167 vssd1 vssd1 vccd1 vccd1 net1127 sky130_fd_sc_hd__buf_2
Xfanout1138 net1139 vssd1 vssd1 vccd1 vccd1 net1138 sky130_fd_sc_hd__clkbuf_4
Xfanout1149 net1150 vssd1 vssd1 vccd1 vccd1 net1149 sky130_fd_sc_hd__buf_2
X_13930_ clknet_leaf_60_clk _01161_ net1142 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[918\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06707__A1 net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout184 _06060_ vssd1 vssd1 vccd1 vccd1 net184 sky130_fd_sc_hd__buf_2
Xfanout195 _06024_ vssd1 vssd1 vccd1 vccd1 net195 sky130_fd_sc_hd__buf_2
X_13861_ clknet_leaf_52_clk _01092_ net1175 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[849\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12812_ net1366 vssd1 vssd1 vccd1 vccd1 _00253_ sky130_fd_sc_hd__clkbuf_1
X_13792_ clknet_leaf_10_clk _01023_ net1098 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[780\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13506__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12743_ _05059_ _06373_ vssd1 vssd1 vccd1 vccd1 _06382_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_80_2923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_2300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12674_ _06324_ net1431 net979 vssd1 vssd1 vccd1 vccd1 _01339_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12008__A2 net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11625_ net216 net630 vssd1 vssd1 vccd1 vccd1 _06170_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_13_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13656__CLK clknet_leaf_65_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11556_ net218 net634 vssd1 vssd1 vccd1 vccd1 _06134_ sky130_fd_sc_hd__and2_1
Xwire541 _01995_ vssd1 vssd1 vccd1 vccd1 net541 sky130_fd_sc_hd__buf_4
XANTENNA__08632__A1 net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_2852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06904__A net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_2863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_2874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_2716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10507_ final_design.CPU_instr_adr\[3\] net1018 net1057 vssd1 vssd1 vccd1 vccd1 _05256_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_69_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_2885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12117__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_2727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11487_ net186 net2392 net308 vssd1 vssd1 vccd1 vccd1 _00365_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_74_2738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_2749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11519__B2 net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13226_ clknet_leaf_60_clk _00457_ net1140 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[214\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09774__X _04693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10438_ _02991_ net593 vssd1 vssd1 vccd1 vccd1 _05203_ sky130_fd_sc_hd__nor2_1
X_13157_ clknet_leaf_49_clk _00388_ net1181 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[145\]
+ sky130_fd_sc_hd__dfrtp_1
X_10369_ net11 net1025 net1008 final_design.data_from_mem\[18\] vssd1 vssd1 vccd1
+ vccd1 _00122_ sky130_fd_sc_hd__a22o_1
X_12108_ net1621 net210 net390 vssd1 vssd1 vccd1 vccd1 _00832_ sky130_fd_sc_hd__mux2_1
XANTENNA__10045__A1_N _04632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13088_ clknet_leaf_12_clk _00319_ net1090 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[76\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_23_clk_A clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13036__CLK clknet_leaf_46_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11257__A net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12039_ net1671 net212 net396 vssd1 vssd1 vccd1 vccd1 _00767_ sky130_fd_sc_hd__mux2_1
XANTENNA__09896__A0 net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12495__A2 net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06600_ final_design.cpu.reg_window\[412\] final_design.cpu.reg_window\[444\] net938
+ vssd1 vssd1 vccd1 vccd1 _01551_ sky130_fd_sc_hd__mux2_1
X_07580_ final_design.cpu.reg_window\[671\] final_design.cpu.reg_window\[703\] net857
+ vssd1 vssd1 vccd1 vccd1 _02531_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_38_clk_A clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13186__CLK clknet_leaf_11_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07470__A _01480_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06531_ _01454_ _01455_ _01458_ _01460_ vssd1 vssd1 vccd1 vccd1 _01482_ sky130_fd_sc_hd__nand4_4
XFILLER_0_73_1082 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09250_ _02670_ _02702_ _02671_ vssd1 vssd1 vccd1 vccd1 _04169_ sky130_fd_sc_hd__o21ba_1
X_06462_ _01405_ _01412_ _00211_ vssd1 vssd1 vccd1 vccd1 _01413_ sky130_fd_sc_hd__a21oi_1
X_08201_ _03148_ _03149_ _03150_ _03151_ net678 net701 vssd1 vssd1 vccd1 vccd1 _03152_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_51_1380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09181_ _04099_ vssd1 vssd1 vccd1 vccd1 _04100_ sky130_fd_sc_hd__inv_2
XANTENNA__08572__Y _03523_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08132_ net720 _03082_ vssd1 vssd1 vccd1 vccd1 _03083_ sky130_fd_sc_hd__nor2_1
XANTENNA__06814__A net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08063_ final_design.cpu.reg_window\[914\] final_design.cpu.reg_window\[946\] net844
+ vssd1 vssd1 vccd1 vccd1 _03014_ sky130_fd_sc_hd__mux2_1
XANTENNA__10430__B2 net245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12027__S net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07014_ _01959_ _01964_ net749 vssd1 vssd1 vccd1 vccd1 _01965_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1022_A _06298_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08965_ _03899_ _03900_ _03903_ net258 net1016 vssd1 vssd1 vccd1 vccd1 _03904_ sky130_fd_sc_hd__a221o_1
XANTENNA__08240__S net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout482_A net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07916_ net617 _02863_ _02865_ _01717_ vssd1 vssd1 vccd1 vccd1 _02867_ sky130_fd_sc_hd__a211oi_2
XANTENNA__10071__A net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08234__S0 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08896_ _02471_ net624 _03839_ _03841_ net256 vssd1 vssd1 vccd1 vccd1 _03842_ sky130_fd_sc_hd__a311o_1
XANTENNA__12486__A2 net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13529__CLK clknet_leaf_54_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11694__B1 net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07847_ _01788_ net617 vssd1 vssd1 vccd1 vccd1 _02798_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout270_X net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_32_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout747_A _01438_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout368_X net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06695__S net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07778_ _02725_ _02726_ _02727_ _02728_ net686 net694 vssd1 vssd1 vccd1 vccd1 _02729_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__09639__B1 net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07380__A _02326_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09517_ net484 _04435_ vssd1 vssd1 vccd1 vccd1 _04436_ sky130_fd_sc_hd__nand2_1
X_06729_ final_design.cpu.reg_window\[600\] final_design.cpu.reg_window\[632\] net942
+ vssd1 vssd1 vccd1 vccd1 _01680_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout914_A net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout535_X net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13679__CLK clknet_leaf_44_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09448_ net486 _04366_ vssd1 vssd1 vccd1 vccd1 _04367_ sky130_fd_sc_hd__nand2_1
XFILLER_0_52_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout702_X net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09379_ net478 _04097_ _04296_ vssd1 vssd1 vccd1 vccd1 _04298_ sky130_fd_sc_hd__or3_1
XPHY_EDGE_ROW_49_Left_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_23_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11410_ net1936 net232 net310 vssd1 vssd1 vccd1 vccd1 _00307_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_23_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12390_ net1767 net186 net271 vssd1 vssd1 vccd1 vccd1 _01101_ sky130_fd_sc_hd__mux2_1
XANTENNA__12410__A2 net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09811__B1 net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1885 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11341_ net432 net574 _06032_ net317 net1899 vssd1 vssd1 vccd1 vccd1 _00298_ sky130_fd_sc_hd__a32o_1
XFILLER_0_50_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14060_ clknet_leaf_16_clk _00022_ net1091 vssd1 vssd1 vccd1 vccd1 final_design.uart.BAUD_counter\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_11272_ _04509_ net653 _05843_ _05971_ vssd1 vssd1 vccd1 vccd1 _05972_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_28_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12174__A1 net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13059__CLK clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13011_ net1342 _00242_ net1228 vssd1 vssd1 vccd1 vccd1 final_design.CPU_instr_adr\[31\]
+ sky130_fd_sc_hd__dfrtp_2
X_10223_ final_design.uart.BAUD_counter\[7\] final_design.uart.BAUD_counter\[8\] _05099_
+ vssd1 vssd1 vccd1 vccd1 _05103_ sky130_fd_sc_hd__and3_1
XANTENNA_input43_A mem_adr_start[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10154_ _01384_ _05048_ vssd1 vssd1 vccd1 vccd1 _05052_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_7_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_58_Left_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_7_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10085_ final_design.VGA_data_control.v_count\[0\] _05000_ final_design.VGA_data_control.v_count\[5\]
+ vssd1 vssd1 vccd1 vccd1 _05001_ sky130_fd_sc_hd__o21ai_1
Xhold7 final_design.cpu.reg_window\[3\] vssd1 vssd1 vccd1 vccd1 net1349 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12477__A2 net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1612 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13913_ clknet_leaf_54_clk _01144_ net1177 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[901\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11364__X _06053_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07561__Y _02512_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13844_ clknet_leaf_8_clk _01075_ net1153 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[832\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_1905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08528__S1 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09725__S0 net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11524__B net196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13775_ clknet_leaf_43_clk _01006_ net1218 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[763\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10987_ _05710_ _05711_ _05713_ net1033 net1381 vssd1 vssd1 vccd1 vccd1 _00198_ sky130_fd_sc_hd__a32o_1
XFILLER_0_69_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12726_ final_design.VGA_data_control.v_count\[1\] _06366_ vssd1 vssd1 vccd1 vccd1
+ _06367_ sky130_fd_sc_hd__and2b_1
XFILLER_0_57_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07656__A2 _02602_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_67_Left_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12657_ final_design.VGA_data_control.ready_data\[16\] net1021 net976 final_design.data_from_mem\[16\]
+ vssd1 vssd1 vccd1 vccd1 _06316_ sky130_fd_sc_hd__a22o_1
XFILLER_0_5_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11540__A net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11608_ net2123 net299 _06161_ net430 vssd1 vssd1 vccd1 vccd1 _00436_ sky130_fd_sc_hd__a22o_1
XANTENNA__07408__A2 net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12588_ net1523 net998 net984 final_design.data_from_mem\[6\] vssd1 vssd1 vccd1 vccd1
+ _01281_ sky130_fd_sc_hd__a22o_1
XANTENNA__12401__A2 net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11204__A3 _05911_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08325__S net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11539_ net232 net2354 net302 vssd1 vssd1 vccd1 vccd1 _00403_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold407 final_design.cpu.reg_window\[479\] vssd1 vssd1 vccd1 vccd1 net1749 sky130_fd_sc_hd__dlygate4sd3_1
Xhold418 final_design.cpu.reg_window\[72\] vssd1 vssd1 vccd1 vccd1 net1760 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09945__A net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold429 final_design.cpu.reg_window\[640\] vssd1 vssd1 vccd1 vccd1 net1771 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_61_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12165__A1 net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13209_ clknet_leaf_57_clk _00440_ net1146 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[197\]
+ sky130_fd_sc_hd__dfrtp_1
X_14189_ net1248 vssd1 vssd1 vccd1 vccd1 gpio_oeb[1] sky130_fd_sc_hd__buf_2
XFILLER_0_42_1346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout909 net910 vssd1 vssd1 vccd1 vccd1 net909 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07592__A1 net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08750_ final_design.CPU_instr_adr\[6\] _02240_ vssd1 vssd1 vccd1 vccd1 _03701_ sky130_fd_sc_hd__or2_1
Xhold1107 final_design.cpu.reg_window\[825\] vssd1 vssd1 vccd1 vccd1 net2449 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1118 final_design.cpu.reg_window\[107\] vssd1 vssd1 vccd1 vccd1 net2460 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1129 final_design.cpu.reg_window\[497\] vssd1 vssd1 vccd1 vccd1 net2471 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12468__A2 net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07701_ final_design.cpu.reg_window\[219\] final_design.cpu.reg_window\[251\] net861
+ vssd1 vssd1 vccd1 vccd1 _02652_ sky130_fd_sc_hd__mux2_1
X_08681_ _02545_ _03610_ _03631_ _02542_ vssd1 vssd1 vccd1 vccd1 _03632_ sky130_fd_sc_hd__a211o_1
XFILLER_0_75_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08567__Y _03518_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07632_ net711 _02582_ vssd1 vssd1 vccd1 vccd1 _02583_ sky130_fd_sc_hd__nor2_1
XANTENNA__07471__Y _02422_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13821__CLK clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12310__S net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_1188 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07404__S net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07563_ _01488_ net734 net728 net662 vssd1 vssd1 vccd1 vccd1 _02514_ sky130_fd_sc_hd__or4_4
XFILLER_0_14_1404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09302_ net497 net594 _04111_ vssd1 vssd1 vccd1 vccd1 _04221_ sky130_fd_sc_hd__and3_1
X_06514_ _01458_ _01460_ _01461_ _01462_ vssd1 vssd1 vccd1 vccd1 _01465_ sky130_fd_sc_hd__a22o_2
XFILLER_0_0_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_17_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08583__X _03534_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07494_ _02129_ _02444_ vssd1 vssd1 vccd1 vccd1 _02445_ sky130_fd_sc_hd__nand2_1
XFILLER_0_64_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_17_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09233_ _03324_ _04151_ _04150_ vssd1 vssd1 vccd1 vccd1 _04152_ sky130_fd_sc_hd__o21ai_1
X_06445_ _01369_ _01398_ vssd1 vssd1 vccd1 vccd1 _01399_ sky130_fd_sc_hd__nand2_1
XANTENNA__13971__CLK clknet_leaf_40_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout230_A net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06950__S0 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11450__A net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout328_A net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09164_ _04080_ _04082_ net467 vssd1 vssd1 vccd1 vccd1 _04083_ sky130_fd_sc_hd__mux2_1
XANTENNA__08235__S net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_40_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08115_ _02064_ net611 vssd1 vssd1 vccd1 vccd1 _03066_ sky130_fd_sc_hd__nor2_1
XANTENNA__10403__B2 net246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09095_ net2525 net1013 _04018_ vssd1 vssd1 vccd1 vccd1 _00215_ sky130_fd_sc_hd__a21bo_1
XANTENNA__13201__CLK clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1237_A net1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09855__A _03627_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08046_ _02994_ _02995_ vssd1 vssd1 vccd1 vccd1 _02997_ sky130_fd_sc_hd__or2_1
Xhold930 final_design.cpu.reg_window\[496\] vssd1 vssd1 vccd1 vccd1 net2272 sky130_fd_sc_hd__dlygate4sd3_1
Xhold941 final_design.cpu.reg_window\[133\] vssd1 vssd1 vccd1 vccd1 net2283 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold952 final_design.cpu.reg_window\[641\] vssd1 vssd1 vccd1 vccd1 net2294 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout697_A net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold963 final_design.cpu.reg_window\[633\] vssd1 vssd1 vccd1 vccd1 net2305 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07258__S1 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold974 final_design.cpu.reg_window\[349\] vssd1 vssd1 vccd1 vccd1 net2316 sky130_fd_sc_hd__dlygate4sd3_1
Xhold985 final_design.cpu.reg_window\[989\] vssd1 vssd1 vccd1 vccd1 net2327 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1025_X net1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold996 final_design.cpu.reg_window\[804\] vssd1 vssd1 vccd1 vccd1 net2338 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13351__CLK clknet_leaf_58_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11609__B net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09997_ _04124_ _04915_ _04914_ _04911_ vssd1 vssd1 vccd1 vccd1 _04916_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout864_A net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08948_ final_design.CPU_instr_adr\[21\] _03888_ net1038 vssd1 vssd1 vccd1 vccd1
+ _00232_ sky130_fd_sc_hd__mux2_1
XANTENNA__08207__S0 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08879_ net621 _03826_ _03824_ net256 vssd1 vssd1 vccd1 vccd1 _03827_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout652_X net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10910_ net1042 _05636_ vssd1 vssd1 vccd1 vccd1 _05640_ sky130_fd_sc_hd__nor2_1
XFILLER_0_73_1829 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11890_ net224 net2293 net273 vssd1 vssd1 vccd1 vccd1 _00632_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07430__S1 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1228 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07314__S net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10841_ net960 _05572_ _05573_ net956 vssd1 vssd1 vccd1 vccd1 _05574_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_79_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout917_X net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13560_ clknet_leaf_65_clk _00791_ net1070 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[548\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12092__B1 net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10772_ _05347_ _05385_ _05502_ _05507_ vssd1 vssd1 vccd1 vccd1 _05508_ sky130_fd_sc_hd__a31oi_4
XFILLER_0_67_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12511_ _06173_ net351 net328 net1896 vssd1 vssd1 vccd1 vccd1 _01216_ sky130_fd_sc_hd__a22o_1
XFILLER_0_81_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13491_ clknet_leaf_39_clk _00722_ net1210 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[479\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12442_ net1635 net217 net334 vssd1 vssd1 vccd1 vccd1 _01149_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_258 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12373_ net1779 net219 net268 vssd1 vssd1 vccd1 vccd1 _01084_ sky130_fd_sc_hd__mux2_1
X_14112_ clknet_leaf_14_clk _01309_ net1103 vssd1 vssd1 vccd1 vccd1 final_design.reqhand.data_from_UART\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_65_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11324_ net589 net649 _06016_ vssd1 vssd1 vccd1 vccd1 _06018_ sky130_fd_sc_hd__and3_1
XFILLER_0_31_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14043_ clknet_leaf_16_clk _00035_ net1094 vssd1 vssd1 vccd1 vccd1 final_design.uart.BAUD_counter\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07556__Y _02507_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11255_ net644 _05953_ _05956_ vssd1 vssd1 vccd1 vccd1 _05957_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_82_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11355__C1 net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10206_ final_design.uart.BAUD_counter\[1\] final_design.uart.BAUD_counter\[0\] final_design.uart.BAUD_counter\[2\]
+ vssd1 vssd1 vccd1 vccd1 _05092_ sky130_fd_sc_hd__a21o_1
X_11186_ net651 _05893_ _05895_ vssd1 vssd1 vccd1 vccd1 _05896_ sky130_fd_sc_hd__and3_1
XFILLER_0_78_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10423__B _05190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10137_ net2544 net954 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.next_state\[1\]
+ sky130_fd_sc_hd__nor2_1
XANTENNA__13844__CLK clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11658__B1 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_13_Right_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10068_ _01495_ net251 _04044_ vssd1 vssd1 vccd1 vccd1 _04987_ sky130_fd_sc_hd__o21a_1
XFILLER_0_76_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13827_ clknet_leaf_1_clk _01058_ net1072 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[815\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13994__CLK clknet_leaf_60_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12083__B1 net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13758_ clknet_leaf_13_clk _00989_ net1099 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[746\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12709_ final_design.VGA_data_control.v_count\[4\] _06338_ _06343_ _06344_ vssd1
+ vssd1 vccd1 vccd1 _06350_ sky130_fd_sc_hd__a22o_1
XANTENNA__06837__B1 _01504_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13689_ clknet_leaf_57_clk _00920_ net1177 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[677\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13224__CLK clknet_leaf_41_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_22_Right_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11189__A2 net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold204 final_design.cpu.reg_window\[155\] vssd1 vssd1 vccd1 vccd1 net1546 sky130_fd_sc_hd__dlygate4sd3_1
Xhold215 final_design.cpu.reg_window\[851\] vssd1 vssd1 vccd1 vccd1 net1557 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold226 final_design.uart.BAUD_counter\[22\] vssd1 vssd1 vccd1 vccd1 net1568 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13374__CLK clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold237 final_design.cpu.reg_window\[584\] vssd1 vssd1 vccd1 vccd1 net1579 sky130_fd_sc_hd__dlygate4sd3_1
Xhold248 final_design.cpu.reg_window\[549\] vssd1 vssd1 vccd1 vccd1 net1590 sky130_fd_sc_hd__dlygate4sd3_1
X_09920_ _04778_ _04834_ net470 vssd1 vssd1 vccd1 vccd1 _04839_ sky130_fd_sc_hd__mux2_1
Xhold259 final_design.cpu.reg_window\[560\] vssd1 vssd1 vccd1 vccd1 net1601 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12305__S net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout706 _01752_ vssd1 vssd1 vccd1 vccd1 net706 sky130_fd_sc_hd__clkbuf_4
X_09851_ _04181_ _04769_ vssd1 vssd1 vccd1 vccd1 _04770_ sky130_fd_sc_hd__or2_1
Xfanout717 net718 vssd1 vssd1 vccd1 vccd1 net717 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08211__C1 net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11897__A0 net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout728 net730 vssd1 vssd1 vccd1 vccd1 net728 sky130_fd_sc_hd__clkbuf_4
XANTENNA_clkload15_A clknet_leaf_15_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1176 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08802_ _03670_ _03752_ vssd1 vssd1 vccd1 vccd1 _03753_ sky130_fd_sc_hd__or2_1
X_09782_ _04697_ _04699_ vssd1 vssd1 vccd1 vccd1 _04701_ sky130_fd_sc_hd__nand2_1
X_06994_ final_design.cpu.reg_window\[463\] final_design.cpu.reg_window\[495\] net891
+ vssd1 vssd1 vccd1 vccd1 _01945_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_31_Right_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_33_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08733_ _03683_ vssd1 vssd1 vccd1 vccd1 _03684_ sky130_fd_sc_hd__inv_2
XANTENNA__09306__A2 net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout180_A _06074_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08738__B _02097_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout278_A net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12040__S net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08664_ _02028_ _02061_ _03613_ vssd1 vssd1 vccd1 vccd1 _03615_ sky130_fd_sc_hd__o21a_1
XANTENNA__10321__B1 net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07134__S net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07615_ final_design.cpu.reg_window\[989\] final_design.cpu.reg_window\[1021\] net870
+ vssd1 vssd1 vccd1 vccd1 _02566_ sky130_fd_sc_hd__mux2_1
X_08595_ final_design.cpu.reg_window\[512\] final_design.cpu.reg_window\[544\] net825
+ vssd1 vssd1 vccd1 vccd1 _03546_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout445_A net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1187_A net1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07546_ final_design.cpu.reg_window\[671\] final_design.cpu.reg_window\[703\] net937
+ vssd1 vssd1 vccd1 vccd1 _02497_ sky130_fd_sc_hd__mux2_1
XANTENNA__12074__B1 net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12613__A2 net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11821__A0 net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout612_A _02513_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07477_ _02426_ _02427_ vssd1 vssd1 vccd1 vccd1 _02428_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_40_Right_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout233_X net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11180__A net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09216_ _03589_ _04134_ vssd1 vssd1 vccd1 vccd1 _04135_ sky130_fd_sc_hd__nand2_1
X_06428_ final_design.VGA_data_control.state\[0\] vssd1 vssd1 vccd1 vccd1 _01383_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_45_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10067__Y _04986_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13717__CLK clknet_leaf_58_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_984 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09147_ _04060_ _04065_ _03484_ vssd1 vssd1 vccd1 vccd1 _04066_ sky130_fd_sc_hd__mux2_2
XANTENNA_fanout400_X net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_1655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09078_ _03655_ _04002_ _04003_ net1037 vssd1 vssd1 vccd1 vccd1 _04004_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_9_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11179__X _05890_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08029_ final_design.cpu.reg_window\[787\] final_design.cpu.reg_window\[819\] net832
+ vssd1 vssd1 vccd1 vccd1 _02980_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_9_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold760 final_design.cpu.reg_window\[338\] vssd1 vssd1 vccd1 vccd1 net2102 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13867__CLK clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold771 final_design.cpu.reg_window\[421\] vssd1 vssd1 vccd1 vccd1 net2113 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11337__C1 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold782 final_design.cpu.reg_window\[267\] vssd1 vssd1 vccd1 vccd1 net2124 sky130_fd_sc_hd__dlygate4sd3_1
X_11040_ net88 _05737_ _05763_ vssd1 vssd1 vccd1 vccd1 _05764_ sky130_fd_sc_hd__a21o_1
XANTENNA__11888__A0 net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09545__A2 net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold793 final_design.cpu.reg_window\[373\] vssd1 vssd1 vccd1 vccd1 net2135 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout867_X net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11352__A2 net235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07833__A net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12891__CLK clknet_leaf_17_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12991_ net1322 _00222_ net1193 vssd1 vssd1 vccd1 vccd1 final_design.CPU_instr_adr\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12301__A1 net240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1773 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11942_ _06143_ net283 net409 net2009 vssd1 vssd1 vccd1 vccd1 _00677_ sky130_fd_sc_hd__a22o_1
XANTENNA__07403__S1 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11873_ net2352 net519 _06244_ net433 vssd1 vssd1 vccd1 vccd1 _00618_ sky130_fd_sc_hd__a22o_1
XANTENNA__13247__CLK clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1058 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13612_ clknet_leaf_45_clk _00843_ net1213 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[600\]
+ sky130_fd_sc_hd__dfrtp_1
X_10824_ net669 _05546_ _05557_ net966 _05556_ vssd1 vssd1 vccd1 vccd1 _05558_ sky130_fd_sc_hd__o221a_1
XANTENNA_input100_X net100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12065__B1 net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06736__X _01687_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11407__A3 _06090_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07167__S0 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13543_ clknet_leaf_62_clk _00774_ net1120 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[531\]
+ sky130_fd_sc_hd__dfrtp_1
X_10755_ _04040_ _05490_ _05491_ _04042_ vssd1 vssd1 vccd1 vccd1 _05492_ sky130_fd_sc_hd__a22o_1
XANTENNA__12080__A3 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11090__A net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13474_ clknet_leaf_4_clk _00705_ net1079 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[462\]
+ sky130_fd_sc_hd__dfrtp_1
X_10686_ net71 net1043 vssd1 vssd1 vccd1 vccd1 _05426_ sky130_fd_sc_hd__xnor2_1
XANTENNA__13397__CLK clknet_leaf_56_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12425_ _06112_ net355 net340 net1951 vssd1 vssd1 vccd1 vccd1 _01134_ sky130_fd_sc_hd__a22o_1
XANTENNA__10379__B1 net1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1608 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12356_ net2449 net362 net352 _06046_ vssd1 vssd1 vccd1 vccd1 _01068_ sky130_fd_sc_hd__a22o_1
XFILLER_0_77_16 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11591__A2 net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11307_ _04570_ net651 net588 _06002_ vssd1 vssd1 vccd1 vccd1 _06003_ sky130_fd_sc_hd__o211a_1
XANTENNA__10434__A _02929_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08419__S0 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12287_ net574 _06217_ net509 net371 net1655 vssd1 vssd1 vccd1 vccd1 _01002_ sky130_fd_sc_hd__a32o_1
XANTENNA__12125__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14026_ clknet_leaf_60_clk _01257_ net1141 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[1014\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11249__B net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11238_ net647 net568 net214 vssd1 vssd1 vccd1 vccd1 _05942_ sky130_fd_sc_hd__and3_1
XANTENNA__11879__B1 net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11169_ _05855_ _05880_ vssd1 vssd1 vccd1 vccd1 _05881_ sky130_fd_sc_hd__nand2_1
XANTENNA__14022__CLK clknet_leaf_51_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11265__A net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_1272 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14172__CLK clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07400_ final_design.cpu.reg_window\[642\] final_design.cpu.reg_window\[674\] net913
+ vssd1 vssd1 vccd1 vccd1 _02351_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07889__S net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08380_ final_design.cpu.reg_window\[326\] final_design.cpu.reg_window\[358\] net831
+ vssd1 vssd1 vccd1 vccd1 _03331_ sky130_fd_sc_hd__mux2_1
XANTENNA__06646__X _01597_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07331_ net749 _02275_ net745 vssd1 vssd1 vccd1 vccd1 _02282_ sky130_fd_sc_hd__o21a_1
XFILLER_0_9_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11803__B1 net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08275__A2 _03224_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12071__A3 net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_0_clk_X clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07262_ net533 _02212_ vssd1 vssd1 vccd1 vccd1 _02213_ sky130_fd_sc_hd__nor2_1
XFILLER_0_61_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09001_ net623 _03934_ _03935_ net255 _03933_ vssd1 vssd1 vccd1 vccd1 _03936_ sky130_fd_sc_hd__a311o_1
X_07193_ final_design.cpu.reg_window\[777\] final_design.cpu.reg_window\[809\] net891
+ vssd1 vssd1 vccd1 vccd1 _02144_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1817 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12035__S net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10790__B1 net1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07129__S net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09903_ net485 _04559_ _04560_ _04262_ _04120_ vssd1 vssd1 vccd1 vccd1 _04822_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_35_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout503 net504 vssd1 vssd1 vccd1 vccd1 net503 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11159__B net251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout514 net515 vssd1 vssd1 vccd1 vccd1 net514 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_67_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07538__A1 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout395_A _06263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout547 _01880_ vssd1 vssd1 vccd1 vccd1 net547 sky130_fd_sc_hd__dlymetal6s2s_1
X_09834_ _03229_ _04087_ net440 _03227_ _04752_ vssd1 vssd1 vccd1 vccd1 _04753_ sky130_fd_sc_hd__a221o_1
Xfanout558 net562 vssd1 vssd1 vccd1 vccd1 net558 sky130_fd_sc_hd__buf_2
XANTENNA_fanout1102_A net1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout569 net571 vssd1 vssd1 vccd1 vccd1 net569 sky130_fd_sc_hd__clkbuf_4
X_09765_ _04393_ _04402_ net470 vssd1 vssd1 vccd1 vccd1 _04684_ sky130_fd_sc_hd__mux2_1
X_06977_ final_design.cpu.reg_window\[912\] final_design.cpu.reg_window\[944\] net923
+ vssd1 vssd1 vccd1 vccd1 _01928_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout562_A net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1913 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08716_ final_design.CPU_instr_adr\[25\] _01660_ vssd1 vssd1 vccd1 vccd1 _03667_
+ sky130_fd_sc_hd__and2_1
XANTENNA__12295__B1 net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09696_ _01382_ _04185_ vssd1 vssd1 vccd1 vccd1 _04615_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_1_243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09160__B1 _03523_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08647_ _01658_ _02765_ vssd1 vssd1 vccd1 vccd1 _03598_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_29_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout350_X net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout827_A net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout448_X net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09138__S1 net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08578_ _03525_ _03526_ _03527_ _03528_ net678 net698 vssd1 vssd1 vccd1 vccd1 _03529_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__06556__X _01507_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12598__B2 final_design.data_from_mem\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07529_ final_design.cpu.reg_window\[479\] final_design.cpu.reg_window\[511\] net939
+ vssd1 vssd1 vccd1 vccd1 _02480_ sky130_fd_sc_hd__mux2_1
XANTENNA__09999__C1 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09299__B _03419_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10540_ net250 _04864_ vssd1 vssd1 vccd1 vccd1 _05287_ sky130_fd_sc_hd__and2b_1
XFILLER_0_0_1917 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10471_ net1438 net1030 net1002 _05222_ vssd1 vssd1 vccd1 vccd1 _00173_ sky130_fd_sc_hd__a22o_1
X_12210_ net577 _06138_ net510 net378 net1916 vssd1 vssd1 vccd1 vccd1 _00928_ sky130_fd_sc_hd__a32o_1
XFILLER_0_81_1917 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13190_ clknet_leaf_51_clk _00421_ net1168 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[178\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout984_X net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11573__A2 net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12141_ net214 net2479 net385 vssd1 vssd1 vccd1 vccd1 _00862_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14045__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12072_ net560 _05935_ net503 net392 net1711 vssd1 vssd1 vccd1 vccd1 _00797_ sky130_fd_sc_hd__a32o_1
Xhold590 final_design.cpu.reg_window\[336\] vssd1 vssd1 vccd1 vccd1 net1932 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11325__A2 net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11023_ _05735_ _05746_ net55 vssd1 vssd1 vccd1 vccd1 _05748_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_70_2582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06878__S net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_2593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11089__B2 net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12974_ clknet_leaf_21_clk _00211_ net1160 vssd1 vssd1 vccd1 vccd1 final_design.reqhand.current_client\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__12286__B1 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_2_clk_X clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11925_ _06128_ net281 net409 net2496 vssd1 vssd1 vccd1 vccd1 _00662_ sky130_fd_sc_hd__a22o_1
XANTENNA__11372__X _06060_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1817 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11856_ net215 net553 vssd1 vssd1 vccd1 vccd1 _06240_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_64_2386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_2397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10807_ _05524_ _05540_ vssd1 vssd1 vccd1 vccd1 _05542_ sky130_fd_sc_hd__nand2b_1
X_11787_ net2438 net414 net286 _05959_ vssd1 vssd1 vccd1 vccd1 _00544_ sky130_fd_sc_hd__a22o_1
XANTENNA__10429__A net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11261__A1 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10738_ net669 _05462_ _05475_ net965 _05474_ vssd1 vssd1 vccd1 vccd1 _05476_ sky130_fd_sc_hd__o221a_1
X_13526_ clknet_leaf_61_clk _00757_ net1137 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[514\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13457_ clknet_leaf_35_clk _00688_ net1240 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[445\]
+ sky130_fd_sc_hd__dfrtp_1
X_10669_ _05408_ _05409_ vssd1 vssd1 vccd1 vccd1 _05410_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_11_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12408_ _06240_ net499 net339 net2256 vssd1 vssd1 vccd1 vccd1 _01118_ sky130_fd_sc_hd__a22o_1
XANTENNA__12210__B1 net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13388_ clknet_leaf_45_clk _00619_ net1216 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[376\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_11_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput106 net106 vssd1 vssd1 vccd1 vccd1 ADR_O[14] sky130_fd_sc_hd__clkbuf_4
XANTENNA__12363__B net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_2179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07768__A1 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput117 net117 vssd1 vssd1 vccd1 vccd1 ADR_O[24] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_11_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput128 net128 vssd1 vssd1 vccd1 vccd1 ADR_O[5] sky130_fd_sc_hd__clkbuf_4
X_12339_ _06231_ net498 net360 net2193 vssd1 vssd1 vccd1 vccd1 _01051_ sky130_fd_sc_hd__a22o_1
Xoutput139 net139 vssd1 vssd1 vccd1 vccd1 DAT_O[14] sky130_fd_sc_hd__buf_2
X_14009_ clknet_leaf_56_clk _01240_ net1147 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[997\]
+ sky130_fd_sc_hd__dfrtp_1
X_06900_ _01468_ net736 net744 vssd1 vssd1 vccd1 vccd1 _01851_ sky130_fd_sc_hd__a21oi_4
XANTENNA__13412__CLK clknet_leaf_52_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07880_ _01504_ _01822_ net605 vssd1 vssd1 vccd1 vccd1 _02831_ sky130_fd_sc_hd__and3_1
XFILLER_0_78_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06831_ _01778_ _01779_ _01780_ _01781_ net778 net783 vssd1 vssd1 vccd1 vccd1 _01782_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__11707__B net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09550_ _04072_ _04468_ _04462_ _04464_ vssd1 vssd1 vccd1 vccd1 _04469_ sky130_fd_sc_hd__or4b_1
XANTENNA__12277__B1 net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06762_ final_design.cpu.reg_window\[599\] final_design.cpu.reg_window\[631\] net926
+ vssd1 vssd1 vccd1 vccd1 _01713_ sky130_fd_sc_hd__mux2_1
X_08501_ _02330_ net595 vssd1 vssd1 vccd1 vccd1 _03452_ sky130_fd_sc_hd__nand2_1
XANTENNA__13562__CLK clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09481_ _04056_ _04399_ vssd1 vssd1 vccd1 vccd1 _04400_ sky130_fd_sc_hd__or2_1
XFILLER_0_77_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06693_ net755 _01637_ net747 vssd1 vssd1 vccd1 vccd1 _01644_ sky130_fd_sc_hd__o21a_1
XFILLER_0_53_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12292__A3 net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08432_ _03377_ _03382_ net715 vssd1 vssd1 vccd1 vccd1 _03383_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08363_ _03310_ _03311_ _03312_ _03313_ net674 net696 vssd1 vssd1 vccd1 vccd1 _03314_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_73_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07314_ _02259_ _02264_ net752 vssd1 vssd1 vccd1 vccd1 _02265_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11252__A1 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07456__B1 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08294_ final_design.cpu.reg_window\[585\] final_design.cpu.reg_window\[617\] net807
+ vssd1 vssd1 vccd1 vccd1 _03245_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07245_ final_design.cpu.reg_window\[455\] final_design.cpu.reg_window\[487\] net892
+ vssd1 vssd1 vccd1 vccd1 _02196_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout310_A _06092_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout408_A net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1761 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12201__B1 net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07176_ net881 _02119_ _02125_ _02107_ _02113_ vssd1 vssd1 vccd1 vccd1 _02127_ sky130_fd_sc_hd__a32o_4
XANTENNA__14068__CLK clknet_leaf_15_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10074__A net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout300 net301 vssd1 vssd1 vccd1 vccd1 net300 sky130_fd_sc_hd__buf_4
XFILLER_0_1_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout311 _06092_ vssd1 vssd1 vccd1 vccd1 net311 sky130_fd_sc_hd__buf_4
XANTENNA_fanout777_A net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13092__CLK clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout398_X net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11307__A2 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout322 net323 vssd1 vssd1 vccd1 vccd1 net322 sky130_fd_sc_hd__buf_4
Xfanout333 _06283_ vssd1 vssd1 vccd1 vccd1 net333 sky130_fd_sc_hd__buf_4
XPHY_EDGE_ROW_21_Left_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout344 net345 vssd1 vssd1 vccd1 vccd1 net344 sky130_fd_sc_hd__clkbuf_4
Xfanout355 net358 vssd1 vssd1 vccd1 vccd1 net355 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09381__A0 net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1105_X net1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout366 net367 vssd1 vssd1 vccd1 vccd1 net366 sky130_fd_sc_hd__buf_6
XANTENNA__11617__B net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout377 _06271_ vssd1 vssd1 vccd1 vccd1 net377 sky130_fd_sc_hd__buf_4
X_09817_ _04378_ _04735_ net497 vssd1 vssd1 vccd1 vccd1 _04736_ sky130_fd_sc_hd__a21o_1
Xfanout388 net389 vssd1 vssd1 vccd1 vccd1 net388 sky130_fd_sc_hd__clkbuf_8
XANTENNA__13905__CLK clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10521__B net250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout399 _06261_ vssd1 vssd1 vccd1 vccd1 net399 sky130_fd_sc_hd__buf_4
XANTENNA_fanout944_A net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12268__B1 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1721 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09748_ _04261_ _04262_ net494 _04097_ vssd1 vssd1 vccd1 vccd1 _04667_ sky130_fd_sc_hd__a211o_1
XFILLER_0_69_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_1765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout732_X net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09679_ _04595_ _04596_ net730 _04594_ vssd1 vssd1 vccd1 vccd1 _04598_ sky130_fd_sc_hd__o211ai_4
XANTENNA__09684__A1 _04097_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12283__A3 net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11710_ net567 net422 _06213_ net295 net1647 vssd1 vssd1 vccd1 vccd1 _00486_ sky130_fd_sc_hd__a32o_1
XANTENNA__11633__A net207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12690_ _01383_ final_design.VGA_data_control.state\[1\] _06332_ vssd1 vssd1 vccd1
+ vccd1 _06333_ sky130_fd_sc_hd__or3_4
XFILLER_0_56_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08418__S net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07322__S net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11641_ net201 net633 vssd1 vssd1 vccd1 vccd1 _06178_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_30_Left_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09436__A1 net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09597__X _04516_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11572_ net203 net637 vssd1 vssd1 vccd1 vccd1 _06142_ sky130_fd_sc_hd__and2_1
XFILLER_0_80_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07998__A1 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13311_ clknet_leaf_7_clk _00542_ net1135 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[299\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput19 DAT_I[25] vssd1 vssd1 vccd1 vccd1 net19 sky130_fd_sc_hd__clkbuf_1
X_10523_ net94 final_design.VGA_adr\[2\] vssd1 vssd1 vccd1 vccd1 _05271_ sky130_fd_sc_hd__or2_1
XFILLER_0_68_1547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11066__A1_N net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13242_ clknet_leaf_1_clk _00473_ net1081 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[230\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input73_A memory_size[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10454_ _02668_ net593 vssd1 vssd1 vccd1 vccd1 _05211_ sky130_fd_sc_hd__nor2_1
XFILLER_0_21_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13173_ clknet_leaf_57_clk _00404_ net1132 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[161\]
+ sky130_fd_sc_hd__dfrtp_1
X_10385_ net1518 net1032 net1004 vssd1 vssd1 vccd1 vccd1 _00136_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_76_2791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13435__CLK clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_53_2010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1889 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_2021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12124_ net2281 net180 net390 vssd1 vssd1 vccd1 vccd1 _00848_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_53_2032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_72_2677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12055_ net2167 net182 net398 vssd1 vssd1 vccd1 vccd1 _00783_ sky130_fd_sc_hd__mux2_1
X_11006_ net53 _05708_ _05712_ vssd1 vssd1 vccd1 vccd1 _05732_ sky130_fd_sc_hd__a21oi_1
XANTENNA__13585__CLK clknet_leaf_34_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11019__S net1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12259__B1 net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08676__X _03627_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_66_2448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12957_ clknet_leaf_29_clk _00195_ net1196 vssd1 vssd1 vccd1 vccd1 net115 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12274__A3 net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1603 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11908_ net804 _06246_ vssd1 vssd1 vccd1 vccd1 _06248_ sky130_fd_sc_hd__nor2_4
XFILLER_0_59_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12888_ clknet_leaf_17_clk _00126_ net1109 vssd1 vssd1 vccd1 vccd1 final_design.data_from_mem\[22\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_73_1297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11839_ net183 net2227 net266 vssd1 vssd1 vccd1 vccd1 _00591_ sky130_fd_sc_hd__mux2_1
XANTENNA__11785__A2 net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13509_ clknet_leaf_49_clk _00740_ net1184 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[497\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08650__A2 _02668_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1901 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07030_ net758 _01980_ vssd1 vssd1 vccd1 vccd1 _01981_ sky130_fd_sc_hd__or2_2
XANTENNA__10606__B final_design.VGA_adr\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14219__1277 vssd1 vssd1 vccd1 vccd1 _14219__1277/HI net1277 sky130_fd_sc_hd__conb_1
XFILLER_0_2_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_1208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08981_ _03793_ _03917_ vssd1 vssd1 vccd1 vccd1 _03918_ sky130_fd_sc_hd__or2_1
XANTENNA__13928__CLK clknet_leaf_41_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_1680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07932_ final_design.cpu.reg_window\[790\] final_design.cpu.reg_window\[822\] net837
+ vssd1 vssd1 vccd1 vccd1 _02883_ sky130_fd_sc_hd__mux2_1
XANTENNA__12313__S net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12498__B1 net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08166__A1 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08299__A net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1120 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_1697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07863_ final_design.cpu.reg_window\[212\] final_design.cpu.reg_window\[244\] net868
+ vssd1 vssd1 vccd1 vccd1 _02814_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_3_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09602_ _04074_ _04440_ _04517_ net497 _04520_ vssd1 vssd1 vccd1 vccd1 _04521_ sky130_fd_sc_hd__o221a_1
X_06814_ net763 _01764_ vssd1 vssd1 vccd1 vccd1 _01765_ sky130_fd_sc_hd__or2_1
XANTENNA__12952__CLK clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07794_ final_design.cpu.reg_window\[89\] final_design.cpu.reg_window\[121\] net855
+ vssd1 vssd1 vccd1 vccd1 _02745_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_1440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09533_ net729 _04429_ _04450_ vssd1 vssd1 vccd1 vccd1 _04452_ sky130_fd_sc_hd__nand3_2
XFILLER_0_79_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06745_ final_design.cpu.reg_window\[407\] final_design.cpu.reg_window\[439\] net929
+ vssd1 vssd1 vccd1 vccd1 _01696_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08469__A2 _03415_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12265__A3 net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout358_A net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09464_ _02735_ _02769_ _04281_ net448 vssd1 vssd1 vccd1 vccd1 _04383_ sky130_fd_sc_hd__a31o_1
X_06676_ net884 _01619_ _01625_ _01612_ _01613_ vssd1 vssd1 vccd1 vccd1 _01627_ sky130_fd_sc_hd__a32o_2
XANTENNA__13308__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08415_ final_design.cpu.reg_window\[69\] final_design.cpu.reg_window\[101\] net840
+ vssd1 vssd1 vccd1 vccd1 _03366_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09418__A1 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09395_ _02576_ _04087_ net442 _02575_ vssd1 vssd1 vccd1 vccd1 _04314_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_47_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11225__A1 final_design.data_from_mem\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08346_ _02212_ net610 vssd1 vssd1 vccd1 vccd1 _03297_ sky130_fd_sc_hd__or2_1
XFILLER_0_80_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12422__B1 net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09969__A2 net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08762__A net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06834__X _01785_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11776__A2 net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08277_ net599 _03224_ _03200_ net537 vssd1 vssd1 vccd1 vccd1 _03228_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout313_X net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13458__CLK clknet_leaf_38_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1055_X net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07228_ final_design.cpu.reg_window\[776\] final_design.cpu.reg_window\[808\] net897
+ vssd1 vssd1 vccd1 vccd1 _02179_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_1433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07159_ final_design.cpu.reg_window\[202\] final_design.cpu.reg_window\[234\] net896
+ vssd1 vssd1 vccd1 vccd1 _02110_ sky130_fd_sc_hd__mux2_1
XANTENNA__09051__C1 net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07827__S1 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10170_ final_design.vga.h_current_state\[0\] _05009_ vssd1 vssd1 vccd1 vccd1 _05062_
+ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout682_X net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1106 net1107 vssd1 vssd1 vccd1 vccd1 net1106 sky130_fd_sc_hd__clkbuf_4
Xfanout1117 net1118 vssd1 vssd1 vccd1 vccd1 net1117 sky130_fd_sc_hd__clkbuf_2
XANTENNA__12489__B1 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1128 net1129 vssd1 vssd1 vccd1 vccd1 net1128 sky130_fd_sc_hd__clkbuf_4
XANTENNA_clkbuf_3_6_0_clk_X clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1139 net1150 vssd1 vssd1 vccd1 vccd1 net1139 sky130_fd_sc_hd__clkbuf_2
Xfanout185 _06060_ vssd1 vssd1 vccd1 vccd1 net185 sky130_fd_sc_hd__clkbuf_2
XANTENNA__11700__A2 net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout196 _06016_ vssd1 vssd1 vccd1 vccd1 net196 sky130_fd_sc_hd__clkbuf_2
X_13860_ clknet_leaf_52_clk _01091_ net1171 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[848\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09106__A0 net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12811_ net1374 vssd1 vssd1 vccd1 vccd1 _00252_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13791_ clknet_leaf_7_clk _01022_ net1130 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[779\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_1404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12256__A3 _06264_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1901 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07560__B _01480_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12742_ _06359_ _06379_ vssd1 vssd1 vccd1 vccd1 _06381_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_80_2924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_2301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07052__S net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_2946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_69_Right_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12673_ final_design.VGA_data_control.ready_data\[24\] net1020 net975 final_design.data_from_mem\[24\]
+ vssd1 vssd1 vccd1 vccd1 _06324_ sky130_fd_sc_hd__a22o_1
XFILLER_0_56_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07987__S net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11624_ net557 net420 _06169_ net298 net1492 vssd1 vssd1 vccd1 vccd1 _00444_ sky130_fd_sc_hd__a32o_1
XANTENNA__12413__B1 net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11216__B2 net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_13_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_1500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11555_ net425 net559 _06133_ net302 net1691 vssd1 vssd1 vccd1 vccd1 _00411_ sky130_fd_sc_hd__a32o_1
XANTENNA__11810__B net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_78_2853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_2230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_2864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10506_ _05235_ _05254_ vssd1 vssd1 vccd1 vccd1 _05255_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_78_2875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_2717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11486_ net186 net640 vssd1 vssd1 vccd1 vccd1 _06111_ sky130_fd_sc_hd__and2_1
XFILLER_0_29_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_74_2728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_74_2739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11519__A2 _06120_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13225_ clknet_leaf_36_clk _00456_ net1229 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[213\]
+ sky130_fd_sc_hd__dfrtp_1
X_10437_ net253 _05202_ net1030 net2540 vssd1 vssd1 vccd1 vccd1 _00159_ sky130_fd_sc_hd__a2bb2o_1
XPHY_EDGE_ROW_78_Right_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13156_ clknet_leaf_55_clk _00387_ net1187 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[144\]
+ sky130_fd_sc_hd__dfrtp_1
X_10368_ net10 net1026 _05170_ final_design.data_from_mem\[17\] vssd1 vssd1 vccd1
+ vccd1 _00121_ sky130_fd_sc_hd__a22o_1
X_12107_ net1766 net212 net388 vssd1 vssd1 vccd1 vccd1 _00831_ sky130_fd_sc_hd__mux2_1
XANTENNA__12975__CLK clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12133__S net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10442__A _02797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13087_ clknet_leaf_8_clk _00318_ net1154 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[75\]
+ sky130_fd_sc_hd__dfrtp_1
X_10299_ _05149_ _05151_ _05152_ _01384_ vssd1 vssd1 vccd1 vccd1 _05153_ sky130_fd_sc_hd__o22a_1
X_12038_ net1648 net214 net397 vssd1 vssd1 vccd1 vccd1 _00766_ sky130_fd_sc_hd__mux2_1
XANTENNA__11257__B net209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09896__A1 net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11152__B1 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07751__A _01626_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13989_ clknet_leaf_49_clk _01220_ net1181 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[977\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12247__A3 net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11273__A net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06530_ _01478_ _01479_ vssd1 vssd1 vccd1 vccd1 _01481_ sky130_fd_sc_hd__and2_2
XANTENNA__12983__RESET_B net1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07470__B net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_1619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06461_ net1057 final_design.reqhand.current_client\[1\] net1041 vssd1 vssd1 vccd1
+ vccd1 _00211_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08200_ final_design.cpu.reg_window\[910\] final_design.cpu.reg_window\[942\] net825
+ vssd1 vssd1 vccd1 vccd1 _03151_ sky130_fd_sc_hd__mux2_1
XANTENNA__11560__X _06136_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13600__CLK clknet_leaf_11_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12404__B1 net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09180_ net478 _04098_ vssd1 vssd1 vccd1 vccd1 _04099_ sky130_fd_sc_hd__or2_1
XFILLER_0_69_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08131_ _03078_ _03079_ _03080_ _03081_ net682 net702 vssd1 vssd1 vccd1 vccd1 _03082_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__12308__S net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08062_ final_design.cpu.reg_window\[978\] final_design.cpu.reg_window\[1010\] net845
+ vssd1 vssd1 vccd1 vccd1 _03013_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkload45_A clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07013_ _01960_ _01961_ _01962_ _01963_ net764 net780 vssd1 vssd1 vccd1 vccd1 _01964_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__13750__CLK clknet_leaf_60_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11391__B1 _01491_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1038 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06493__S0 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12043__S net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08964_ _03902_ vssd1 vssd1 vccd1 vccd1 _03903_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout1015_A net1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07915_ net606 _02863_ _02839_ _01717_ vssd1 vssd1 vccd1 vccd1 _02866_ sky130_fd_sc_hd__o211a_1
X_08895_ net624 _03840_ vssd1 vssd1 vccd1 vccd1 _03841_ sky130_fd_sc_hd__nor2_1
XANTENNA__09887__A1 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08234__S1 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11143__B1 net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout475_A net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11694__A1 net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07846_ net877 _02796_ _02785_ _02784_ vssd1 vssd1 vccd1 vccd1 _02797_ sky130_fd_sc_hd__o2bb2a_2
XTAP_TAPCELL_ROW_32_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13130__CLK clknet_leaf_61_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09205__X _04124_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07777_ final_design.cpu.reg_window\[536\] final_design.cpu.reg_window\[568\] net855
+ vssd1 vssd1 vccd1 vccd1 _02728_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout642_A _05946_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12238__A3 net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout263_X net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06728_ _01675_ _01676_ _01677_ _01678_ net775 net784 vssd1 vssd1 vccd1 vccd1 _01679_
+ sky130_fd_sc_hd__mux4_1
X_09516_ _04337_ _04434_ net472 vssd1 vssd1 vccd1 vccd1 _04435_ sky130_fd_sc_hd__mux2_2
XFILLER_0_79_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07745__S0 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11997__A2 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09447_ net478 _04362_ _04363_ _04365_ _04293_ vssd1 vssd1 vccd1 vccd1 _04366_ sky130_fd_sc_hd__o32a_2
XFILLER_0_52_1156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06659_ final_design.cpu.reg_window\[26\] final_design.cpu.reg_window\[58\] net942
+ vssd1 vssd1 vccd1 vccd1 _01610_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout430_X net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_42_clk_X clknet_leaf_42_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout907_A net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13280__CLK clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09378_ net462 _04103_ _04257_ _04223_ net454 vssd1 vssd1 vccd1 vccd1 _04297_ sky130_fd_sc_hd__a32o_1
XANTENNA__12848__CLK clknet_leaf_18_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_23_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08329_ _03276_ _03277_ _03278_ _03279_ net675 net697 vssd1 vssd1 vccd1 vccd1 _03280_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_23_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11340_ net650 net193 vssd1 vssd1 vccd1 vccd1 _06032_ sky130_fd_sc_hd__and2_1
XFILLER_0_1_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_57_clk_X clknet_leaf_57_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11271_ net645 _05967_ _05970_ vssd1 vssd1 vccd1 vccd1 _05971_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09024__C1 net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13010_ net1341 _00241_ net1231 vssd1 vssd1 vccd1 vccd1 final_design.CPU_instr_adr\[30\]
+ sky130_fd_sc_hd__dfrtp_2
X_10222_ final_design.uart.BAUD_counter\[7\] final_design.uart.BAUD_counter\[6\] _05098_
+ final_design.uart.BAUD_counter\[8\] vssd1 vssd1 vccd1 vccd1 _05102_ sky130_fd_sc_hd__a31o_1
XFILLER_0_43_1859 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11382__B1 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10153_ _05050_ vssd1 vssd1 vccd1 vccd1 _05051_ sky130_fd_sc_hd__inv_2
XANTENNA__06484__S0 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input36_A mem_adr_start[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10084_ net1051 final_design.VGA_data_control.v_count\[2\] final_design.VGA_data_control.v_count\[3\]
+ final_design.VGA_data_control.v_count\[1\] vssd1 vssd1 vccd1 vccd1 _05000_ sky130_fd_sc_hd__or4_2
Xhold8 final_design.cpu.reg_window\[27\] vssd1 vssd1 vccd1 vccd1 net1350 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_1624 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13912_ clknet_leaf_64_clk _01143_ net1074 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[900\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_67_2510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06739__X _01690_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13843_ clknet_leaf_40_clk _01074_ net1211 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[831\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13623__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10986_ net1005 _05712_ vssd1 vssd1 vccd1 vccd1 _05713_ sky130_fd_sc_hd__nor2_1
X_13774_ clknet_leaf_43_clk _01005_ net1221 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[762\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09725__S1 net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11524__C _06116_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14218__1276 vssd1 vssd1 vccd1 vccd1 _14218__1276/HI net1276 sky130_fd_sc_hd__conb_1
XFILLER_0_15_1917 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14177__Q final_design.VGA_adr\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11988__A2 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12725_ _06363_ _06365_ _06361_ vssd1 vssd1 vccd1 vccd1 _06366_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_31_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11380__X _06067_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06864__A1 net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12656_ _06315_ net1440 net979 vssd1 vssd1 vccd1 vccd1 _01330_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08833__C net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13773__CLK clknet_leaf_48_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11540__B net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11607_ net228 net566 net631 vssd1 vssd1 vccd1 vccd1 _06161_ sky130_fd_sc_hd__and3_1
X_12587_ net2388 net998 net984 final_design.data_from_mem\[5\] vssd1 vssd1 vccd1 vccd1
+ _01280_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06616__A1 net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11538_ net671 _05848_ _06124_ vssd1 vssd1 vccd1 vccd1 _06125_ sky130_fd_sc_hd__or3_4
XFILLER_0_0_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold408 final_design.cpu.reg_window\[559\] vssd1 vssd1 vccd1 vccd1 net1750 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold419 final_design.cpu.reg_window\[837\] vssd1 vssd1 vccd1 vccd1 net1761 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14129__CLK clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11469_ net209 net2453 net308 vssd1 vssd1 vccd1 vccd1 _00352_ sky130_fd_sc_hd__mux2_1
XANTENNA__09015__C1 net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09566__A0 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13208_ clknet_leaf_65_clk _00439_ net1073 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[196\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14188_ net1247 vssd1 vssd1 vccd1 vccd1 gpio_oeb[0] sky130_fd_sc_hd__buf_2
XANTENNA__06650__A _01596_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13139_ clknet_leaf_37_clk _00370_ net1228 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[127\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_1781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07592__A2 _02540_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13153__CLK clknet_leaf_49_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1108 final_design.cpu.reg_window\[1020\] vssd1 vssd1 vccd1 vccd1 net2450 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1119 final_design.cpu.reg_window\[318\] vssd1 vssd1 vccd1 vccd1 net2461 sky130_fd_sc_hd__dlygate4sd3_1
X_07700_ final_design.cpu.reg_window\[27\] final_design.cpu.reg_window\[59\] net861
+ vssd1 vssd1 vccd1 vccd1 _02651_ sky130_fd_sc_hd__mux2_1
X_08680_ _03617_ net594 vssd1 vssd1 vccd1 vccd1 _03631_ sky130_fd_sc_hd__nand2_4
XANTENNA__06796__S net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11676__B2 net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07631_ _02578_ _02579_ _02580_ _02581_ net687 net705 vssd1 vssd1 vccd1 vccd1 _02582_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__11715__B net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07562_ _01489_ net731 net725 net660 vssd1 vssd1 vccd1 vccd1 _02513_ sky130_fd_sc_hd__and4_2
XFILLER_0_53_1443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09301_ net497 _04111_ vssd1 vssd1 vccd1 vccd1 _04220_ sky130_fd_sc_hd__nand2_1
XFILLER_0_49_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06513_ _01461_ _01462_ vssd1 vssd1 vccd1 vccd1 _01464_ sky130_fd_sc_hd__nand2_1
XFILLER_0_18_1574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11979__A2 net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07493_ _02130_ _02159_ _02443_ vssd1 vssd1 vccd1 vccd1 _02444_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_17_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_17_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09232_ _03325_ _03355_ vssd1 vssd1 vccd1 vccd1 _04151_ sky130_fd_sc_hd__nor2_1
X_06444_ final_design.VGA_data_control.v_count\[7\] final_design.VGA_data_control.v_count\[6\]
+ vssd1 vssd1 vccd1 vccd1 _01398_ sky130_fd_sc_hd__nor2_1
XFILLER_0_29_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09201__A net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06950__S1 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11450__B net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09163_ net552 net458 _04081_ vssd1 vssd1 vccd1 vccd1 _04082_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_25_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12038__S net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08114_ _03052_ _03053_ _03064_ net874 vssd1 vssd1 vccd1 vccd1 _03065_ sky130_fd_sc_hd__a22oi_4
XTAP_TAPCELL_ROW_40_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09094_ net255 _04016_ _04017_ _04013_ net1013 vssd1 vssd1 vccd1 vccd1 _04018_ sky130_fd_sc_hd__a221o_1
X_08045_ _02994_ _02995_ vssd1 vssd1 vccd1 vccd1 _02996_ sky130_fd_sc_hd__nor2_1
XANTENNA__10781__S net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold920 final_design.cpu.reg_window\[788\] vssd1 vssd1 vccd1 vccd1 net2262 sky130_fd_sc_hd__dlygate4sd3_1
Xhold931 final_design.cpu.reg_window\[999\] vssd1 vssd1 vccd1 vccd1 net2273 sky130_fd_sc_hd__dlygate4sd3_1
Xhold942 final_design.cpu.reg_window\[490\] vssd1 vssd1 vccd1 vccd1 net2284 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold953 final_design.cpu.reg_window\[552\] vssd1 vssd1 vccd1 vccd1 net2295 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08251__S net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold964 final_design.cpu.reg_window\[1012\] vssd1 vssd1 vccd1 vccd1 net2306 sky130_fd_sc_hd__dlygate4sd3_1
Xhold975 final_design.cpu.reg_window\[663\] vssd1 vssd1 vccd1 vccd1 net2317 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout592_A net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold986 final_design.cpu.reg_window\[566\] vssd1 vssd1 vccd1 vccd1 net2328 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold997 final_design.cpu.reg_window\[352\] vssd1 vssd1 vccd1 vccd1 net2339 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09996_ _02738_ _03594_ vssd1 vssd1 vccd1 vccd1 _04915_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout1018_X net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07943__X _02894_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08947_ _03885_ _03887_ net258 vssd1 vssd1 vccd1 vccd1 _03888_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout380_X net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08207__S1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout857_A net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13646__CLK clknet_leaf_44_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10810__A net1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08878_ _03775_ _03825_ vssd1 vssd1 vccd1 vccd1 _03826_ sky130_fd_sc_hd__nor2_1
XFILLER_0_38_1917 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11625__B net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07829_ final_design.cpu.reg_window\[277\] final_design.cpu.reg_window\[309\] net858
+ vssd1 vssd1 vccd1 vccd1 _02780_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout645_X net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10840_ final_design.CPU_instr_adr\[19\] _03903_ net1060 vssd1 vssd1 vccd1 vccd1
+ _05573_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_15_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13796__CLK clknet_leaf_51_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10771_ _05403_ _05502_ _05505_ _05506_ vssd1 vssd1 vccd1 vccd1 _05507_ sky130_fd_sc_hd__a211o_1
XANTENNA__12092__A1 net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10956__S net1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12510_ _06172_ net344 net326 net1573 vssd1 vssd1 vccd1 vccd1 _01215_ sky130_fd_sc_hd__a22o_1
XFILLER_0_26_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13490_ clknet_leaf_39_clk _00721_ net1205 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[478\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12441_ net1866 net219 net334 vssd1 vssd1 vccd1 vccd1 _01148_ sky130_fd_sc_hd__mux2_1
XANTENNA__09111__A final_design.CPU_instr_adr\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_22_clk_A clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13026__CLK clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08143__S0 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08599__A1 net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09796__B1 net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12372_ net2309 net221 net268 vssd1 vssd1 vccd1 vccd1 _01083_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11323_ net589 net196 vssd1 vssd1 vccd1 vccd1 _06017_ sky130_fd_sc_hd__and2_2
X_14111_ clknet_leaf_13_clk _01308_ net1100 vssd1 vssd1 vccd1 vccd1 final_design.reqhand.data_from_UART\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10691__S net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14042_ clknet_leaf_15_clk _00034_ net1095 vssd1 vssd1 vccd1 vccd1 final_design.uart.BAUD_counter\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_11254_ _02030_ net641 _05954_ _05955_ net658 vssd1 vssd1 vccd1 vccd1 _05956_ sky130_fd_sc_hd__a221o_1
XANTENNA__13176__CLK clknet_leaf_65_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_37_clk_A clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11088__A net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10205_ _05083_ net799 _05091_ vssd1 vssd1 vccd1 vccd1 _00017_ sky130_fd_sc_hd__and3_1
XFILLER_0_66_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11185_ _05855_ _05894_ vssd1 vssd1 vccd1 vccd1 _05895_ sky130_fd_sc_hd__nand2_1
X_10136_ _01383_ final_design.VGA_data_control.state\[1\] net954 vssd1 vssd1 vccd1
+ vccd1 final_design.VGA_data_control.next_state\[0\] sky130_fd_sc_hd__a21o_1
X_10067_ _04198_ _04983_ _04984_ _04985_ vssd1 vssd1 vccd1 vccd1 _04986_ sky130_fd_sc_hd__nand4_4
XANTENNA__11122__A3 net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09720__B1 net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10330__B2 final_design.data_from_mem\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkload1_A clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12607__B1 net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13826_ clknet_leaf_4_clk _01057_ net1084 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[814\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09079__A2 net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07709__S0 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12083__A1 net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13757_ clknet_leaf_2_clk _00988_ net1065 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[745\]
+ sky130_fd_sc_hd__dfrtp_1
X_10969_ _04385_ net249 net669 vssd1 vssd1 vccd1 vccd1 _05696_ sky130_fd_sc_hd__a21o_1
XANTENNA__08826__A2 _01539_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08382__S0 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12708_ final_design.VGA_data_control.v_count\[3\] _06348_ _06347_ vssd1 vssd1 vccd1
+ vccd1 _06349_ sky130_fd_sc_hd__o21ba_1
X_13688_ clknet_leaf_65_clk _00919_ net1073 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[676\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08039__B1 net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12639_ final_design.VGA_data_control.ready_data\[7\] net1021 net976 final_design.data_from_mem\[7\]
+ vssd1 vssd1 vccd1 vccd1 _06307_ sky130_fd_sc_hd__a22o_1
XFILLER_0_26_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13519__CLK clknet_leaf_42_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold205 final_design.cpu.reg_window\[135\] vssd1 vssd1 vccd1 vccd1 net1547 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07747__Y _02698_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold216 final_design.cpu.reg_window\[681\] vssd1 vssd1 vccd1 vccd1 net1558 sky130_fd_sc_hd__dlygate4sd3_1
Xhold227 final_design.cpu.reg_window\[721\] vssd1 vssd1 vccd1 vccd1 net1569 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09539__A0 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold238 final_design.VGA_data_control.data_to_VGA\[8\] vssd1 vssd1 vccd1 vccd1 net1580
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold249 final_design.cpu.reg_window\[857\] vssd1 vssd1 vccd1 vccd1 net1591 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_46_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09850_ net98 _04180_ vssd1 vssd1 vccd1 vccd1 _04769_ sky130_fd_sc_hd__nor2_1
XANTENNA__13669__CLK clknet_leaf_49_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout707 net709 vssd1 vssd1 vccd1 vccd1 net707 sky130_fd_sc_hd__clkbuf_4
Xfanout718 _01720_ vssd1 vssd1 vccd1 vccd1 net718 sky130_fd_sc_hd__buf_4
Xfanout729 net730 vssd1 vssd1 vccd1 vccd1 net729 sky130_fd_sc_hd__buf_4
X_08801_ _03671_ _03751_ _03672_ vssd1 vssd1 vccd1 vccd1 _03752_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_42_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09781_ _04697_ _04699_ vssd1 vssd1 vccd1 vccd1 _04700_ sky130_fd_sc_hd__nor2_1
X_06993_ final_design.cpu.reg_window\[271\] final_design.cpu.reg_window\[303\] net891
+ vssd1 vssd1 vccd1 vccd1 _01944_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_1431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11285__X _05983_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08732_ _03681_ _03682_ vssd1 vssd1 vccd1 vccd1 _03683_ sky130_fd_sc_hd__and2_1
XANTENNA__12321__S net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09841__D _04759_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07415__S net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08663_ _01999_ _02061_ _02029_ vssd1 vssd1 vccd1 vccd1 _03614_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10321__B2 final_design.data_from_mem\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07614_ final_design.cpu.reg_window\[797\] final_design.cpu.reg_window\[829\] net871
+ vssd1 vssd1 vccd1 vccd1 _02565_ sky130_fd_sc_hd__mux2_1
X_08594_ final_design.cpu.reg_window\[576\] final_design.cpu.reg_window\[608\] net827
+ vssd1 vssd1 vccd1 vccd1 _03545_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07545_ final_design.cpu.reg_window\[735\] final_design.cpu.reg_window\[767\] net937
+ vssd1 vssd1 vccd1 vccd1 _02496_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13049__CLK clknet_leaf_56_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout340_A net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1082_A net1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout438_A _04095_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10624__A2 net247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07476_ _02390_ _02394_ vssd1 vssd1 vccd1 vccd1 _02427_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_23_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06555__A net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06427_ net73 vssd1 vssd1 vccd1 vccd1 _01382_ sky130_fd_sc_hd__inv_2
X_09215_ _02997_ _03029_ vssd1 vssd1 vccd1 vccd1 _04134_ sky130_fd_sc_hd__nor2_1
X_09146_ net465 _04064_ _04062_ vssd1 vssd1 vccd1 vccd1 _04065_ sky130_fd_sc_hd__o21a_1
XFILLER_0_60_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13199__CLK clknet_leaf_42_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11585__B1 net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09077_ net620 _04001_ _03999_ net254 vssd1 vssd1 vccd1 vccd1 _04003_ sky130_fd_sc_hd__a211o_1
XFILLER_0_62_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08028_ final_design.cpu.reg_window\[851\] final_design.cpu.reg_window\[883\] net830
+ vssd1 vssd1 vccd1 vccd1 _02979_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_9_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold750 final_design.cpu.reg_window\[387\] vssd1 vssd1 vccd1 vccd1 net2092 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout974_A _06299_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11337__B1 _06028_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold761 final_design.cpu.reg_window\[690\] vssd1 vssd1 vccd1 vccd1 net2103 sky130_fd_sc_hd__dlygate4sd3_1
X_14217__1275 vssd1 vssd1 vccd1 vccd1 _14217__1275/HI net1275 sky130_fd_sc_hd__conb_1
Xhold772 final_design.cpu.reg_window\[500\] vssd1 vssd1 vccd1 vccd1 net2114 sky130_fd_sc_hd__dlygate4sd3_1
Xhold783 final_design.cpu.reg_window\[485\] vssd1 vssd1 vccd1 vccd1 net2125 sky130_fd_sc_hd__dlygate4sd3_1
Xhold794 final_design.cpu.reg_window\[884\] vssd1 vssd1 vccd1 vccd1 net2136 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout762_X net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09979_ _04896_ _04897_ _04890_ _04894_ vssd1 vssd1 vccd1 vccd1 _04898_ sky130_fd_sc_hd__a211o_1
X_12990_ net1321 _00221_ net1193 vssd1 vssd1 vccd1 vccd1 final_design.CPU_instr_adr\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07325__S net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11941_ _06142_ net285 net410 net2375 vssd1 vssd1 vccd1 vccd1 _00676_ sky130_fd_sc_hd__a22o_1
XFILLER_0_77_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11872_ net193 net554 vssd1 vssd1 vccd1 vccd1 _06244_ sky130_fd_sc_hd__and2_1
XANTENNA__09540__S net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13611_ clknet_leaf_52_clk _00842_ net1183 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[599\]
+ sky130_fd_sc_hd__dfrtp_1
X_10823_ net1055 _05553_ net1000 final_design.CPU_instr_adr\[18\] vssd1 vssd1 vccd1
+ vccd1 _05557_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__07167__S1 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13542_ clknet_leaf_50_clk _00773_ net1172 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[530\]
+ sky130_fd_sc_hd__dfrtp_1
X_10754_ _01363_ _03930_ net1060 vssd1 vssd1 vccd1 vccd1 _05491_ sky130_fd_sc_hd__mux2_1
XANTENNA__07492__A1 net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10685_ _05410_ _05411_ _05408_ vssd1 vssd1 vccd1 vccd1 _05425_ sky130_fd_sc_hd__o21ba_1
X_13473_ clknet_leaf_49_clk _00704_ net1186 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[461\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_63_760 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09769__B1 net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12424_ _06111_ net355 net340 net2142 vssd1 vssd1 vccd1 vccd1 _01133_ sky130_fd_sc_hd__a22o_1
XANTENNA__08680__A _03617_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10379__B2 final_design.data_from_mem\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12355_ net2260 net362 net356 _06039_ vssd1 vssd1 vccd1 vccd1 _01067_ sky130_fd_sc_hd__a22o_1
XANTENNA__06471__Y _01422_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13811__CLK clknet_leaf_40_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11306_ net645 _05998_ _06001_ vssd1 vssd1 vccd1 vccd1 _06002_ sky130_fd_sc_hd__a21o_1
XFILLER_0_77_28 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12286_ net570 _06216_ net507 net369 net1609 vssd1 vssd1 vccd1 vccd1 _01001_ sky130_fd_sc_hd__a32o_1
XANTENNA__11328__B1 net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10434__B net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08419__S1 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14025_ clknet_leaf_37_clk _01256_ net1231 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[1013\]
+ sky130_fd_sc_hd__dfrtp_1
X_11237_ net591 _05939_ _05940_ vssd1 vssd1 vccd1 vccd1 _05941_ sky130_fd_sc_hd__and3_1
XFILLER_0_43_1486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12540__A2 net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11168_ final_design.reqhand.data_from_UART\[3\] final_design.data_from_mem\[3\]
+ net247 vssd1 vssd1 vccd1 vccd1 _05880_ sky130_fd_sc_hd__mux2_1
XANTENNA__10551__A1 _04042_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13961__CLK clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10551__B2 net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10119_ final_design.VGA_data_control.v_count\[6\] _05026_ vssd1 vssd1 vccd1 vccd1
+ _05029_ sky130_fd_sc_hd__or2_1
XANTENNA__11546__A net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12141__S net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06850__S0 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11099_ _05801_ _05805_ _05804_ vssd1 vssd1 vccd1 vccd1 _05820_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10450__A _02763_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07235__S net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11265__B net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_1246 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13809_ clknet_leaf_34_clk _01040_ net1243 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[797\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07330_ net757 _02280_ vssd1 vssd1 vccd1 vccd1 _02281_ sky130_fd_sc_hd__or2_1
XANTENNA__11281__A net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11803__B2 _06046_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13341__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07261_ net666 _01598_ vssd1 vssd1 vccd1 vccd1 _02212_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_41_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1891 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09000_ _02452_ _02454_ vssd1 vssd1 vccd1 vccd1 _03935_ sky130_fd_sc_hd__nand2_1
XANTENNA__12909__CLK clknet_leaf_61_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08107__S0 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12359__A2 net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09686__A net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_3_7_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_3_7_0_clk sky130_fd_sc_hd__clkbuf_8
X_07192_ final_design.cpu.reg_window\[841\] final_design.cpu.reg_window\[873\] net901
+ vssd1 vssd1 vccd1 vccd1 _02143_ sky130_fd_sc_hd__mux2_1
XANTENNA__11567__B1 net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12316__S net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13491__CLK clknet_leaf_39_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07918__B net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1829 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08983__A1 net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10790__A1 _05508_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09902_ _04340_ _04817_ _04818_ _04277_ _04118_ vssd1 vssd1 vccd1 vccd1 _04821_ sky130_fd_sc_hd__a32o_1
XFILLER_0_6_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout504 net516 vssd1 vssd1 vccd1 vccd1 net504 sky130_fd_sc_hd__clkbuf_4
Xfanout515 net516 vssd1 vssd1 vccd1 vccd1 net515 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12531__A2 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout537 _02126_ vssd1 vssd1 vccd1 vccd1 net537 sky130_fd_sc_hd__buf_2
X_09833_ _03228_ net444 vssd1 vssd1 vccd1 vccd1 _04752_ sky130_fd_sc_hd__nor2_1
Xfanout548 _01850_ vssd1 vssd1 vccd1 vccd1 net548 sky130_fd_sc_hd__buf_2
XANTENNA_fanout290_A _06228_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout559 net561 vssd1 vssd1 vccd1 vccd1 net559 sky130_fd_sc_hd__buf_2
XANTENNA_fanout388_A net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12051__S net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09764_ _04394_ _04396_ net475 vssd1 vssd1 vccd1 vccd1 _04683_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06976_ final_design.cpu.reg_window\[976\] final_design.cpu.reg_window\[1008\] net923
+ vssd1 vssd1 vccd1 vccd1 _01927_ sky130_fd_sc_hd__mux2_1
X_08715_ final_design.CPU_instr_adr\[25\] _01660_ vssd1 vssd1 vccd1 vccd1 _03666_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_74_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11098__A2 net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12295__A1 net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09695_ net729 _04613_ vssd1 vssd1 vccd1 vccd1 _04614_ sky130_fd_sc_hd__and2_1
XANTENNA__11890__S net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout555_A _05869_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout176_X net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08646_ _01686_ _02733_ vssd1 vssd1 vccd1 vccd1 _03597_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_29_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12047__A1 net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout722_A net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout343_X net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08577_ final_design.cpu.reg_window\[384\] final_design.cpu.reg_window\[416\] net828
+ vssd1 vssd1 vccd1 vccd1 _03528_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout1085_X net1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10058__B1 _04905_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07528_ final_design.cpu.reg_window\[287\] final_design.cpu.reg_window\[319\] net939
+ vssd1 vssd1 vccd1 vccd1 _02479_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout510_X net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07459_ final_design.cpu.reg_window\[960\] final_design.cpu.reg_window\[992\] net909
+ vssd1 vssd1 vccd1 vccd1 _02410_ sky130_fd_sc_hd__mux2_1
XANTENNA__11270__A2 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13834__CLK clknet_leaf_59_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10470_ net36 _05220_ vssd1 vssd1 vccd1 vccd1 _05222_ sky130_fd_sc_hd__xor2_1
X_09129_ _02771_ _03594_ vssd1 vssd1 vccd1 vccd1 _04048_ sky130_fd_sc_hd__nand2_1
XFILLER_0_33_988 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12140_ net216 net2189 net384 vssd1 vssd1 vccd1 vccd1 _00861_ sky130_fd_sc_hd__mux2_1
XANTENNA__13984__CLK clknet_leaf_11_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12071_ net556 _05929_ net502 net392 net1723 vssd1 vssd1 vccd1 vccd1 _00796_ sky130_fd_sc_hd__a32o_1
XFILLER_0_44_1773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold580 final_design.cpu.reg_window\[139\] vssd1 vssd1 vccd1 vccd1 net1922 sky130_fd_sc_hd__dlygate4sd3_1
Xhold591 final_design.cpu.reg_window\[448\] vssd1 vssd1 vccd1 vccd1 net1933 sky130_fd_sc_hd__dlygate4sd3_1
X_11022_ _05735_ _05746_ net55 vssd1 vssd1 vccd1 vccd1 _05747_ sky130_fd_sc_hd__o21bai_1
XANTENNA__12522__A2 net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09923__B1 _04838_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10533__A1 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_2583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10533__B2 net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11730__B1 net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_70_2594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13214__CLK clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07055__S net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12973_ net1312 _00210_ net1155 vssd1 vssd1 vccd1 vccd1 final_design.CPU_instr_adr\[1\]
+ sky130_fd_sc_hd__dfrtp_2
X_11924_ _06127_ net282 net409 net1948 vssd1 vssd1 vccd1 vccd1 _00661_ sky130_fd_sc_hd__a22o_1
XANTENNA__06894__S net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07162__B1 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13364__CLK clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11855_ _06105_ net279 net517 net2093 vssd1 vssd1 vccd1 vccd1 _00605_ sky130_fd_sc_hd__a22o_1
XFILLER_0_5_1829 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_2376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_2387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12589__A2 net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10806_ _05522_ _05525_ _05540_ vssd1 vssd1 vccd1 vccd1 _05541_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_64_2398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11786_ net2407 net412 net278 _05952_ vssd1 vssd1 vccd1 vccd1 _00543_ sky130_fd_sc_hd__a22o_1
XANTENNA__10429__B _05190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13525_ clknet_leaf_58_clk _00756_ net1132 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[513\]
+ sky130_fd_sc_hd__dfrtp_1
X_10737_ net1055 _05471_ net1000 final_design.CPU_instr_adr\[14\] vssd1 vssd1 vccd1
+ vccd1 _05475_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_67_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13456_ clknet_leaf_37_clk _00687_ net1232 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[444\]
+ sky130_fd_sc_hd__dfrtp_1
X_10668_ net69 final_design.VGA_adr\[8\] _05407_ vssd1 vssd1 vccd1 vccd1 _05409_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11549__B1 net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12407_ _06105_ net345 net338 net1935 vssd1 vssd1 vccd1 vccd1 _01117_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_11_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12136__S net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12210__A1 net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10599_ net65 _05330_ _05342_ vssd1 vssd1 vccd1 vccd1 _05344_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_11_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13387_ clknet_leaf_38_clk _00618_ net1189 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[375\]
+ sky130_fd_sc_hd__dfrtp_1
Xoutput107 net107 vssd1 vssd1 vccd1 vccd1 ADR_O[15] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_51_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput118 net118 vssd1 vssd1 vccd1 vccd1 ADR_O[25] sky130_fd_sc_hd__clkbuf_4
XANTENNA__08965__B2 net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput129 net129 vssd1 vssd1 vccd1 vccd1 ADR_O[6] sky130_fd_sc_hd__clkbuf_4
X_12338_ net2417 net360 net342 _05911_ vssd1 vssd1 vccd1 vccd1 _01050_ sky130_fd_sc_hd__a22o_1
XANTENNA__10490__A1_N net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09953__B net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12269_ net569 _06199_ net507 net369 net2372 vssd1 vssd1 vccd1 vccd1 _00984_ sky130_fd_sc_hd__a32o_1
X_14008_ clknet_leaf_63_clk _01239_ net1076 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[996\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12513__A2 net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09914__B1 net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11276__A net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06830_ final_design.cpu.reg_window\[533\] final_design.cpu.reg_window\[565\] net940
+ vssd1 vssd1 vccd1 vccd1 _01781_ sky130_fd_sc_hd__mux2_1
XANTENNA__12277__A1 net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13707__CLK clknet_leaf_52_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06761_ final_design.cpu.reg_window\[663\] final_design.cpu.reg_window\[695\] net929
+ vssd1 vssd1 vccd1 vccd1 _01712_ sky130_fd_sc_hd__mux2_1
X_08500_ _02330_ net608 vssd1 vssd1 vccd1 vccd1 _03451_ sky130_fd_sc_hd__nor2_1
X_06692_ net762 _01642_ vssd1 vssd1 vccd1 vccd1 _01643_ sky130_fd_sc_hd__or2_1
X_09480_ _04395_ _04398_ net491 vssd1 vssd1 vccd1 vccd1 _04399_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11723__B net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08431_ _03378_ _03379_ _03380_ _03381_ net680 net692 vssd1 vssd1 vccd1 vccd1 _03382_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_59_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06900__B1 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14216__1274 vssd1 vssd1 vccd1 vccd1 _14216__1274/HI net1274 sky130_fd_sc_hd__conb_1
XFILLER_0_74_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13857__CLK clknet_leaf_48_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08362_ final_design.cpu.reg_window\[903\] final_design.cpu.reg_window\[935\] net811
+ vssd1 vssd1 vccd1 vccd1 _03313_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_1221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07313_ _02260_ _02261_ _02262_ _02263_ net770 net789 vssd1 vssd1 vccd1 vccd1 _02264_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__07456__A1 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08293_ net716 _03243_ vssd1 vssd1 vccd1 vccd1 _03244_ sky130_fd_sc_hd__nor2_1
X_07244_ final_design.cpu.reg_window\[263\] final_design.cpu.reg_window\[295\] net892
+ vssd1 vssd1 vccd1 vccd1 _02195_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12881__CLK clknet_leaf_17_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07175_ net882 _02119_ _02125_ _02107_ _02113_ vssd1 vssd1 vccd1 vccd1 _02126_ sky130_fd_sc_hd__a32oi_4
XFILLER_0_67_1773 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12046__S net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout303_A _06125_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12752__A2 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11960__B1 net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11885__S net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13237__CLK clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1212_A net1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout301 _06159_ vssd1 vssd1 vccd1 vccd1 net301 sky130_fd_sc_hd__buf_4
XANTENNA__12504__A2 net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout312 net313 vssd1 vssd1 vccd1 vccd1 net312 sky130_fd_sc_hd__clkbuf_8
Xfanout323 _06285_ vssd1 vssd1 vccd1 vccd1 net323 sky130_fd_sc_hd__buf_4
Xfanout334 net335 vssd1 vssd1 vccd1 vccd1 net334 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_61_1394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout293_X net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11712__B1 net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout345 net350 vssd1 vssd1 vccd1 vccd1 net345 sky130_fd_sc_hd__buf_2
Xfanout356 net358 vssd1 vssd1 vccd1 vccd1 net356 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09381__A1 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11186__A net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09816_ net489 _04459_ _04734_ vssd1 vssd1 vccd1 vccd1 _04735_ sky130_fd_sc_hd__a21o_1
Xfanout367 _06275_ vssd1 vssd1 vccd1 vccd1 net367 sky130_fd_sc_hd__buf_6
XANTENNA_fanout1000_X net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout378 net379 vssd1 vssd1 vccd1 vccd1 net378 sky130_fd_sc_hd__buf_4
Xfanout389 _06265_ vssd1 vssd1 vccd1 vccd1 net389 sky130_fd_sc_hd__clkbuf_4
XANTENNA__13387__CLK clknet_leaf_38_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12268__A1 net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09747_ net484 _04664_ _04665_ vssd1 vssd1 vccd1 vccd1 _04666_ sky130_fd_sc_hd__a21oi_1
X_06959_ _01909_ vssd1 vssd1 vccd1 vccd1 _01910_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout937_A net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1733 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11914__A final_design.cpu.reg_window\[411\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09678_ _04595_ _04596_ _04594_ vssd1 vssd1 vccd1 vccd1 _04597_ sky130_fd_sc_hd__o21a_1
XFILLER_0_74_1777 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08341__C1 _02184_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11633__B net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08629_ net599 _03065_ _03041_ _02059_ vssd1 vssd1 vccd1 vccd1 _03580_ sky130_fd_sc_hd__o211a_1
XFILLER_0_51_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout725_X net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11228__C1 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11640_ net575 net424 _06177_ net301 net1575 vssd1 vssd1 vccd1 vccd1 _00452_ sky130_fd_sc_hd__a32o_1
XANTENNA__11779__B1 net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_2_0_clk_X clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11571_ net432 net572 _06141_ net305 net1566 vssd1 vssd1 vccd1 vccd1 _00419_ sky130_fd_sc_hd__a32o_1
XANTENNA__12440__A1 net221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10451__B1 net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13310_ clknet_leaf_9_clk _00541_ net1100 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[298\]
+ sky130_fd_sc_hd__dfrtp_1
X_10522_ net94 final_design.VGA_adr\[2\] vssd1 vssd1 vccd1 vccd1 _05270_ sky130_fd_sc_hd__nand2_1
XANTENNA__14012__CLK clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10453_ net1451 net1035 _05210_ net248 vssd1 vssd1 vccd1 vccd1 _00167_ sky130_fd_sc_hd__a22o_1
X_13241_ clknet_leaf_56_clk _00472_ net1146 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[229\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_1737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input66_A mem_adr_start[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1857 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13172_ clknet_leaf_12_clk _00403_ net1088 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[160\]
+ sky130_fd_sc_hd__dfrtp_1
X_10384_ net1 net1029 vssd1 vssd1 vccd1 vccd1 _05173_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_76_2792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_2011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06958__B1 _01821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11951__B1 net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_2022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12123_ net2248 net183 net390 vssd1 vssd1 vccd1 vccd1 _00847_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_72_2656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_2033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14162__CLK clknet_leaf_18_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_2678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12054_ net2331 net184 net398 vssd1 vssd1 vccd1 vccd1 _00782_ sky130_fd_sc_hd__mux2_1
XFILLER_0_40_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_1622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11005_ _05729_ _05730_ vssd1 vssd1 vccd1 vccd1 _05731_ sky130_fd_sc_hd__or2_1
XFILLER_0_74_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout890 net899 vssd1 vssd1 vccd1 vccd1 net890 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_5_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12956_ clknet_leaf_29_clk _00194_ net1196 vssd1 vssd1 vccd1 vccd1 net114 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11907_ net195 net2056 net273 vssd1 vssd1 vccd1 vccd1 _00649_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12887_ clknet_leaf_18_clk _00125_ net1107 vssd1 vssd1 vccd1 vccd1 final_design.data_from_mem\[21\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_5_1615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13136__RESET_B net1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11838_ net185 net2145 net267 vssd1 vssd1 vccd1 vccd1 _00590_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09427__A2 _04088_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07438__A1 net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11769_ net230 net2332 net412 vssd1 vssd1 vccd1 vccd1 _00531_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_40_clk clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_40_clk sky130_fd_sc_hd__clkbuf_8
X_13508_ clknet_leaf_54_clk _00739_ net1179 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[496\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13439_ clknet_leaf_7_clk _00670_ net1149 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[427\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_64_1913 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08938__A1 net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10745__B2 net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11942__B1 net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1367 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08980_ final_design.CPU_instr_adr\[17\] _03792_ vssd1 vssd1 vccd1 vccd1 _03917_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_48_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07931_ final_design.cpu.reg_window\[854\] final_design.cpu.reg_window\[886\] net837
+ vssd1 vssd1 vccd1 vccd1 _02882_ sky130_fd_sc_hd__mux2_1
XANTENNA__12498__A1 net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1132 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07862_ final_design.cpu.reg_window\[20\] final_design.cpu.reg_window\[52\] net868
+ vssd1 vssd1 vccd1 vccd1 _02813_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_3_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire526_X net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13906__RESET_B net1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09601_ _02705_ _04088_ net443 _02703_ vssd1 vssd1 vccd1 vccd1 _04520_ sky130_fd_sc_hd__o22a_1
XFILLER_0_78_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06813_ _01760_ _01761_ _01762_ _01763_ net778 net784 vssd1 vssd1 vccd1 vccd1 _01764_
+ sky130_fd_sc_hd__mux4_1
X_07793_ _02740_ _02741_ _02742_ _02743_ net684 net703 vssd1 vssd1 vccd1 vccd1 _02744_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__09115__A1 final_design.CPU_instr_adr\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09532_ _04429_ _04450_ vssd1 vssd1 vccd1 vccd1 _04451_ sky130_fd_sc_hd__and2_1
X_06744_ final_design.cpu.reg_window\[471\] final_design.cpu.reg_window\[503\] net929
+ vssd1 vssd1 vccd1 vccd1 _01695_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_1403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_1452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_1917 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08746__C _01598_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06675_ net884 _01619_ _01625_ _01612_ _01613_ vssd1 vssd1 vccd1 vccd1 _01626_ sky130_fd_sc_hd__a32oi_4
X_09463_ _02735_ _04281_ _02769_ vssd1 vssd1 vccd1 vccd1 _04382_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_56_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout253_A _04961_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08414_ _03361_ _03362_ _03363_ _03364_ net680 net700 vssd1 vssd1 vccd1 vccd1 _03365_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_59_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09394_ net494 _04312_ _04231_ vssd1 vssd1 vccd1 vccd1 _04313_ sky130_fd_sc_hd__a21o_1
XANTENNA__14035__CLK clknet_leaf_40_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08345_ _03103_ _03166_ _03231_ _03295_ vssd1 vssd1 vccd1 vccd1 _03296_ sky130_fd_sc_hd__and4_1
XANTENNA_fanout420_A net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_31_clk clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_31_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout1162_A net1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout518_A net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08276_ net611 _03224_ _03225_ net537 vssd1 vssd1 vccd1 vccd1 _03227_ sky130_fd_sc_hd__a211oi_2
X_07227_ final_design.cpu.reg_window\[840\] final_design.cpu.reg_window\[872\] net897
+ vssd1 vssd1 vccd1 vccd1 _02178_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14185__CLK clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout306_X net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07158_ final_design.cpu.reg_window\[10\] final_design.cpu.reg_window\[42\] net896
+ vssd1 vssd1 vccd1 vccd1 _02109_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_1_clk_X clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11933__B1 net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout887_A net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07089_ final_design.cpu.reg_window\[12\] final_design.cpu.reg_window\[44\] net895
+ vssd1 vssd1 vccd1 vccd1 _02040_ sky130_fd_sc_hd__mux2_1
XFILLER_0_41_1721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11187__Y _05897_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1107 net1116 vssd1 vssd1 vccd1 vccd1 net1107 sky130_fd_sc_hd__clkbuf_4
Xfanout1118 net100 vssd1 vssd1 vccd1 vccd1 net1118 sky130_fd_sc_hd__buf_2
Xfanout1129 net1131 vssd1 vssd1 vccd1 vccd1 net1129 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout675_X net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout186 net187 vssd1 vssd1 vccd1 vccd1 net186 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_22_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout197 net198 vssd1 vssd1 vccd1 vccd1 net197 sky130_fd_sc_hd__buf_2
XANTENNA_fanout842_X net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12810_ net1344 vssd1 vssd1 vccd1 vccd1 _00251_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13790_ clknet_leaf_13_clk _01021_ net1100 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[778\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12741_ final_design.VGA_adr\[3\] net796 _06380_ _05039_ vssd1 vssd1 vccd1 vccd1
+ _01350_ sky130_fd_sc_hd__a22o_1
XFILLER_0_6_1913 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_2925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12661__B2 final_design.data_from_mem\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_2302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06457__B net1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_2947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10672__B1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12672_ _06323_ net1420 net978 vssd1 vssd1 vccd1 vccd1 _01338_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11623_ net219 net630 vssd1 vssd1 vccd1 vccd1 _06169_ sky130_fd_sc_hd__and2_1
XANTENNA__11216__A2 net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_22_clk clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_22_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_13_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13402__CLK clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08672__B _01505_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_13_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10424__B1 _05195_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11554_ net220 net634 vssd1 vssd1 vccd1 vccd1 _06133_ sky130_fd_sc_hd__and2_1
XANTENNA__09290__B1 net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_59_2220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_2854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire543 _01966_ vssd1 vssd1 vccd1 vccd1 net543 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_59_2231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_2865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10505_ _05251_ _05253_ vssd1 vssd1 vccd1 vccd1 _05254_ sky130_fd_sc_hd__nand2_1
XFILLER_0_29_1318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_78_2876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11485_ net189 net2319 net308 vssd1 vssd1 vccd1 vccd1 _00364_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_74_2718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_74_2729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13224_ clknet_leaf_41_clk _00455_ net1220 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[212\]
+ sky130_fd_sc_hd__dfrtp_1
X_10436_ _03022_ net593 vssd1 vssd1 vccd1 vccd1 _05202_ sky130_fd_sc_hd__or2_1
XANTENNA__13552__CLK clknet_leaf_36_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11924__B1 net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11378__X _06065_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13155_ clknet_leaf_0_clk _00386_ net1061 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[143\]
+ sky130_fd_sc_hd__dfrtp_1
X_10367_ net9 net1023 net1006 final_design.data_from_mem\[16\] vssd1 vssd1 vccd1 vccd1
+ _00120_ sky130_fd_sc_hd__o22a_1
X_12106_ net1820 net214 net389 vssd1 vssd1 vccd1 vccd1 _00830_ sky130_fd_sc_hd__mux2_1
X_14215__1273 vssd1 vssd1 vccd1 vccd1 _14215__1273/HI net1273 sky130_fd_sc_hd__conb_1
X_10298_ final_design.VGA_data_control.data_to_VGA\[3\] final_design.VGA_data_control.data_to_VGA\[2\]
+ final_design.VGA_data_control.data_to_VGA\[1\] final_design.VGA_data_control.data_to_VGA\[0\]
+ final_design.VGA_data_control.h_count\[1\] net1049 vssd1 vssd1 vccd1 vccd1 _05152_
+ sky130_fd_sc_hd__mux4_1
X_13086_ clknet_leaf_13_clk _00317_ net1099 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[74\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10442__B net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08148__A2 _03096_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12037_ net1851 net216 net396 vssd1 vssd1 vccd1 vccd1 _00765_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07591__X _02542_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11554__A net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13988_ clknet_leaf_54_clk _01219_ net1178 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[976\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14058__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1002 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12939_ clknet_leaf_22_clk _00177_ net1163 vssd1 vssd1 vccd1 vccd1 net127 sky130_fd_sc_hd__dfrtp_1
XANTENNA__07470__C net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06460_ _01405_ _01412_ vssd1 vssd1 vccd1 vccd1 _00002_ sky130_fd_sc_hd__and2_1
XFILLER_0_69_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09959__A net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13082__CLK clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_13_clk clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_13_clk sky130_fd_sc_hd__clkbuf_8
X_08130_ final_design.cpu.reg_window\[141\] final_design.cpu.reg_window\[173\] net850
+ vssd1 vssd1 vccd1 vccd1 _03081_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12952__RESET_B net1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09281__A0 net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08061_ final_design.cpu.reg_window\[786\] final_design.cpu.reg_window\[818\] net845
+ vssd1 vssd1 vccd1 vccd1 _03012_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07012_ final_design.cpu.reg_window\[527\] final_design.cpu.reg_window\[559\] net890
+ vssd1 vssd1 vccd1 vccd1 _01963_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_1765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11915__B1 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1885 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkload38_A clknet_leaf_28_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12324__S net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11391__A1 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08963_ _03794_ _03901_ vssd1 vssd1 vccd1 vccd1 _03902_ sky130_fd_sc_hd__or2_1
XANTENNA__11448__B net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06493__S1 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07914_ _01722_ net617 vssd1 vssd1 vccd1 vccd1 _02865_ sky130_fd_sc_hd__nor2_1
X_08894_ _03664_ _03772_ vssd1 vssd1 vccd1 vccd1 _03840_ sky130_fd_sc_hd__xnor2_1
XANTENNA__11143__A1 _04939_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09887__A2 _04805_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12340__B1 net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1008_A _05170_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07845_ _02790_ _02795_ net712 vssd1 vssd1 vccd1 vccd1 _02796_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout370_A net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11694__A2 net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11464__A net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout468_A net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1861 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07776_ final_design.cpu.reg_window\[600\] final_design.cpu.reg_window\[632\] net862
+ vssd1 vssd1 vccd1 vccd1 _02727_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09639__A2 net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06558__A _01453_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07153__S net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09515_ net550 net549 net548 net546 net453 net463 vssd1 vssd1 vccd1 vccd1 _04434_
+ sky130_fd_sc_hd__mux4_1
X_06727_ final_design.cpu.reg_window\[792\] final_design.cpu.reg_window\[824\] net944
+ vssd1 vssd1 vccd1 vccd1 _01678_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12643__B2 final_design.data_from_mem\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout635_A _06123_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13425__CLK clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07745__S1 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09446_ net472 _04223_ vssd1 vssd1 vccd1 vccd1 _04365_ sky130_fd_sc_hd__or2_1
X_06658_ final_design.cpu.reg_window\[90\] final_design.cpu.reg_window\[122\] net941
+ vssd1 vssd1 vccd1 vccd1 _01609_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout423_X net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09377_ net453 _04223_ _04293_ vssd1 vssd1 vccd1 vccd1 _04296_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10808__A _05508_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06589_ _01535_ _01538_ vssd1 vssd1 vccd1 vccd1 _01540_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout1165_X net1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08328_ final_design.cpu.reg_window\[904\] final_design.cpu.reg_window\[936\] net816
+ vssd1 vssd1 vccd1 vccd1 _03279_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_23_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10957__A1 _04040_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13575__CLK clknet_leaf_62_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09811__A2 net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10957__B2 _04042_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08259_ final_design.cpu.reg_window\[138\] final_design.cpu.reg_window\[170\] net814
+ vssd1 vssd1 vccd1 vccd1 _03210_ sky130_fd_sc_hd__mux2_1
XANTENNA__09621__A_N _04342_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_1821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11270_ _01967_ net641 _05968_ _05969_ net658 vssd1 vssd1 vccd1 vccd1 _05970_ sky130_fd_sc_hd__a221o_2
XANTENNA_fanout792_X net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11906__A0 net196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10221_ net2441 _05099_ _05101_ vssd1 vssd1 vccd1 vccd1 _00035_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11382__A1 net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06740__B net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07328__S net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10152_ _01384_ _05048_ vssd1 vssd1 vccd1 vccd1 _05050_ sky130_fd_sc_hd__nor2_1
XFILLER_0_24_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06484__S1 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10083_ final_design.VGA_data_control.v_count\[8\] _04998_ _01404_ vssd1 vssd1 vccd1
+ vccd1 _04999_ sky130_fd_sc_hd__a21boi_2
Xhold9 final_design.cpu.reg_window\[31\] vssd1 vssd1 vccd1 vccd1 net1351 sky130_fd_sc_hd__dlygate4sd3_1
X_13911_ clknet_leaf_6_clk _01142_ net1128 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[899\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_67_2500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1636 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input29_A DAT_I[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_2511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08667__B _02061_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13842_ clknet_leaf_44_clk _01073_ net1209 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[830\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_1901 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13773_ clknet_leaf_48_clk _01004_ net1200 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[761\]
+ sky130_fd_sc_hd__dfrtp_1
X_10985_ _05690_ _05709_ vssd1 vssd1 vccd1 vccd1 _05712_ sky130_fd_sc_hd__nor2_1
XFILLER_0_74_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12724_ final_design.VGA_data_control.v_count\[1\] _06364_ vssd1 vssd1 vccd1 vccd1
+ _06365_ sky130_fd_sc_hd__nor2_1
XFILLER_0_6_1743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13918__CLK clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12655_ final_design.VGA_data_control.ready_data\[15\] net1020 net975 final_design.data_from_mem\[15\]
+ vssd1 vssd1 vccd1 vccd1 _06315_ sky130_fd_sc_hd__a22o_1
XANTENNA__12398__B1 net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11606_ net229 net631 vssd1 vssd1 vccd1 vccd1 _06160_ sky130_fd_sc_hd__and2_1
XFILLER_0_25_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12586_ net2555 net998 net984 final_design.data_from_mem\[4\] vssd1 vssd1 vccd1 vccd1
+ _01279_ sky130_fd_sc_hd__a22o_1
XFILLER_0_81_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11537_ net803 _02359_ net805 vssd1 vssd1 vccd1 vccd1 _06124_ sky130_fd_sc_hd__or3b_1
XFILLER_0_41_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold409 final_design.cpu.reg_window\[84\] vssd1 vssd1 vccd1 vccd1 net1751 sky130_fd_sc_hd__dlygate4sd3_1
X_11468_ net210 net640 vssd1 vssd1 vccd1 vccd1 _06106_ sky130_fd_sc_hd__and2_1
XFILLER_0_61_1905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13207_ clknet_leaf_6_clk _00438_ net1128 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[195\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09566__A1 net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10419_ _03224_ _05190_ vssd1 vssd1 vccd1 vccd1 _05193_ sky130_fd_sc_hd__nor2_1
X_14187_ net133 vssd1 vssd1 vccd1 vccd1 net170 sky130_fd_sc_hd__clkbuf_1
XANTENNA__12144__S net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06650__B _01599_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11399_ net663 _03781_ net738 vssd1 vssd1 vccd1 vccd1 _06083_ sky130_fd_sc_hd__a21oi_1
X_13138_ clknet_leaf_39_clk _00369_ net1209 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[126\]
+ sky130_fd_sc_hd__dfrtp_1
X_13069_ clknet_leaf_44_clk _00300_ net1202 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[57\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1109 final_design.cpu.reg_window\[370\] vssd1 vssd1 vccd1 vccd1 net2451 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_2_clk clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_2_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_75_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11676__A2 net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13151__RESET_B net1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13448__CLK clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07630_ final_design.cpu.reg_window\[412\] final_design.cpu.reg_window\[444\] net858
+ vssd1 vssd1 vccd1 vccd1 _02581_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07561_ net744 _01481_ vssd1 vssd1 vccd1 vccd1 _02512_ sky130_fd_sc_hd__nand2_2
XFILLER_0_53_1433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09300_ net494 _04112_ vssd1 vssd1 vccd1 vccd1 _04219_ sky130_fd_sc_hd__nor2_1
X_06512_ _01461_ _01462_ vssd1 vssd1 vccd1 vccd1 _01463_ sky130_fd_sc_hd__and2_2
X_07492_ net536 _02157_ _02439_ _02440_ _02187_ vssd1 vssd1 vccd1 vccd1 _02443_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_17_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09231_ _03388_ _03421_ _03389_ vssd1 vssd1 vccd1 vccd1 _04150_ sky130_fd_sc_hd__a21o_1
X_06443_ final_design.vga.v_current_state\[1\] final_design.vga.v_current_state\[0\]
+ vssd1 vssd1 vccd1 vccd1 _01397_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_17_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11731__B net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12319__S net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1190 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09162_ net614 _03550_ _01658_ _02423_ vssd1 vssd1 vccd1 vccd1 _04081_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_25_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10347__B net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07002__A net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08113_ _03058_ _03063_ net708 vssd1 vssd1 vccd1 vccd1 _03064_ sky130_fd_sc_hd__mux2_1
XANTENNA__06544__C _01480_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09093_ net619 _04014_ net255 vssd1 vssd1 vccd1 vccd1 _04017_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout216_A net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08044_ net618 _02991_ _02992_ _01850_ vssd1 vssd1 vccd1 vccd1 _02995_ sky130_fd_sc_hd__a211oi_2
Xhold910 final_design.cpu.reg_window\[111\] vssd1 vssd1 vccd1 vccd1 net2252 sky130_fd_sc_hd__dlygate4sd3_1
Xhold921 final_design.cpu.reg_window\[262\] vssd1 vssd1 vccd1 vccd1 net2263 sky130_fd_sc_hd__dlygate4sd3_1
Xhold932 final_design.cpu.reg_window\[410\] vssd1 vssd1 vccd1 vccd1 net2274 sky130_fd_sc_hd__dlygate4sd3_1
Xhold943 final_design.cpu.reg_window\[796\] vssd1 vssd1 vccd1 vccd1 net2285 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12054__S net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold954 final_design.cpu.reg_window\[511\] vssd1 vssd1 vccd1 vccd1 net2296 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1125_A net1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold965 final_design.cpu.reg_window\[430\] vssd1 vssd1 vccd1 vccd1 net2307 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12561__B1 net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold976 final_design.cpu.reg_window\[488\] vssd1 vssd1 vccd1 vccd1 net2318 sky130_fd_sc_hd__dlygate4sd3_1
Xhold987 final_design.cpu.reg_window\[667\] vssd1 vssd1 vccd1 vccd1 net2329 sky130_fd_sc_hd__dlygate4sd3_1
Xhold998 final_design.cpu.reg_window\[492\] vssd1 vssd1 vccd1 vccd1 net2340 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11178__B _05886_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09995_ net320 _04684_ _04781_ net318 _04913_ vssd1 vssd1 vccd1 vccd1 _04914_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_38_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout585_A net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11893__S net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08946_ _03886_ vssd1 vssd1 vccd1 vccd1 _03887_ sky130_fd_sc_hd__inv_2
XANTENNA__09871__B net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08877_ _03659_ _03774_ vssd1 vssd1 vccd1 vccd1 _03825_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout373_X net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout752_A _01427_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07828_ final_design.cpu.reg_window\[341\] final_design.cpu.reg_window\[373\] net858
+ vssd1 vssd1 vccd1 vccd1 _02779_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07759_ final_design.cpu.reg_window\[472\] final_design.cpu.reg_window\[504\] net864
+ vssd1 vssd1 vccd1 vccd1 _02710_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout540_X net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout638_X net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10770_ _05440_ _05501_ vssd1 vssd1 vccd1 vccd1 _05506_ sky130_fd_sc_hd__nor2_1
XFILLER_0_67_747 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11641__B net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09429_ _04225_ _04343_ _04339_ vssd1 vssd1 vccd1 vccd1 _04348_ sky130_fd_sc_hd__o21a_1
XFILLER_0_54_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout805_X net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14214__1272 vssd1 vssd1 vccd1 vccd1 _14214__1272/HI net1272 sky130_fd_sc_hd__conb_1
X_12440_ net1625 net221 net334 vssd1 vssd1 vccd1 vccd1 _01147_ sky130_fd_sc_hd__mux2_1
XANTENNA__09886__X _04805_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08143__S1 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12371_ net1844 net244 net268 vssd1 vssd1 vccd1 vccd1 _01082_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14110_ clknet_leaf_14_clk _01307_ net1110 vssd1 vssd1 vccd1 vccd1 final_design.reqhand.data_from_UART\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07847__A _01788_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11322_ _04597_ _06015_ net652 vssd1 vssd1 vccd1 vccd1 _06016_ sky130_fd_sc_hd__mux2_2
XFILLER_0_22_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14229__1283 vssd1 vssd1 vccd1 vccd1 _14229__1283/HI net1283 sky130_fd_sc_hd__conb_1
XANTENNA__09548__A1 net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14041_ clknet_leaf_15_clk _00033_ net1095 vssd1 vssd1 vccd1 vccd1 final_design.uart.BAUD_counter\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09548__B2 net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11253_ net736 _03950_ vssd1 vssd1 vccd1 vccd1 _05955_ sky130_fd_sc_hd__nand2_1
XANTENNA__12552__B1 net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1072 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10204_ final_design.uart.BAUD_counter\[1\] final_design.uart.BAUD_counter\[0\] vssd1
+ vssd1 vccd1 vccd1 _05091_ sky130_fd_sc_hd__nand2_1
X_11184_ final_design.reqhand.data_from_UART\[5\] final_design.data_from_mem\[5\]
+ net247 vssd1 vssd1 vccd1 vccd1 _05894_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_1709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10135_ final_design.VGA_data_control.state\[1\] _01402_ _05038_ final_design.VGA_data_control.state\[0\]
+ vssd1 vssd1 vccd1 vccd1 _05039_ sky130_fd_sc_hd__and4b_1
XANTENNA__08678__A _03617_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07582__A net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10066_ _04550_ _04551_ vssd1 vssd1 vccd1 vccd1 _04985_ sky130_fd_sc_hd__nand2_1
XANTENNA__11658__A2 net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13825_ clknet_leaf_47_clk _01056_ net1203 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[813\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13740__CLK clknet_leaf_46_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12607__B2 final_design.data_from_mem\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08684__Y _03635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07709__S1 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13756_ clknet_leaf_2_clk _00987_ net1065 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[744\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_50_1606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10968_ net1474 net1033 _05694_ _05695_ vssd1 vssd1 vccd1 vccd1 _00197_ sky130_fd_sc_hd__a22o_1
XFILLER_0_35_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12707_ _01391_ _06338_ _06343_ _06346_ vssd1 vssd1 vccd1 vccd1 _06348_ sky130_fd_sc_hd__o31ai_2
XANTENNA__09302__A net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08382__S1 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06837__A2 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11291__B1 _05843_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10448__A _02731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12139__S net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13687_ clknet_leaf_4_clk _00918_ net1084 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[675\]
+ sky130_fd_sc_hd__dfrtp_1
X_10899_ _05593_ _05612_ _05628_ vssd1 vssd1 vccd1 vccd1 _05629_ sky130_fd_sc_hd__a21o_1
XFILLER_0_13_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08039__A1 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13890__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12638_ _06306_ net1439 net980 vssd1 vssd1 vccd1 vccd1 _01321_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12795__26 clknet_leaf_31_clk vssd1 vssd1 vccd1 vccd1 net1336 sky130_fd_sc_hd__inv_2
XFILLER_0_31_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12569_ net2259 _06289_ _06286_ vssd1 vssd1 vccd1 vccd1 _01269_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06661__A net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold206 final_design.cpu.reg_window\[707\] vssd1 vssd1 vccd1 vccd1 net1548 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_1568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07893__S0 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold217 final_design.cpu.reg_window\[223\] vssd1 vssd1 vccd1 vccd1 net1559 sky130_fd_sc_hd__dlygate4sd3_1
Xhold228 final_design.cpu.reg_window\[688\] vssd1 vssd1 vccd1 vccd1 net1570 sky130_fd_sc_hd__dlygate4sd3_1
X_14239_ net1293 vssd1 vssd1 vccd1 vccd1 gpio_out[17] sky130_fd_sc_hd__buf_2
Xhold239 final_design.cpu.reg_window\[675\] vssd1 vssd1 vccd1 vccd1 net1581 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_1844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_894 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12543__B1 net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08211__A1 net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout708 net709 vssd1 vssd1 vccd1 vccd1 net708 sky130_fd_sc_hd__clkbuf_2
Xfanout719 net720 vssd1 vssd1 vccd1 vccd1 net719 sky130_fd_sc_hd__clkbuf_4
X_08800_ _03675_ _03676_ _03749_ _03673_ vssd1 vssd1 vccd1 vccd1 _03751_ sky130_fd_sc_hd__o31ai_2
XANTENNA_clkbuf_leaf_41_clk_X clknet_leaf_41_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13270__CLK clknet_leaf_57_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09780_ _04187_ _04698_ vssd1 vssd1 vccd1 vccd1 _04699_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_7_Right_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06992_ final_design.cpu.reg_window\[335\] final_design.cpu.reg_window\[367\] net901
+ vssd1 vssd1 vccd1 vccd1 _01943_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_33_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12838__CLK clknet_leaf_18_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08731_ final_design.CPU_instr_adr\[14\] _02000_ vssd1 vssd1 vccd1 vccd1 _03682_
+ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_33_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08662_ _01998_ _02029_ _02062_ vssd1 vssd1 vccd1 vccd1 _03613_ sky130_fd_sc_hd__or3_2
XANTENNA__07846__A1_N net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10321__A2 net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_56_clk_X clknet_leaf_56_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07613_ final_design.cpu.reg_window\[861\] final_design.cpu.reg_window\[893\] net870
+ vssd1 vssd1 vccd1 vccd1 _02564_ sky130_fd_sc_hd__mux2_1
X_08593_ final_design.cpu.reg_window\[640\] final_design.cpu.reg_window\[672\] net826
+ vssd1 vssd1 vccd1 vccd1 _03544_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07544_ net753 _02494_ vssd1 vssd1 vccd1 vccd1 _02495_ sky130_fd_sc_hd__or2_2
XFILLER_0_72_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12074__A2 _05952_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_822 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_27_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09570__S0 net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12049__S net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07475_ _02419_ _02424_ vssd1 vssd1 vccd1 vccd1 _02426_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout333_A _06283_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06555__B _01505_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09214_ _02803_ _02836_ _04128_ _04132_ vssd1 vssd1 vccd1 vccd1 _04133_ sky130_fd_sc_hd__a31oi_2
X_06426_ final_design.data_from_mem\[20\] vssd1 vssd1 vccd1 vccd1 _01381_ sky130_fd_sc_hd__inv_2
XFILLER_0_63_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11888__S net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09145_ net528 net456 _04063_ vssd1 vssd1 vccd1 vccd1 _04064_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout500_A net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1624 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1242_A net1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout219_X net219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11585__A1 net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11386__A2_N _06071_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_12_Left_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09076_ final_design.CPU_instr_adr\[6\] _03785_ vssd1 vssd1 vccd1 vccd1 _04002_ sky130_fd_sc_hd__xor2_1
XANTENNA__08262__S net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1668 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06461__A0 net1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08027_ net717 _02977_ vssd1 vssd1 vccd1 vccd1 _02978_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_9_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1030_X net1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold740 final_design.cpu.reg_window\[282\] vssd1 vssd1 vccd1 vccd1 net2082 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13613__CLK clknet_leaf_48_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold751 final_design.cpu.reg_window\[362\] vssd1 vssd1 vccd1 vccd1 net2093 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11337__A1 _01722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12534__B1 net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold762 final_design.cpu.reg_window\[814\] vssd1 vssd1 vccd1 vccd1 net2104 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11337__B2 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold773 final_design.cpu.reg_window\[260\] vssd1 vssd1 vccd1 vccd1 net2115 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12792__23_A clknet_leaf_27_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold784 final_design.cpu.reg_window\[143\] vssd1 vssd1 vccd1 vccd1 net2126 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout490_X net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold795 final_design.cpu.reg_window\[472\] vssd1 vssd1 vccd1 vccd1 net2137 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout588_X net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08753__A2 _01659_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09978_ _03327_ _04895_ _04046_ vssd1 vssd1 vccd1 vccd1 _04897_ sky130_fd_sc_hd__o21a_1
XFILLER_0_60_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13002__RESET_B net1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08929_ final_design.CPU_instr_adr\[23\] net1014 _03867_ _03871_ vssd1 vssd1 vccd1
+ vccd1 _00234_ sky130_fd_sc_hd__a22o_1
XANTENNA__13763__CLK clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout755_X net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08505__A2 _03450_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11940_ _06141_ net287 net410 net1905 vssd1 vssd1 vccd1 vccd1 _00675_ sky130_fd_sc_hd__a22o_1
XFILLER_0_19_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_1748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11871_ net432 net195 net554 net518 net1606 vssd1 vssd1 vccd1 vccd1 _00617_ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout922_X net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14119__CLK clknet_leaf_17_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13610_ clknet_leaf_60_clk _00841_ net1168 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[598\]
+ sky130_fd_sc_hd__dfrtp_1
X_10822_ net966 _05555_ vssd1 vssd1 vccd1 vccd1 _05556_ sky130_fd_sc_hd__nand2_1
XANTENNA__12065__A2 net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09466__B1 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10076__A1 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13541_ clknet_leaf_50_clk _00772_ net1172 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[529\]
+ sky130_fd_sc_hd__dfrtp_1
X_10753_ _05484_ _05488_ vssd1 vssd1 vccd1 vccd1 _05490_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_3_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input96_A memory_size[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13472_ clknet_leaf_11_clk _00703_ net1097 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[460\]
+ sky130_fd_sc_hd__dfrtp_1
X_10684_ net253 _04654_ vssd1 vssd1 vccd1 vccd1 _05424_ sky130_fd_sc_hd__and2b_1
XANTENNA__13143__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12423_ _06245_ _06264_ net340 net2015 vssd1 vssd1 vccd1 vccd1 _01132_ sky130_fd_sc_hd__a22o_1
XANTENNA__09313__S0 net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10379__A2 net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08680__B net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12354_ net2409 net362 net352 _06032_ vssd1 vssd1 vccd1 vccd1 _01066_ sky130_fd_sc_hd__a22o_1
X_11305_ _01853_ net641 _05999_ _06000_ net656 vssd1 vssd1 vccd1 vccd1 _06001_ sky130_fd_sc_hd__a221o_4
XANTENNA__13293__CLK clknet_leaf_44_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12285_ net586 _06215_ net513 net371 net2314 vssd1 vssd1 vccd1 vccd1 _01000_ sky130_fd_sc_hd__a32o_1
XANTENNA__11328__A1 final_design.data_from_mem\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12525__B1 net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14024_ clknet_leaf_41_clk _01255_ net1224 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[1012\]
+ sky130_fd_sc_hd__dfrtp_1
X_11236_ _04676_ net655 vssd1 vssd1 vccd1 vccd1 _05940_ sky130_fd_sc_hd__nand2_1
XANTENNA__11879__A2 net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11167_ net731 _04022_ _05878_ vssd1 vssd1 vccd1 vccd1 _05879_ sky130_fd_sc_hd__o21ai_1
X_10118_ _05003_ _05027_ _05028_ vssd1 vssd1 vccd1 vccd1 final_design.vga.v_next_count\[5\]
+ sky130_fd_sc_hd__and3_1
XANTENNA__11546__B net240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11098_ _04177_ net253 _04990_ vssd1 vssd1 vccd1 vccd1 _05819_ sky130_fd_sc_hd__o21ai_1
XANTENNA__10450__B net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06850__S1 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10049_ _04452_ _04454_ vssd1 vssd1 vccd1 vccd1 _04968_ sky130_fd_sc_hd__xnor2_1
XANTENNA__08052__S0 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11265__C net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_19_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11562__A net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09303__Y _04222_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13808_ clknet_leaf_34_clk _01039_ net1239 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[796\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07251__S net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11264__B1 net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13739_ clknet_leaf_53_clk _00970_ net1187 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[727\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11803__A2 net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07260_ _02193_ _02199_ _02210_ net881 vssd1 vssd1 vccd1 vccd1 _02211_ sky130_fd_sc_hd__a22oi_4
XTAP_TAPCELL_ROW_41_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08107__S1 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07191_ net749 _02135_ net745 vssd1 vssd1 vccd1 vccd1 _02142_ sky130_fd_sc_hd__o21a_1
XANTENNA__13636__CLK clknet_leaf_54_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10625__B final_design.VGA_adr\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12788__19_A clknet_leaf_30_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12516__B1 net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09901_ _04124_ _04812_ _04813_ vssd1 vssd1 vccd1 vccd1 _04820_ sky130_fd_sc_hd__or3_1
XFILLER_0_22_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_35_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkload20_A clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13786__CLK clknet_leaf_58_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout505 net516 vssd1 vssd1 vccd1 vccd1 net505 sky130_fd_sc_hd__clkbuf_4
Xfanout516 _06259_ vssd1 vssd1 vccd1 vccd1 net516 sky130_fd_sc_hd__buf_4
X_09832_ net69 _04182_ vssd1 vssd1 vccd1 vccd1 _04751_ sky130_fd_sc_hd__xnor2_1
Xfanout527 _02502_ vssd1 vssd1 vccd1 vccd1 net527 sky130_fd_sc_hd__buf_4
Xfanout538 _02091_ vssd1 vssd1 vccd1 vccd1 net538 sky130_fd_sc_hd__buf_2
Xfanout549 _01815_ vssd1 vssd1 vccd1 vccd1 net549 sky130_fd_sc_hd__clkbuf_4
X_14213__1271 vssd1 vssd1 vccd1 vccd1 _14213__1271/HI net1271 sky130_fd_sc_hd__conb_1
XANTENNA__07426__S net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11456__B net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09763_ _03585_ _03589_ vssd1 vssd1 vccd1 vccd1 _04682_ sky130_fd_sc_hd__nand2_1
X_06975_ final_design.cpu.reg_window\[784\] final_design.cpu.reg_window\[816\] net923
+ vssd1 vssd1 vccd1 vccd1 _01926_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout283_A net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_21_clk_A clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13016__CLK clknet_leaf_62_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08714_ final_design.CPU_instr_adr\[25\] _01660_ vssd1 vssd1 vccd1 vccd1 _03665_
+ sky130_fd_sc_hd__nor2_1
X_09694_ net447 _04600_ _04610_ _04612_ vssd1 vssd1 vccd1 vccd1 _04613_ sky130_fd_sc_hd__o22a_2
XANTENNA__08499__B2 net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09160__A2 net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08645_ _02772_ _03593_ vssd1 vssd1 vccd1 vccd1 _03596_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_1_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout450_A _04069_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1192_A net1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout548_A _01850_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06837__Y _01788_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14228__1282 vssd1 vssd1 vccd1 vccd1 _14228__1282/HI net1282 sky130_fd_sc_hd__conb_1
X_08576_ final_design.cpu.reg_window\[448\] final_design.cpu.reg_window\[480\] net827
+ vssd1 vssd1 vccd1 vccd1 _03527_ sky130_fd_sc_hd__mux2_1
XANTENNA__13166__CLK clknet_leaf_45_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_36_clk_A clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10058__A1 _04529_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07527_ final_design.cpu.reg_window\[351\] final_design.cpu.reg_window\[383\] net939
+ vssd1 vssd1 vccd1 vccd1 _02478_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout336_X net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07458_ final_design.cpu.reg_window\[768\] final_design.cpu.reg_window\[800\] net909
+ vssd1 vssd1 vccd1 vccd1 _02409_ sky130_fd_sc_hd__mux2_1
X_06409_ final_design.CPU_instr_adr\[14\] vssd1 vssd1 vccd1 vccd1 _01364_ sky130_fd_sc_hd__inv_2
XFILLER_0_49_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07389_ final_design.cpu.reg_window\[194\] final_design.cpu.reg_window\[226\] net913
+ vssd1 vssd1 vccd1 vccd1 _02340_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout503_X net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1245_X net1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11411__S net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09128_ net659 _04045_ vssd1 vssd1 vccd1 vccd1 _04047_ sky130_fd_sc_hd__nand2_2
X_09059_ _03787_ _03986_ vssd1 vssd1 vccd1 vccd1 _03987_ sky130_fd_sc_hd__or2_1
XFILLER_0_66_1487 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12507__B1 net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12070_ net2295 net392 net498 _05922_ vssd1 vssd1 vccd1 vccd1 _00795_ sky130_fd_sc_hd__a22o_1
Xhold570 final_design.cpu.reg_window\[76\] vssd1 vssd1 vccd1 vccd1 net1912 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout872_X net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold581 final_design.cpu.reg_window\[581\] vssd1 vssd1 vccd1 vccd1 net1923 sky130_fd_sc_hd__dlygate4sd3_1
Xhold592 final_design.cpu.reg_window\[666\] vssd1 vssd1 vccd1 vccd1 net1934 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08499__Y _03450_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11021_ net966 _05743_ _05745_ vssd1 vssd1 vccd1 vccd1 _05746_ sky130_fd_sc_hd__o21a_1
XANTENNA__09923__A1 _04109_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11647__A net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09923__B2 _04222_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_2584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11730__A1 net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_2595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08021__A net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07563__C net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09687__A0 net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12972_ net1311 _00209_ net1166 vssd1 vssd1 vccd1 vccd1 final_design.CPU_instr_adr\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA_input11_A DAT_I[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13509__CLK clknet_leaf_49_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07860__A net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11923_ _06126_ net282 net409 net2485 vssd1 vssd1 vccd1 vccd1 _00660_ sky130_fd_sc_hd__a22o_1
XANTENNA__07162__A1 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09123__Y _04042_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11854_ _06104_ net277 net517 net1897 vssd1 vssd1 vccd1 vccd1 _00604_ sky130_fd_sc_hd__a22o_1
XFILLER_0_55_1870 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07071__S net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14091__CLK clknet_leaf_19_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_2377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10805_ net44 _05539_ vssd1 vssd1 vccd1 vccd1 _05540_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_64_2388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_1865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_64_2399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11785_ net2480 net412 _06232_ net429 vssd1 vssd1 vccd1 vccd1 _00542_ sky130_fd_sc_hd__a22o_1
XFILLER_0_32_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11797__B2 net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13524_ clknet_leaf_10_clk _00755_ net1102 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[512\]
+ sky130_fd_sc_hd__dfrtp_1
X_10736_ net964 _05473_ vssd1 vssd1 vccd1 vccd1 _05474_ sky130_fd_sc_hd__nand2_1
X_13455_ clknet_leaf_42_clk _00686_ net1224 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[443\]
+ sky130_fd_sc_hd__dfrtp_1
X_10667_ net69 final_design.VGA_adr\[8\] _05407_ vssd1 vssd1 vccd1 vccd1 _05408_ sky130_fd_sc_hd__and3_1
XANTENNA__11549__A1 net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12406_ _06104_ net343 net338 net2100 vssd1 vssd1 vccd1 vccd1 _01116_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_11_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13386_ clknet_leaf_51_clk _00617_ net1170 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[374\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10598_ _05330_ _05342_ net65 vssd1 vssd1 vccd1 vccd1 _05343_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_11_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07100__A net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput108 net108 vssd1 vssd1 vccd1 vccd1 ADR_O[16] sky130_fd_sc_hd__clkbuf_4
X_12337_ net2534 net360 net346 _05905_ vssd1 vssd1 vccd1 vccd1 _01049_ sky130_fd_sc_hd__a22o_1
XANTENNA__07622__C1 _01535_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput119 net119 vssd1 vssd1 vccd1 vccd1 ADR_O[26] sky130_fd_sc_hd__clkbuf_4
XANTENNA__07594__X _02545_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12268_ net563 _06198_ net505 net369 net2164 vssd1 vssd1 vccd1 vccd1 _00983_ sky130_fd_sc_hd__a32o_1
XFILLER_0_43_1251 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14007_ clknet_leaf_6_clk _01238_ net1129 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[995\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13039__CLK clknet_leaf_42_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11219_ final_design.data_from_mem\[9\] _05914_ _05917_ vssd1 vssd1 vccd1 vccd1 _05925_
+ sky130_fd_sc_hd__a21o_1
XANTENNA__12152__S net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12199_ net566 _06127_ net506 net377 net1964 vssd1 vssd1 vccd1 vccd1 _00917_ sky130_fd_sc_hd__a32o_1
XANTENNA__07246__S net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11991__S net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06760_ final_design.cpu.reg_window\[727\] final_design.cpu.reg_window\[759\] net929
+ vssd1 vssd1 vccd1 vccd1 _01711_ sky130_fd_sc_hd__mux2_1
XANTENNA__13189__CLK clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09314__X _04233_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09142__A2 _03549_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06691_ _01638_ _01639_ _01640_ _01641_ net774 net792 vssd1 vssd1 vccd1 vccd1 _01642_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_76_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11292__A net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08430_ final_design.cpu.reg_window\[517\] final_design.cpu.reg_window\[549\] net843
+ vssd1 vssd1 vccd1 vccd1 _03381_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06900__A1 _01468_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08361_ final_design.cpu.reg_window\[967\] final_design.cpu.reg_window\[999\] net811
+ vssd1 vssd1 vccd1 vccd1 _03312_ sky130_fd_sc_hd__mux2_1
XANTENNA__08102__B1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07312_ final_design.cpu.reg_window\[645\] final_design.cpu.reg_window\[677\] net921
+ vssd1 vssd1 vccd1 vccd1 _02263_ sky130_fd_sc_hd__mux2_1
XANTENNA__09697__A net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08292_ _03239_ _03240_ _03241_ _03242_ net674 net696 vssd1 vssd1 vccd1 vccd1 _03243_
+ sky130_fd_sc_hd__mux4_1
X_07243_ final_design.cpu.reg_window\[327\] final_design.cpu.reg_window\[359\] net900
+ vssd1 vssd1 vccd1 vccd1 _02194_ sky130_fd_sc_hd__mux2_1
XANTENNA__12327__S net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07174_ net757 _02124_ vssd1 vssd1 vccd1 vccd1 _02125_ sky130_fd_sc_hd__or2_1
XANTENNA__07839__S0 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12201__A2 net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_1785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1038_A _01410_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout302 net303 vssd1 vssd1 vccd1 vccd1 net302 sky130_fd_sc_hd__buf_4
XANTENNA_fanout498_A net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout313 _06092_ vssd1 vssd1 vccd1 vccd1 net313 sky130_fd_sc_hd__buf_4
XANTENNA__12062__S net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout324 net325 vssd1 vssd1 vccd1 vccd1 net324 sky130_fd_sc_hd__buf_4
XFILLER_0_61_1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11712__A1 net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout335 net337 vssd1 vssd1 vccd1 vccd1 net335 sky130_fd_sc_hd__clkbuf_8
Xfanout346 net347 vssd1 vssd1 vccd1 vccd1 net346 sky130_fd_sc_hd__clkbuf_4
XANTENNA_input3_A DAT_I[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09815_ net482 _04733_ _04112_ vssd1 vssd1 vccd1 vccd1 _04734_ sky130_fd_sc_hd__a21o_1
Xfanout357 net358 vssd1 vssd1 vccd1 vccd1 net357 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09381__A2 net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout368 net369 vssd1 vssd1 vccd1 vccd1 net368 sky130_fd_sc_hd__buf_4
Xfanout379 _06271_ vssd1 vssd1 vccd1 vccd1 net379 sky130_fd_sc_hd__buf_4
XANTENNA_fanout286_X net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout665_A _01503_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09746_ net491 _04559_ _04341_ vssd1 vssd1 vccd1 vccd1 _04665_ sky130_fd_sc_hd__a21o_1
XFILLER_0_74_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06958_ net784 net664 _01821_ vssd1 vssd1 vccd1 vccd1 _01909_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_69_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11914__B _05845_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1745 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09677_ _02803_ _02834_ _04330_ net449 vssd1 vssd1 vccd1 vccd1 _04596_ sky130_fd_sc_hd__a31o_1
X_06889_ final_design.cpu.reg_window\[979\] final_design.cpu.reg_window\[1011\] net911
+ vssd1 vssd1 vccd1 vccd1 _01840_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout453_X net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1195_X net1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08628_ _02026_ _03072_ _03097_ vssd1 vssd1 vccd1 vccd1 _03579_ sky130_fd_sc_hd__and3b_1
XFILLER_0_74_1789 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13801__CLK clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08559_ final_design.cpu.reg_window\[513\] final_design.cpu.reg_window\[545\] net831
+ vssd1 vssd1 vccd1 vccd1 _03510_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout620_X net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout718_X net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11930__A net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11779__B2 _05911_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11570_ net223 net637 vssd1 vssd1 vccd1 vccd1 _06141_ sky130_fd_sc_hd__and2_1
XFILLER_0_0_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10521_ _04847_ net250 vssd1 vssd1 vccd1 vccd1 _05269_ sky130_fd_sc_hd__nor2_1
XANTENNA__13951__CLK clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1749 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11141__S net245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13240_ clknet_leaf_62_clk _00471_ net1073 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[228\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_33_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10452_ _02698_ net593 vssd1 vssd1 vccd1 vccd1 _05210_ sky130_fd_sc_hd__nor2_1
XFILLER_0_66_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1705 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11844__C_N net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13171_ clknet_leaf_37_clk _00402_ net1206 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[159\]
+ sky130_fd_sc_hd__dfrtp_1
X_10383_ _01372_ _04995_ vssd1 vssd1 vccd1 vccd1 _05172_ sky130_fd_sc_hd__nand2_4
XFILLER_0_81_1749 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06958__A1 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_2793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_2170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12122_ net1733 net184 net390 vssd1 vssd1 vccd1 vccd1 _00846_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_53_2012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_2023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input59_A mem_adr_start[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_2657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_2034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12053_ net2127 net187 net398 vssd1 vssd1 vccd1 vccd1 _00781_ sky130_fd_sc_hd__mux2_1
XFILLER_0_40_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07066__S net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11004_ net54 _05728_ vssd1 vssd1 vccd1 vccd1 _05730_ sky130_fd_sc_hd__nor2_1
XANTENNA__13331__CLK clknet_leaf_40_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1891 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout891 net892 vssd1 vssd1 vccd1 vccd1 net891 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_5_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08686__A _02325_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_3_6_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_3_6_0_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_5_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07590__A _02504_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11467__A0 net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input14_X net14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12955_ clknet_leaf_29_clk _00193_ net1195 vssd1 vssd1 vccd1 vccd1 net113 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06569__S0 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13481__CLK clknet_leaf_36_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11906_ net196 net2324 net274 vssd1 vssd1 vccd1 vccd1 _00648_ sky130_fd_sc_hd__mux2_1
X_12886_ clknet_leaf_17_clk _00124_ net1109 vssd1 vssd1 vccd1 vccd1 final_design.data_from_mem\[20\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__07686__A2 _02635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11837_ net186 net1816 net267 vssd1 vssd1 vccd1 vccd1 _00589_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07589__X _02540_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08635__A1 net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11768_ net673 _05850_ _06118_ vssd1 vssd1 vccd1 vccd1 _06227_ sky130_fd_sc_hd__or3_1
X_14212__1270 vssd1 vssd1 vccd1 vccd1 _14212__1270/HI net1270 sky130_fd_sc_hd__conb_1
X_10719_ _05438_ _05441_ _05457_ vssd1 vssd1 vccd1 vccd1 _05458_ sky130_fd_sc_hd__nand3_1
X_13507_ clknet_leaf_1_clk _00738_ net1071 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[495\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12147__S net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11699_ net207 net626 vssd1 vssd1 vccd1 vccd1 _06208_ sky130_fd_sc_hd__and2_1
XANTENNA__10456__A _02602_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13438_ clknet_leaf_9_clk _00669_ net1097 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[426\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12195__A1 net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13369_ clknet_leaf_55_clk _00600_ net1148 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[357\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14227__1281 vssd1 vssd1 vccd1 vccd1 _14227__1281/HI net1281 sky130_fd_sc_hd__conb_1
XFILLER_0_80_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07930_ net718 _02880_ vssd1 vssd1 vccd1 vccd1 _02881_ sky130_fd_sc_hd__nor2_1
XFILLER_0_48_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12498__A2 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07861_ final_design.cpu.reg_window\[84\] final_design.cpu.reg_window\[116\] net868
+ vssd1 vssd1 vccd1 vccd1 _02812_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07374__A1 net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09600_ net473 _04211_ _04518_ _04109_ vssd1 vssd1 vccd1 vccd1 _04519_ sky130_fd_sc_hd__a211o_1
XFILLER_0_58_1718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06812_ final_design.cpu.reg_window\[21\] final_design.cpu.reg_window\[53\] net939
+ vssd1 vssd1 vccd1 vccd1 _01763_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07792_ final_design.cpu.reg_window\[409\] final_design.cpu.reg_window\[441\] net854
+ vssd1 vssd1 vccd1 vccd1 _02743_ sky130_fd_sc_hd__mux2_1
XANTENNA__13824__CLK clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1019 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09531_ net321 _04430_ _04431_ _04449_ vssd1 vssd1 vccd1 vccd1 _04450_ sky130_fd_sc_hd__o31ai_2
X_06743_ final_design.cpu.reg_window\[279\] final_design.cpu.reg_window\[311\] net931
+ vssd1 vssd1 vccd1 vccd1 _01694_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09462_ _04048_ _04360_ _04361_ _04380_ vssd1 vssd1 vccd1 vccd1 _04381_ sky130_fd_sc_hd__a31o_1
X_06674_ net761 _01624_ vssd1 vssd1 vccd1 vccd1 _01625_ sky130_fd_sc_hd__or2_1
X_08413_ final_design.cpu.reg_window\[389\] final_design.cpu.reg_window\[421\] net838
+ vssd1 vssd1 vccd1 vccd1 _03364_ sky130_fd_sc_hd__mux2_1
XANTENNA__13974__CLK clknet_leaf_59_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09393_ _04227_ _04295_ vssd1 vssd1 vccd1 vccd1 _04312_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout246_A net247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09418__A3 net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1041 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08344_ _03259_ _03260_ _03290_ _03292_ vssd1 vssd1 vccd1 vccd1 _03295_ sky130_fd_sc_hd__o22a_1
XFILLER_0_58_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12422__A2 net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10433__B2 net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12057__S net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11630__B1 net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08275_ net599 _03224_ _03200_ vssd1 vssd1 vccd1 vccd1 _03226_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout413_A net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1155_A net1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07226_ net757 _02176_ vssd1 vssd1 vccd1 vccd1 _02177_ sky130_fd_sc_hd__or2_1
XFILLER_0_67_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12186__A1 net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11896__S net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07157_ final_design.cpu.reg_window\[74\] final_design.cpu.reg_window\[106\] net898
+ vssd1 vssd1 vccd1 vccd1 _02108_ sky130_fd_sc_hd__mux2_1
XANTENNA__09051__A1 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08485__S0 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13354__CLK clknet_leaf_51_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11909__B _05845_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07088_ final_design.cpu.reg_window\[76\] final_design.cpu.reg_window\[108\] net895
+ vssd1 vssd1 vccd1 vccd1 _02039_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_1599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout782_A _01419_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1108 net1109 vssd1 vssd1 vccd1 vccd1 net1108 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_11_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12489__A2 net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1119 net1127 vssd1 vssd1 vccd1 vccd1 net1119 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout668_X net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout176 _06089_ vssd1 vssd1 vccd1 vccd1 net176 sky130_fd_sc_hd__buf_2
Xfanout187 _06052_ vssd1 vssd1 vccd1 vccd1 net187 sky130_fd_sc_hd__buf_2
Xfanout198 _06010_ vssd1 vssd1 vccd1 vccd1 net198 sky130_fd_sc_hd__buf_2
XANTENNA__11449__A0 net242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07614__S net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09729_ _03071_ net446 net438 _03068_ _04640_ vssd1 vssd1 vccd1 vccd1 _04648_ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout835_X net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06738__B net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12740_ _06366_ _06377_ vssd1 vssd1 vccd1 vccd1 _06380_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_39_1695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_61_2303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06457__C net34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_2937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12671_ final_design.VGA_data_control.ready_data\[23\] net1019 net974 final_design.data_from_mem\[23\]
+ vssd1 vssd1 vccd1 vccd1 _06323_ sky130_fd_sc_hd__a22o_1
XFILLER_0_77_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06971__S0 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11622_ net559 net420 _06168_ net298 net1884 vssd1 vssd1 vccd1 vccd1 _00443_ sky130_fd_sc_hd__a32o_1
XANTENNA__09814__A0 _04618_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12413__A2 net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08672__C _01537_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1879 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11553_ net2194 net302 _06132_ net420 vssd1 vssd1 vccd1 vccd1 _00410_ sky130_fd_sc_hd__a22o_1
XANTENNA__10424__B2 net245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_2210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10504_ net93 final_design.VGA_adr\[1\] vssd1 vssd1 vccd1 vccd1 _05253_ sky130_fd_sc_hd__or2_1
XFILLER_0_29_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_59_2221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_2855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_2232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_2866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11484_ net190 net2444 net308 vssd1 vssd1 vccd1 vccd1 _00363_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_78_2877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_2719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13223_ clknet_leaf_62_clk _00454_ net1120 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[211\]
+ sky130_fd_sc_hd__dfrtp_1
X_10435_ net1461 net1028 _05201_ net246 vssd1 vssd1 vccd1 vccd1 _00158_ sky130_fd_sc_hd__a22o_1
X_13154_ clknet_leaf_11_clk _00385_ net1086 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[142\]
+ sky130_fd_sc_hd__dfrtp_1
X_10366_ net8 net1023 net1007 final_design.data_from_mem\[15\] vssd1 vssd1 vccd1 vccd1
+ _00119_ sky130_fd_sc_hd__o22a_1
X_12105_ net1971 net216 net388 vssd1 vssd1 vccd1 vccd1 _00829_ sky130_fd_sc_hd__mux2_1
X_13085_ clknet_leaf_2_clk _00316_ net1064 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[73\]
+ sky130_fd_sc_hd__dfrtp_1
X_10297_ final_design.VGA_data_control.data_to_VGA\[4\] _05013_ _05150_ final_design.VGA_data_control.h_count\[3\]
+ vssd1 vssd1 vccd1 vccd1 _05151_ sky130_fd_sc_hd__a211o_1
XANTENNA__13847__CLK clknet_leaf_58_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_0_Left_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_1806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12036_ net2184 net218 net396 vssd1 vssd1 vccd1 vccd1 _00764_ sky130_fd_sc_hd__mux2_1
XANTENNA__11688__B1 net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11394__X _06079_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10360__B1 net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09305__A _02503_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12871__CLK clknet_leaf_25_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13997__CLK clknet_leaf_44_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11554__B net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07108__A1 net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13987_ clknet_leaf_0_clk _01218_ net1071 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[975\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08305__B1 net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09502__C1 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12938_ clknet_leaf_22_clk _00176_ net1163 vssd1 vssd1 vccd1 vccd1 net126 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_34_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10885__S net1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11860__B1 net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13227__CLK clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12869_ clknet_leaf_9_clk _00107_ net1152 vssd1 vssd1 vccd1 vccd1 final_design.data_from_mem\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__11570__A net223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12404__A2 net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06619__B1 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11612__B1 net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07816__C1 _01657_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09281__A1 net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08060_ final_design.cpu.reg_window\[850\] final_design.cpu.reg_window\[882\] net845
+ vssd1 vssd1 vccd1 vccd1 _03011_ sky130_fd_sc_hd__mux2_1
XANTENNA__13377__CLK clknet_leaf_47_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12168__A1 net240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07011_ final_design.cpu.reg_window\[591\] final_design.cpu.reg_window\[623\] net887
+ vssd1 vssd1 vccd1 vccd1 _01962_ sky130_fd_sc_hd__mux2_1
XANTENNA__11915__A1 _06060_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11915__B2 final_design.cpu.reg_window\[411\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1777 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11729__B net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06603__S net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12902__Q net169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08962_ final_design.CPU_instr_adr\[18\] _03793_ final_design.CPU_instr_adr\[19\]
+ vssd1 vssd1 vccd1 vccd1 _03901_ sky130_fd_sc_hd__a21oi_1
X_07913_ net606 _02863_ vssd1 vssd1 vccd1 vccd1 _02864_ sky130_fd_sc_hd__or2_1
X_08893_ _01631_ _01632_ _01662_ _02470_ vssd1 vssd1 vccd1 vccd1 _03839_ sky130_fd_sc_hd__a211o_1
XANTENNA__11143__A2 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout196_A _06016_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07844_ _02791_ _02792_ _02793_ _02794_ net685 net694 vssd1 vssd1 vccd1 vccd1 _02795_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__10351__B1 net1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06839__A _01785_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07434__S net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14002__CLK clknet_leaf_44_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11464__B net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07775_ final_design.cpu.reg_window\[664\] final_design.cpu.reg_window\[696\] net862
+ vssd1 vssd1 vccd1 vccd1 _02726_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06558__B _01507_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_1873 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09514_ _03029_ net445 net442 _03027_ _04432_ vssd1 vssd1 vccd1 vccd1 _04433_ sky130_fd_sc_hd__o221a_1
XFILLER_0_78_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06726_ final_design.cpu.reg_window\[856\] final_design.cpu.reg_window\[888\] net944
+ vssd1 vssd1 vccd1 vccd1 _01677_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_1737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09502__X _04421_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09445_ _04362_ _04363_ vssd1 vssd1 vccd1 vccd1 _04364_ sky130_fd_sc_hd__nor2_1
XANTENNA__10654__B2 net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11851__B1 net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06657_ final_design.cpu.reg_window\[154\] final_design.cpu.reg_window\[186\] net941
+ vssd1 vssd1 vccd1 vccd1 _01608_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12576__A net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout628_A net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout249_X net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14152__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08265__S net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09376_ net492 _04225_ _04294_ vssd1 vssd1 vccd1 vccd1 _04295_ sky130_fd_sc_hd__or3b_1
X_06588_ net742 _01537_ net665 vssd1 vssd1 vccd1 vccd1 _01539_ sky130_fd_sc_hd__a21o_2
X_08327_ final_design.cpu.reg_window\[968\] final_design.cpu.reg_window\[1000\] net816
+ vssd1 vssd1 vccd1 vccd1 _03278_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1060_X net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout416_X net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08258_ final_design.cpu.reg_window\[202\] final_design.cpu.reg_window\[234\] net814
+ vssd1 vssd1 vccd1 vccd1 _03209_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07209_ final_design.cpu.reg_window\[328\] final_design.cpu.reg_window\[360\] net901
+ vssd1 vssd1 vccd1 vccd1 _02160_ sky130_fd_sc_hd__mux2_1
XANTENNA__09024__A1 net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1833 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_18_Left_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08189_ _03136_ _03137_ _03138_ _03139_ net676 net698 vssd1 vssd1 vccd1 vccd1 _03140_
+ sky130_fd_sc_hd__mux4_1
X_10220_ final_design.uart.BAUD_counter\[7\] _05099_ net799 vssd1 vssd1 vccd1 vccd1
+ _05101_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_82_1877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11639__B net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout785_X net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11382__A2 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10151_ _05046_ _05048_ _05049_ vssd1 vssd1 vccd1 vccd1 final_design.vga.h_next_count\[2\]
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_7_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12894__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10082_ final_design.VGA_data_control.v_count\[7\] final_design.VGA_data_control.v_count\[5\]
+ final_design.VGA_data_control.v_count\[6\] vssd1 vssd1 vccd1 vccd1 _04998_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout952_X net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13910_ clknet_leaf_59_clk _01141_ net1126 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[898\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_67_2501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07344__S net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_27_Left_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13841_ clknet_leaf_34_clk _01072_ net1243 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[829\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_1913 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13772_ clknet_leaf_46_clk _01003_ net1214 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[760\]
+ sky130_fd_sc_hd__dfrtp_1
X_10984_ _05694_ _05709_ vssd1 vssd1 vccd1 vccd1 _05711_ sky130_fd_sc_hd__or2_1
XANTENNA__10645__A1 net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11842__A0 net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12723_ final_design.VGA_data_control.v_count\[2\] _06359_ vssd1 vssd1 vccd1 vccd1
+ _06364_ sky130_fd_sc_hd__xor2_2
X_14226__1280 vssd1 vssd1 vccd1 vccd1 _14226__1280/HI net1280 sky130_fd_sc_hd__conb_1
X_12654_ _06314_ net1421 net979 vssd1 vssd1 vccd1 vccd1 _01329_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11605_ net232 net2369 net298 vssd1 vssd1 vccd1 vccd1 _00435_ sky130_fd_sc_hd__mux2_1
X_12585_ net1813 net997 net983 final_design.data_from_mem\[3\] vssd1 vssd1 vccd1 vccd1
+ _01278_ sky130_fd_sc_hd__a22o_1
XFILLER_0_68_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11536_ net803 _02358_ _02095_ vssd1 vssd1 vccd1 vccd1 _06123_ sky130_fd_sc_hd__and3b_4
XANTENNA__08471__C1 _02294_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06771__X _01722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14255_ net1309 vssd1 vssd1 vccd1 vccd1 gpio_out[33] sky130_fd_sc_hd__buf_2
X_11467_ net212 net2435 net306 vssd1 vssd1 vccd1 vccd1 _00351_ sky130_fd_sc_hd__mux2_1
X_13206_ clknet_leaf_60_clk _00437_ net1138 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[194\]
+ sky130_fd_sc_hd__dfrtp_1
X_10418_ net1456 net1027 _05192_ net246 vssd1 vssd1 vccd1 vccd1 _00150_ sky130_fd_sc_hd__a22o_1
XANTENNA__09566__A2 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1917 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14186_ net169 vssd1 vssd1 vccd1 vccd1 net168 sky130_fd_sc_hd__clkbuf_1
X_11398_ net436 net583 _06082_ net317 net1998 vssd1 vssd1 vccd1 vccd1 _00305_ sky130_fd_sc_hd__a32o_1
XANTENNA__07121__S0 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13137_ clknet_leaf_34_clk _00368_ net1242 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[125\]
+ sky130_fd_sc_hd__dfrtp_1
X_10349_ wb_manage.BUSY_O wb_manage.prev_BUSY_O net1023 vssd1 vssd1 vccd1 vccd1 _05170_
+ sky130_fd_sc_hd__and3b_2
XFILLER_0_0_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13068_ clknet_leaf_47_clk _00299_ net1203 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[56\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14025__CLK clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12322__A1 net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12019_ _06221_ net293 net403 net1928 vssd1 vssd1 vccd1 vccd1 _00750_ sky130_fd_sc_hd__a22o_1
XANTENNA__12160__S net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14175__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12086__B1 net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07560_ net741 _01480_ vssd1 vssd1 vccd1 vccd1 _02511_ sky130_fd_sc_hd__nor2_1
XFILLER_0_18_1543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06511_ final_design.data_from_mem\[6\] net1040 net994 net991 vssd1 vssd1 vccd1 vccd1
+ _01462_ sky130_fd_sc_hd__or4_1
XANTENNA__11833__A0 net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_0_clk_X clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1554 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07491_ _02439_ _02440_ _02187_ vssd1 vssd1 vccd1 vccd1 _02442_ sky130_fd_sc_hd__o21a_1
XFILLER_0_76_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12396__A net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11504__S net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09230_ _03423_ _04148_ vssd1 vssd1 vccd1 vccd1 _04149_ sky130_fd_sc_hd__nand2_2
X_06442_ final_design.reqhand.current_client\[1\] net1041 _01395_ vssd1 vssd1 vccd1
+ vccd1 _01396_ sky130_fd_sc_hd__o21ai_2
XTAP_TAPCELL_ROW_17_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12776__7_A clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1107 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12389__A1 net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09161_ _04078_ _04079_ vssd1 vssd1 vccd1 vccd1 _04080_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_20_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08112_ _03059_ _03060_ _03061_ _03062_ net675 net691 vssd1 vssd1 vccd1 vccd1 _03063_
+ sky130_fd_sc_hd__mux4_1
X_09092_ _03784_ _04015_ vssd1 vssd1 vccd1 vccd1 _04016_ sky130_fd_sc_hd__or2_1
XANTENNA__11299__X _05996_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08043_ net602 _02991_ _02966_ _01850_ vssd1 vssd1 vccd1 vccd1 _02994_ sky130_fd_sc_hd__o211a_1
Xhold900 final_design.cpu.reg_window\[272\] vssd1 vssd1 vccd1 vccd1 net2242 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold911 final_design.cpu.reg_window\[394\] vssd1 vssd1 vccd1 vccd1 net2253 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout209_A net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold922 final_design.cpu.reg_window\[941\] vssd1 vssd1 vccd1 vccd1 net2264 sky130_fd_sc_hd__dlygate4sd3_1
Xhold933 final_design.cpu.reg_window\[356\] vssd1 vssd1 vccd1 vccd1 net2275 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12010__B1 net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold944 final_design.cpu.reg_window\[151\] vssd1 vssd1 vccd1 vccd1 net2286 sky130_fd_sc_hd__dlygate4sd3_1
Xhold955 final_design.cpu.reg_window\[1011\] vssd1 vssd1 vccd1 vccd1 net2297 sky130_fd_sc_hd__dlygate4sd3_1
Xhold966 final_design.cpu.reg_window\[957\] vssd1 vssd1 vccd1 vccd1 net2308 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold977 final_design.cpu.reg_window\[121\] vssd1 vssd1 vccd1 vccd1 net2319 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10021__C1 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1020_A _06298_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold988 final_design.cpu.reg_window\[449\] vssd1 vssd1 vccd1 vccd1 net2330 sky130_fd_sc_hd__dlygate4sd3_1
X_09994_ net477 _04411_ _04912_ net319 vssd1 vssd1 vccd1 vccd1 _04913_ sky130_fd_sc_hd__o211a_1
Xhold999 final_design.cpu.reg_window\[611\] vssd1 vssd1 vccd1 vccd1 net2341 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1118_A net100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1861 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08945_ final_design.CPU_instr_adr\[21\] _03795_ vssd1 vssd1 vccd1 vccd1 _03886_
+ sky130_fd_sc_hd__xnor2_1
XANTENNA__08401__X _03352_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout480_A _03484_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout578_A net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13961__RESET_B net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08876_ _03823_ _02474_ vssd1 vssd1 vccd1 vccd1 _03824_ sky130_fd_sc_hd__and2b_1
XANTENNA__07164__S net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07827_ _02774_ _02775_ _02776_ _02777_ net685 net693 vssd1 vssd1 vccd1 vccd1 _02778_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__11194__B _05900_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout366_X net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout745_A net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12077__B1 net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07758_ final_design.cpu.reg_window\[280\] final_design.cpu.reg_window\[312\] net864
+ vssd1 vssd1 vccd1 vccd1 _02709_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11824__A0 net209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13542__CLK clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06709_ net743 _01659_ net665 vssd1 vssd1 vccd1 vccd1 _01660_ sky130_fd_sc_hd__a21o_2
XANTENNA_fanout912_A net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07689_ _02637_ _02639_ vssd1 vssd1 vccd1 vccd1 _02640_ sky130_fd_sc_hd__nor2_1
XFILLER_0_71_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12092__A3 net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11414__S net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09428_ _04334_ _04335_ _04346_ net262 vssd1 vssd1 vccd1 vccd1 _04347_ sky130_fd_sc_hd__o211a_1
XFILLER_0_63_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout700_X net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09359_ net489 _04277_ _04276_ vssd1 vssd1 vccd1 vccd1 _04278_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_10_1827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13692__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12370_ net1819 net238 net269 vssd1 vssd1 vccd1 vccd1 _01081_ sky130_fd_sc_hd__mux2_1
XANTENNA__09796__A2 net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_976 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11321_ _01788_ net642 _06014_ net643 _06013_ vssd1 vssd1 vccd1 vccd1 _06015_ sky130_fd_sc_hd__a221o_1
X_14040_ clknet_leaf_15_clk _00032_ net1095 vssd1 vssd1 vccd1 vccd1 final_design.uart.BAUD_counter\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_11252_ net660 _03944_ net732 vssd1 vssd1 vccd1 vccd1 _05954_ sky130_fd_sc_hd__o21ai_1
XANTENNA__12001__B1 net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09548__A2 _04373_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14048__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10203_ final_design.uart.BAUD_counter\[0\] net798 vssd1 vssd1 vccd1 vccd1 _00006_
+ sky130_fd_sc_hd__and2b_1
X_11183_ net735 _04009_ _05892_ vssd1 vssd1 vccd1 vccd1 _05893_ sky130_fd_sc_hd__a21o_1
XFILLER_0_63_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input41_A mem_adr_start[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10134_ final_design.VGA_data_control.h_count\[0\] _05037_ vssd1 vssd1 vccd1 vccd1
+ _05038_ sky130_fd_sc_hd__or2_1
XANTENNA__12304__A1 net244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13072__CLK clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08678__B net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10065_ _04510_ _04511_ _04550_ _04551_ vssd1 vssd1 vccd1 vccd1 _04984_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__09126__Y _04045_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07074__S net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10866__B2 net1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12068__B1 net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13824_ clknet_leaf_10_clk _01055_ net1098 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[812\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12607__A2 net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08694__A _02772_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07802__S net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10967_ _05673_ _05692_ net1003 vssd1 vssd1 vccd1 vccd1 _05695_ sky130_fd_sc_hd__o21a_1
XFILLER_0_70_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13755_ clknet_leaf_65_clk _00986_ net1070 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[743\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10288__X final_design.cpu.Error vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12083__A3 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12706_ _06340_ _06346_ _06345_ net1051 vssd1 vssd1 vccd1 vccd1 _06347_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_35_1186 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09302__B net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10898_ _05590_ _05612_ _05611_ vssd1 vssd1 vccd1 vccd1 _05628_ sky130_fd_sc_hd__a21bo_1
X_13686_ clknet_leaf_61_clk _00917_ net1137 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[674\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_31_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10448__B net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12637_ final_design.VGA_data_control.ready_data\[6\] net1021 net976 final_design.data_from_mem\[6\]
+ vssd1 vssd1 vccd1 vccd1 _06306_ sky130_fd_sc_hd__a22o_1
XFILLER_0_25_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12240__B1 net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12568_ final_design.uart.receiving final_design.uart.working_data\[4\] vssd1 vssd1
+ vccd1 vccd1 _06289_ sky130_fd_sc_hd__and2_1
XFILLER_0_14_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11519_ net2206 _06120_ _06121_ net433 vssd1 vssd1 vccd1 vccd1 _00387_ sky130_fd_sc_hd__a22o_1
XANTENNA__12155__S net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10464__A _04940_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12499_ _06160_ net349 net327 net1810 vssd1 vssd1 vccd1 vccd1 _01204_ sky130_fd_sc_hd__a22o_1
XANTENNA__07893__S1 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold207 final_design.cpu.reg_window\[732\] vssd1 vssd1 vccd1 vccd1 net1549 sky130_fd_sc_hd__dlygate4sd3_1
Xhold218 final_design.cpu.reg_window\[646\] vssd1 vssd1 vccd1 vccd1 net1560 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_65_1861 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold229 final_design.cpu.reg_window\[518\] vssd1 vssd1 vccd1 vccd1 net1571 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09539__A2 net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14238_ net1292 vssd1 vssd1 vccd1 vccd1 gpio_out[16] sky130_fd_sc_hd__buf_2
X_14169_ clknet_leaf_20_clk _01343_ net1158 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.data_to_VGA\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13415__CLK clknet_leaf_63_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08211__A2 _03160_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1889 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout709 net710 vssd1 vssd1 vccd1 vccd1 net709 sky130_fd_sc_hd__buf_4
XFILLER_0_0_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06991_ _01940_ _01941_ vssd1 vssd1 vccd1 vccd1 _01942_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_77_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_33_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11295__A net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08730_ final_design.CPU_instr_adr\[14\] _02000_ vssd1 vssd1 vccd1 vccd1 _03681_
+ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_33_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13565__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08661_ _02545_ _03610_ _02542_ vssd1 vssd1 vccd1 vccd1 _03612_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_56_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07612_ _02559_ _02560_ _02561_ _02562_ net688 net705 vssd1 vssd1 vccd1 vccd1 _02563_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_72_1821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08592_ final_design.cpu.reg_window\[704\] final_design.cpu.reg_window\[736\] net826
+ vssd1 vssd1 vccd1 vccd1 _03543_ sky130_fd_sc_hd__mux2_1
XANTENNA__06676__X _01627_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06930__C1 _01821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07543_ _02490_ _02491_ _02492_ _02493_ net774 net792 vssd1 vssd1 vccd1 vccd1 _02494_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__11806__B1 net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12074__A3 net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07474_ net741 _01497_ _02420_ _02421_ vssd1 vssd1 vccd1 vccd1 _02425_ sky130_fd_sc_hd__a211o_2
XFILLER_0_14_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07581__S0 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09213_ _02866_ _04129_ _04130_ _04128_ vssd1 vssd1 vccd1 vccd1 _04132_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_57_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06425_ final_design.reqhand.instruction\[20\] vssd1 vssd1 vccd1 vccd1 _01380_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout326_A net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1068_A net1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09144_ net595 net525 _02325_ _02422_ vssd1 vssd1 vccd1 vccd1 _04063_ sky130_fd_sc_hd__o211a_1
XANTENNA__12231__B1 net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08543__S net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11585__A2 net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09075_ _03723_ _04000_ vssd1 vssd1 vccd1 vccd1 _04001_ sky130_fd_sc_hd__and2_1
XFILLER_0_31_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1235_A net1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1901 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08026_ _02973_ _02974_ _02975_ _02976_ net679 net699 vssd1 vssd1 vccd1 vccd1 _02977_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_60_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_9_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold730 final_design.cpu.reg_window\[615\] vssd1 vssd1 vccd1 vccd1 net2072 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold741 final_design.cpu.reg_window\[427\] vssd1 vssd1 vccd1 vccd1 net2083 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13095__CLK clknet_leaf_62_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold752 final_design.cpu.reg_window\[762\] vssd1 vssd1 vccd1 vccd1 net2094 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09935__C1 _04341_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold763 final_design.cpu.reg_window\[277\] vssd1 vssd1 vccd1 vccd1 net2105 sky130_fd_sc_hd__dlygate4sd3_1
Xhold774 final_design.cpu.reg_window\[439\] vssd1 vssd1 vccd1 vccd1 net2116 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1023_X net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold785 final_design.cpu.reg_window\[538\] vssd1 vssd1 vccd1 vccd1 net2127 sky130_fd_sc_hd__dlygate4sd3_1
Xhold796 final_design.cpu.reg_window\[385\] vssd1 vssd1 vccd1 vccd1 net2138 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07410__B1 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout862_A net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09977_ _03327_ _04895_ vssd1 vssd1 vccd1 vccd1 _04896_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout483_X net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13908__CLK clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08928_ net257 _03869_ net1014 vssd1 vssd1 vccd1 vccd1 _03871_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10841__A1_N net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout650_X net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08859_ net624 _03806_ _03808_ net256 vssd1 vssd1 vccd1 vccd1 _03809_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout748_X net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11870_ _06017_ net640 net288 net519 net2135 vssd1 vssd1 vccd1 vccd1 _00616_ sky130_fd_sc_hd__a32o_1
XANTENNA__06586__X _01537_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10821_ net960 _05553_ _05554_ _04042_ vssd1 vssd1 vccd1 vccd1 _05555_ sky130_fd_sc_hd__a22o_1
XFILLER_0_51_1905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout915_X net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11144__S net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1861 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10752_ _05467_ _05470_ _05488_ vssd1 vssd1 vccd1 vccd1 _05489_ sky130_fd_sc_hd__o21ba_1
X_13540_ clknet_leaf_54_clk _00771_ net1177 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[528\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12470__B1 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13471_ clknet_leaf_7_clk _00702_ net1134 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[459\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07883__A_N net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10683_ net1411 net1031 net1003 _05423_ vssd1 vssd1 vccd1 vccd1 _00184_ sky130_fd_sc_hd__a22o_1
XFILLER_0_82_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12422_ _06110_ net356 net341 net2107 vssd1 vssd1 vccd1 vccd1 _01131_ sky130_fd_sc_hd__a22o_1
XFILLER_0_30_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12222__B1 net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09313__S1 net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09769__A2 net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input89_A memory_size[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08306__X _03257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07324__S0 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12353_ _06236_ net500 net361 net2201 vssd1 vssd1 vccd1 vccd1 _01065_ sky130_fd_sc_hd__a22o_1
XFILLER_0_23_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13438__CLK clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06988__C1 _01821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11304_ net738 _03902_ vssd1 vssd1 vccd1 vccd1 _06000_ sky130_fd_sc_hd__nand2_1
XANTENNA__07069__S net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12284_ net585 _06214_ net512 net370 net1703 vssd1 vssd1 vccd1 vccd1 _00999_ sky130_fd_sc_hd__a32o_1
XANTENNA__11328__A2 net235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14023_ clknet_leaf_63_clk _01254_ net1123 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[1011\]
+ sky130_fd_sc_hd__dfrtp_1
X_11235_ net644 _05936_ _05937_ _05938_ net655 vssd1 vssd1 vccd1 vccd1 _05939_ sky130_fd_sc_hd__a221o_1
XANTENNA__13812__RESET_B net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13588__CLK clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11166_ net662 _04020_ net734 vssd1 vssd1 vccd1 vccd1 _05878_ sky130_fd_sc_hd__a21o_1
X_10117_ net1051 _05023_ final_design.VGA_data_control.v_count\[5\] vssd1 vssd1 vccd1
+ vccd1 _05028_ sky130_fd_sc_hd__a21o_1
XANTENNA__12289__B1 net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11097_ _05798_ _05815_ _05814_ vssd1 vssd1 vccd1 vccd1 _05818_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11546__C net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10048_ _04529_ _04530_ _04616_ vssd1 vssd1 vccd1 vccd1 _04967_ sky130_fd_sc_hd__o21ba_1
XANTENNA__08052__S1 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold90 final_design.VGA_data_control.data_to_VGA\[29\] vssd1 vssd1 vccd1 vccd1 net1432
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11843__A net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07532__S net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13807_ clknet_leaf_42_clk _01038_ net1223 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[795\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11562__B net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11999_ _06201_ net276 net400 net1883 vssd1 vssd1 vccd1 vccd1 _00730_ sky130_fd_sc_hd__a22o_1
XFILLER_0_50_1415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11264__A1 _04613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13738_ clknet_leaf_50_clk _00969_ net1168 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[726\]
+ sky130_fd_sc_hd__dfrtp_1
X_14249__1303 vssd1 vssd1 vccd1 vccd1 _14249__1303/HI net1303 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_41_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13669_ clknet_leaf_49_clk _00900_ net1181 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[657\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_41_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07190_ net757 _02140_ vssd1 vssd1 vccd1 vccd1 _02141_ sky130_fd_sc_hd__or2_1
XANTENNA__12213__B1 net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11567__A2 net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_1219 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09900_ _03638_ _04087_ net440 _03637_ _04811_ vssd1 vssd1 vccd1 vccd1 _04819_ sky130_fd_sc_hd__a221o_1
XFILLER_0_50_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_1555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout506 net507 vssd1 vssd1 vccd1 vccd1 net506 sky130_fd_sc_hd__buf_4
XFILLER_0_6_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09831_ _04745_ _04747_ vssd1 vssd1 vccd1 vccd1 _04750_ sky130_fd_sc_hd__xnor2_1
Xfanout517 net518 vssd1 vssd1 vccd1 vccd1 net517 sky130_fd_sc_hd__buf_4
XFILLER_0_22_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout528 _02356_ vssd1 vssd1 vccd1 vccd1 net528 sky130_fd_sc_hd__buf_2
Xfanout539 _02058_ vssd1 vssd1 vccd1 vccd1 net539 sky130_fd_sc_hd__buf_2
XANTENNA__07943__A1 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12955__CLK clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06974_ final_design.cpu.reg_window\[848\] final_design.cpu.reg_window\[880\] net923
+ vssd1 vssd1 vccd1 vccd1 _01925_ sky130_fd_sc_hd__mux2_1
X_09762_ _04426_ _04680_ net448 vssd1 vssd1 vccd1 vccd1 _04681_ sky130_fd_sc_hd__a21o_1
XFILLER_0_20_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08713_ _03662_ _03663_ vssd1 vssd1 vccd1 vccd1 _03664_ sky130_fd_sc_hd__and2_1
X_09693_ _03164_ _04498_ _04611_ _03649_ _04045_ vssd1 vssd1 vccd1 vccd1 _04612_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_20_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12295__A3 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout276_A net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08644_ _03040_ _02772_ vssd1 vssd1 vccd1 vccd1 _03595_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_1_246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09791__S1 net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08575_ final_design.cpu.reg_window\[256\] final_design.cpu.reg_window\[288\] net827
+ vssd1 vssd1 vccd1 vccd1 _03526_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout443_A net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10058__A2 _04530_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07526_ _01509_ _02476_ _01508_ vssd1 vssd1 vccd1 vccd1 _02477_ sky130_fd_sc_hd__a21o_1
XANTENNA__11255__A1 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11899__S net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07457_ final_design.cpu.reg_window\[832\] final_design.cpu.reg_window\[864\] net915
+ vssd1 vssd1 vccd1 vccd1 _02408_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout231_X net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout610_A net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout329_X net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout708_A net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06408_ final_design.CPU_instr_adr\[15\] vssd1 vssd1 vccd1 vccd1 _01363_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12204__B1 net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07388_ final_design.cpu.reg_window\[2\] final_design.cpu.reg_window\[34\] net918
+ vssd1 vssd1 vccd1 vccd1 _02339_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09127_ net659 _04045_ vssd1 vssd1 vccd1 vccd1 _04046_ sky130_fd_sc_hd__and2_4
XFILLER_0_60_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09058_ final_design.CPU_instr_adr\[8\] _03786_ vssd1 vssd1 vccd1 vccd1 _03986_ sky130_fd_sc_hd__nor2_1
XFILLER_0_66_1499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13730__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08009_ _02954_ _02959_ net714 vssd1 vssd1 vccd1 vccd1 _02960_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout698_X net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07684__Y _02635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold560 final_design.cpu.reg_window\[689\] vssd1 vssd1 vccd1 vccd1 net1902 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10518__B1 net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold571 final_design.cpu.reg_window\[208\] vssd1 vssd1 vccd1 vccd1 net1913 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09384__A0 net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11020_ _04040_ _05742_ _05744_ _04042_ net963 vssd1 vssd1 vccd1 vccd1 _05745_ sky130_fd_sc_hd__a221o_1
Xhold582 final_design.cpu.reg_window\[880\] vssd1 vssd1 vccd1 vccd1 net1924 sky130_fd_sc_hd__dlygate4sd3_1
Xhold593 final_design.cpu.reg_window\[874\] vssd1 vssd1 vccd1 vccd1 net1935 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_1805 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11647__B net196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout865_X net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_2585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_1849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_2596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13880__CLK clknet_leaf_63_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07563__D net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10978__S net1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12971_ clknet_leaf_19_clk net1343 net1156 vssd1 vssd1 vccd1 vccd1 wb_manage.prev_BUSY_O
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09687__A1 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12286__A3 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11922_ net230 net2494 net408 vssd1 vssd1 vccd1 vccd1 _00659_ sky130_fd_sc_hd__mux2_1
XANTENNA__12691__B1 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08448__S net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13110__CLK clknet_leaf_61_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07793__S0 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07205__X _02156_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11853_ _06103_ net279 net517 net1894 vssd1 vssd1 vccd1 vccd1 _00603_ sky130_fd_sc_hd__a22o_1
XFILLER_0_55_1882 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_2378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10804_ net669 _05527_ _05538_ vssd1 vssd1 vccd1 vccd1 _05539_ sky130_fd_sc_hd__o21ai_1
XANTENNA__11246__A1 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11784_ net648 net555 net215 vssd1 vssd1 vccd1 vccd1 _06232_ sky130_fd_sc_hd__and3_1
XFILLER_0_51_1746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_2389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14082__RESET_B net1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11797__A2 net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13523_ clknet_leaf_39_clk _00754_ net1210 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[511\]
+ sky130_fd_sc_hd__dfrtp_1
X_10735_ net960 _05471_ _05472_ _04042_ vssd1 vssd1 vccd1 vccd1 _05473_ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_40_clk_X clknet_leaf_40_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13260__CLK clknet_leaf_46_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10666_ net70 final_design.VGA_adr\[9\] vssd1 vssd1 vccd1 vccd1 _05407_ sky130_fd_sc_hd__xnor2_1
X_13454_ clknet_leaf_43_clk _00685_ net1222 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[442\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11549__A2 net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12405_ _06103_ net343 net338 net2478 vssd1 vssd1 vccd1 vccd1 _01115_ sky130_fd_sc_hd__a22o_1
X_13385_ clknet_leaf_36_clk _00616_ net1236 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[373\]
+ sky130_fd_sc_hd__dfrtp_1
X_10597_ _05340_ _05341_ net961 vssd1 vssd1 vccd1 vccd1 _05342_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_11_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12210__A3 net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput109 net109 vssd1 vssd1 vccd1 vccd1 ADR_O[17] sky130_fd_sc_hd__clkbuf_4
X_12336_ net2270 net361 net348 _05898_ vssd1 vssd1 vccd1 vccd1 _01048_ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_55_clk_X clknet_leaf_55_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12433__S net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12267_ net565 _06197_ net505 net369 net1985 vssd1 vssd1 vccd1 vccd1 _00982_ sky130_fd_sc_hd__a32o_1
XANTENNA__12978__CLK clknet_leaf_19_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08178__B2 net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14006_ clknet_leaf_59_clk _01237_ net1138 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[994\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11218_ net731 _03981_ _05923_ vssd1 vssd1 vccd1 vccd1 _05924_ sky130_fd_sc_hd__o21a_1
XANTENNA__09308__A net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09914__A2 net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12198_ net566 _06126_ net506 net377 net2358 vssd1 vssd1 vccd1 vccd1 _00916_ sky130_fd_sc_hd__a32o_1
XANTENNA__11182__B1 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11149_ net651 _05860_ _05862_ vssd1 vssd1 vccd1 vccd1 _05863_ sky130_fd_sc_hd__and3_1
XFILLER_0_37_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12277__A3 net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06690_ final_design.cpu.reg_window\[153\] final_design.cpu.reg_window\[185\] net935
+ vssd1 vssd1 vccd1 vccd1 _01641_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06900__A2 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13603__CLK clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08360_ final_design.cpu.reg_window\[775\] final_design.cpu.reg_window\[807\] net811
+ vssd1 vssd1 vccd1 vccd1 _03311_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07311_ final_design.cpu.reg_window\[709\] final_design.cpu.reg_window\[741\] net921
+ vssd1 vssd1 vccd1 vccd1 _02262_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07536__S0 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09697__B _04613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08291_ final_design.cpu.reg_window\[137\] final_design.cpu.reg_window\[169\] net807
+ vssd1 vssd1 vccd1 vccd1 _03242_ sky130_fd_sc_hd__mux2_1
XANTENNA__11512__S net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07242_ net757 _02192_ vssd1 vssd1 vccd1 vccd1 _02193_ sky130_fd_sc_hd__or2_1
XFILLER_0_27_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08093__S net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12737__A1 _05058_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13753__CLK clknet_leaf_56_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07173_ _02120_ _02121_ _02122_ _02123_ net765 net780 vssd1 vssd1 vccd1 vccd1 _02124_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__09984__Y _04903_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09602__B2 net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07839__S1 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11960__A2 net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14109__CLK clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_1472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout303 _06125_ vssd1 vssd1 vccd1 vccd1 net303 sky130_fd_sc_hd__buf_4
Xfanout314 net315 vssd1 vssd1 vccd1 vccd1 net314 sky130_fd_sc_hd__buf_4
Xfanout325 _06285_ vssd1 vssd1 vccd1 vccd1 net325 sky130_fd_sc_hd__buf_4
XANTENNA__11173__B1 net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout393_A _06263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout336 net337 vssd1 vssd1 vccd1 vccd1 net336 sky130_fd_sc_hd__buf_6
XANTENNA__11712__A2 net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09814_ _04618_ _04732_ net470 vssd1 vssd1 vccd1 vccd1 _04733_ sky130_fd_sc_hd__mux2_1
Xfanout347 net350 vssd1 vssd1 vccd1 vccd1 net347 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09381__A3 net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout358 net359 vssd1 vssd1 vccd1 vccd1 net358 sky130_fd_sc_hd__buf_2
XANTENNA__11186__C _05895_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout369 _06274_ vssd1 vssd1 vccd1 vccd1 net369 sky130_fd_sc_hd__buf_4
XANTENNA_fanout1100_A net1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10920__B1 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13133__CLK clknet_leaf_45_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09745_ _04485_ _04663_ net471 vssd1 vssd1 vccd1 vccd1 _04664_ sky130_fd_sc_hd__mux2_1
X_06957_ net886 _01907_ _01896_ _01895_ vssd1 vssd1 vccd1 vccd1 _01908_ sky130_fd_sc_hd__o2bb2a_2
XANTENNA_fanout560_A net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12268__A3 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout279_X net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout658_A _05142_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06888_ final_design.cpu.reg_window\[787\] final_design.cpu.reg_window\[819\] net913
+ vssd1 vssd1 vccd1 vccd1 _01839_ sky130_fd_sc_hd__mux2_1
X_09676_ _02834_ _04330_ _02803_ vssd1 vssd1 vccd1 vccd1 _04595_ sky130_fd_sc_hd__a21oi_2
XANTENNA__06577__A net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08627_ _03572_ _03577_ _03167_ vssd1 vssd1 vccd1 vccd1 _03578_ sky130_fd_sc_hd__a21oi_1
XANTENNA__13283__CLK clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout446_X net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout825_A net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1090_X net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11228__A1 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12425__B1 net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08558_ final_design.cpu.reg_window\[577\] final_design.cpu.reg_window\[609\] net831
+ vssd1 vssd1 vccd1 vccd1 _03509_ sky130_fd_sc_hd__mux2_1
XANTENNA__06864__X _01815_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08629__C1 _02059_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_2990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11779__A2 net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11930__B net244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07509_ _01855_ _02459_ _01856_ vssd1 vssd1 vccd1 vccd1 _02460_ sky130_fd_sc_hd__o21a_1
XANTENNA__10386__X _05174_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08489_ final_design.cpu.reg_window\[771\] final_design.cpu.reg_window\[803\] net831
+ vssd1 vssd1 vccd1 vccd1 _03440_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout613_X net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10987__B1 net1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11422__S net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10520_ _05249_ _05264_ _05263_ vssd1 vssd1 vccd1 vccd1 _05268_ sky130_fd_sc_hd__a21o_1
XFILLER_0_11_1752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10451_ net253 _05209_ net1035 net1396 vssd1 vssd1 vccd1 vccd1 _00166_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_81_1717 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13170_ clknet_leaf_39_clk _00401_ net1210 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[158\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11400__A1 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10382_ net26 net1023 net1007 final_design.data_from_mem\[31\] vssd1 vssd1 vccd1
+ vccd1 _00135_ sky130_fd_sc_hd__o22a_1
XFILLER_0_62_1116 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_2160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_2794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12121_ net1850 net187 net390 vssd1 vssd1 vccd1 vccd1 _00845_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_53_2002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_2171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06958__A2 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11951__A2 net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_2013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_2024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_2035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12052_ net1992 net188 net398 vssd1 vssd1 vccd1 vccd1 _00780_ sky130_fd_sc_hd__mux2_1
XANTENNA__09128__A net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold390 final_design.cpu.reg_window\[246\] vssd1 vssd1 vccd1 vccd1 net1732 sky130_fd_sc_hd__dlygate4sd3_1
X_11003_ net54 _05728_ vssd1 vssd1 vccd1 vccd1 _05729_ sky130_fd_sc_hd__and2_1
X_14248__1302 vssd1 vssd1 vccd1 vccd1 _14248__1302/HI net1302 sky130_fd_sc_hd__conb_1
XANTENNA__10911__B1 net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout870 net871 vssd1 vssd1 vccd1 vccd1 net870 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_79_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout881 net882 vssd1 vssd1 vccd1 vccd1 net881 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_5_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout892 net899 vssd1 vssd1 vccd1 vccd1 net892 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_5_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12259__A3 net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08686__B net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09134__Y _04053_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12954_ clknet_leaf_29_clk _00192_ net1195 vssd1 vssd1 vccd1 vccd1 net111 sky130_fd_sc_hd__dfrtp_1
XANTENNA__06487__A net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1090 final_design.cpu.reg_window\[652\] vssd1 vssd1 vccd1 vccd1 net2432 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_73_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07766__S0 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06569__S1 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11905_ net197 net2310 net274 vssd1 vssd1 vccd1 vccd1 _00647_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12885_ clknet_leaf_19_clk _00123_ net1157 vssd1 vssd1 vccd1 vccd1 final_design.data_from_mem\[19\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_34_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11219__A1 final_design.data_from_mem\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09798__A _04072_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12416__B1 net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11836_ net189 net2043 net267 vssd1 vssd1 vccd1 vccd1 _00588_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13776__CLK clknet_leaf_34_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11767_ net177 net2312 net418 vssd1 vssd1 vccd1 vccd1 _00530_ sky130_fd_sc_hd__mux2_1
XANTENNA__08635__A2 _02961_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06646__A1 net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13506_ clknet_leaf_4_clk _00737_ net1079 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[494\]
+ sky130_fd_sc_hd__dfrtp_1
X_10718_ net40 _05456_ vssd1 vssd1 vccd1 vccd1 _05457_ sky130_fd_sc_hd__xor2_1
X_11698_ net434 net578 _06207_ net296 net1856 vssd1 vssd1 vccd1 vccd1 _00480_ sky130_fd_sc_hd__a32o_1
XANTENNA__10456__B net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_20_clk_A clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13437_ clknet_leaf_2_clk _00668_ net1077 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[425\]
+ sky130_fd_sc_hd__dfrtp_1
X_10649_ _05368_ _05390_ vssd1 vssd1 vccd1 vccd1 _05391_ sky130_fd_sc_hd__nand2_1
X_13368_ clknet_leaf_64_clk _00599_ net1121 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[356\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11942__A2 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12319_ net2174 net195 net365 vssd1 vssd1 vccd1 vccd1 _01033_ sky130_fd_sc_hd__mux2_1
X_13299_ clknet_leaf_40_clk _00530_ net1219 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[287\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09348__B1 net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13156__CLK clknet_leaf_55_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_35_clk_A clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_1694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07860_ net712 _02810_ vssd1 vssd1 vccd1 vccd1 _02811_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_3_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07781__A _01690_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06811_ final_design.cpu.reg_window\[85\] final_design.cpu.reg_window\[117\] net947
+ vssd1 vssd1 vccd1 vccd1 _01762_ sky130_fd_sc_hd__mux2_1
X_07791_ final_design.cpu.reg_window\[473\] final_design.cpu.reg_window\[505\] net853
+ vssd1 vssd1 vccd1 vccd1 _02742_ sky130_fd_sc_hd__mux2_1
XANTENNA__11507__S net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06742_ final_design.cpu.reg_window\[343\] final_design.cpu.reg_window\[375\] net931
+ vssd1 vssd1 vccd1 vccd1 _01693_ sky130_fd_sc_hd__mux2_1
X_09530_ net261 _04433_ _04445_ _04448_ vssd1 vssd1 vccd1 vccd1 _04449_ sky130_fd_sc_hd__and4_1
XFILLER_0_17_1416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09461_ _04231_ _04367_ _04372_ _04379_ net261 vssd1 vssd1 vccd1 vccd1 _04380_ sky130_fd_sc_hd__o2111ai_2
X_06673_ _01620_ _01621_ _01622_ _01623_ net775 net793 vssd1 vssd1 vccd1 vccd1 _01624_
+ sky130_fd_sc_hd__mux4_1
X_08412_ final_design.cpu.reg_window\[453\] final_design.cpu.reg_window\[485\] net838
+ vssd1 vssd1 vccd1 vccd1 _03363_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09392_ _04056_ _04310_ vssd1 vssd1 vccd1 vccd1 _04311_ sky130_fd_sc_hd__nand2b_1
XANTENNA__12407__B1 net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08343_ _03293_ vssd1 vssd1 vccd1 vccd1 _03294_ sky130_fd_sc_hd__inv_2
XANTENNA__09284__C1 _02422_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10969__B1 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout239_A net240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09995__X _04914_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07834__B1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11630__A1 net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08274_ _02128_ net611 vssd1 vssd1 vccd1 vccd1 _03225_ sky130_fd_sc_hd__nor2_1
XFILLER_0_7_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07225_ _02172_ _02173_ _02174_ _02175_ net764 net780 vssd1 vssd1 vccd1 vccd1 _02176_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_61_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout406_A _06255_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1148_A net1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07156_ net750 _02106_ vssd1 vssd1 vccd1 vccd1 _02107_ sky130_fd_sc_hd__or2_1
XFILLER_0_15_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12581__B net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08485__S1 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11394__B1 _06078_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11933__A2 net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11478__A net197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11277__A2_N _05947_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07087_ _02034_ _02035_ _02036_ _02037_ net765 net785 vssd1 vssd1 vccd1 vccd1 _02038_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__14081__CLK clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1109 net1116 vssd1 vssd1 vccd1 vccd1 net1109 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout775_A net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout396_X net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13649__CLK clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08562__A1 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07996__S0 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout177 _06089_ vssd1 vssd1 vccd1 vccd1 net177 sky130_fd_sc_hd__buf_2
XFILLER_0_76_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout188 _06045_ vssd1 vssd1 vccd1 vccd1 net188 sky130_fd_sc_hd__buf_2
Xfanout199 net200 vssd1 vssd1 vccd1 vccd1 net199 sky130_fd_sc_hd__buf_2
XANTENNA_fanout942_A net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07989_ final_design.cpu.reg_window\[464\] final_design.cpu.reg_window\[496\] net846
+ vssd1 vssd1 vccd1 vccd1 _02940_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout563_X net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_29_Right_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11417__S net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09728_ _04643_ _04646_ net491 vssd1 vssd1 vccd1 vccd1 _04647_ sky130_fd_sc_hd__mux2_1
XANTENNA__13799__CLK clknet_leaf_61_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_65_2440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09659_ net480 _04458_ vssd1 vssd1 vccd1 vccd1 _04578_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout730_X net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout828_X net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_2927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_2304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12670_ _06322_ net1445 net978 vssd1 vssd1 vccd1 vccd1 _01337_ sky130_fd_sc_hd__mux2_1
XANTENNA__10672__A2 net1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_2949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11621_ net220 net630 vssd1 vssd1 vccd1 vccd1 _06168_ sky130_fd_sc_hd__and2_1
XANTENNA__06971__S1 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13029__CLK clknet_leaf_49_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11552_ net558 net243 net634 vssd1 vssd1 vccd1 vccd1 _06132_ sky130_fd_sc_hd__and3_1
XANTENNA__08027__A net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_38_Right_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09290__A2 net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_2211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10503_ net93 final_design.VGA_adr\[1\] vssd1 vssd1 vccd1 vccd1 _05252_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_59_2222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_2856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11483_ net191 net640 vssd1 vssd1 vccd1 vccd1 _06110_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_59_2233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_2867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_2878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input71_A memory_size[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10434_ _02929_ net592 vssd1 vssd1 vccd1 vccd1 _05201_ sky130_fd_sc_hd__nor2_2
X_13222_ clknet_leaf_50_clk _00453_ net1169 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[210\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07866__A net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11924__A2 net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10365_ net7 net1025 net1008 final_design.data_from_mem\[14\] vssd1 vssd1 vccd1 vccd1
+ _00118_ sky130_fd_sc_hd__a22o_1
X_13153_ clknet_leaf_49_clk _00384_ net1184 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[141\]
+ sky130_fd_sc_hd__dfrtp_1
X_12104_ net1907 net218 net388 vssd1 vssd1 vccd1 vccd1 _00828_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13084_ clknet_leaf_3_clk _00315_ net1068 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[72\]
+ sky130_fd_sc_hd__dfrtp_1
X_10296_ final_design.VGA_data_control.h_count\[1\] net1049 final_design.VGA_data_control.data_to_VGA\[5\]
+ vssd1 vssd1 vccd1 vccd1 _05150_ sky130_fd_sc_hd__and3b_1
XANTENNA__11137__B1 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12035_ net1925 net220 net396 vssd1 vssd1 vccd1 vccd1 _00763_ sky130_fd_sc_hd__mux2_1
XANTENNA__11688__A1 net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06769__X _01720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_47_Right_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09750__B1 _04222_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10360__B2 final_design.data_from_mem\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09305__B net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13986_ clknet_leaf_4_clk _01217_ net1080 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[974\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08305__A1 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07106__A net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12937_ clknet_leaf_22_clk _00175_ net1163 vssd1 vssd1 vccd1 vccd1 net123 sky130_fd_sc_hd__dfrtp_2
XFILLER_0_76_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_1594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12868_ clknet_leaf_25_clk _00106_ net1151 vssd1 vssd1 vccd1 vccd1 final_design.data_from_mem\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_31_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11570__B net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11819_ net221 net1967 net264 vssd1 vssd1 vccd1 vccd1 _00571_ sky130_fd_sc_hd__mux2_1
XANTENNA__12158__S net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_56_Right_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08164__S0 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13397__RESET_B net1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11612__A1 net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09281__A2 net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07010_ final_design.cpu.reg_window\[655\] final_design.cpu.reg_window\[687\] net887
+ vssd1 vssd1 vccd1 vccd1 _01961_ sky130_fd_sc_hd__mux2_1
XANTENNA__06680__A _01627_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11915__A2 _06248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07044__A1 net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1789 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08961_ net621 _03896_ net258 vssd1 vssd1 vccd1 vccd1 _03900_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_65_Right_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07912_ _02850_ _02851_ _02862_ net879 vssd1 vssd1 vccd1 vccd1 _02863_ sky130_fd_sc_hd__a22oi_4
XANTENNA__12621__S _05080_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08892_ final_design.CPU_instr_adr\[27\] net1015 _03836_ _03838_ vssd1 vssd1 vccd1
+ vccd1 _00238_ sky130_fd_sc_hd__a22o_1
XANTENNA__06679__X _01630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12340__A2 net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07843_ final_design.cpu.reg_window\[533\] final_design.cpu.reg_window\[565\] net860
+ vssd1 vssd1 vccd1 vccd1 _02794_ sky130_fd_sc_hd__mux2_1
XANTENNA__10351__A1 net2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13941__CLK clknet_leaf_57_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07752__C1 _01626_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06839__B _01788_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout189_A _06045_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07774_ final_design.cpu.reg_window\[728\] final_design.cpu.reg_window\[760\] net862
+ vssd1 vssd1 vccd1 vccd1 _02725_ sky130_fd_sc_hd__mux2_1
X_09513_ _03025_ _04094_ vssd1 vssd1 vccd1 vccd1 _04432_ sky130_fd_sc_hd__nand2_1
XFILLER_0_71_1705 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06725_ final_design.cpu.reg_window\[920\] final_design.cpu.reg_window\[952\] net944
+ vssd1 vssd1 vccd1 vccd1 _01676_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_1885 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout356_A net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1098_A net1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1749 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06656_ final_design.cpu.reg_window\[218\] final_design.cpu.reg_window\[250\] net942
+ vssd1 vssd1 vccd1 vccd1 _01607_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09444_ net468 _04078_ _04102_ vssd1 vssd1 vccd1 vccd1 _04363_ sky130_fd_sc_hd__and3_1
XANTENNA__08546__S net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_74_Right_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09375_ net473 _04293_ vssd1 vssd1 vccd1 vccd1 _04294_ sky130_fd_sc_hd__nand2_1
X_06587_ net742 _01537_ net665 vssd1 vssd1 vccd1 vccd1 _01538_ sky130_fd_sc_hd__a21oi_4
XANTENNA_fanout523_A net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08326_ final_design.cpu.reg_window\[776\] final_design.cpu.reg_window\[808\] net816
+ vssd1 vssd1 vccd1 vccd1 _03277_ sky130_fd_sc_hd__mux2_1
X_14247__1301 vssd1 vssd1 vccd1 vccd1 _14247__1301/HI net1301 sky130_fd_sc_hd__conb_1
XANTENNA__10096__B net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13321__CLK clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08257_ final_design.cpu.reg_window\[10\] final_design.cpu.reg_window\[42\] net815
+ vssd1 vssd1 vccd1 vccd1 _03208_ sky130_fd_sc_hd__mux2_1
XANTENNA__09009__C1 net1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout311_X net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1053_X net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout409_X net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_3_5_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_3_5_0_clk sky130_fd_sc_hd__clkbuf_8
X_07208_ net536 _02157_ vssd1 vssd1 vccd1 vccd1 _02159_ sky130_fd_sc_hd__and2_1
XANTENNA__06590__A _01536_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08188_ final_design.cpu.reg_window\[398\] final_design.cpu.reg_window\[430\] net817
+ vssd1 vssd1 vccd1 vccd1 _03139_ sky130_fd_sc_hd__mux2_1
XANTENNA__10383__Y _05172_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout892_A net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07139_ _02084_ _02089_ net751 vssd1 vssd1 vccd1 vccd1 _02090_ sky130_fd_sc_hd__mux2_2
XFILLER_0_63_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13471__CLK clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_1889 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10150_ final_design.VGA_data_control.h_count\[0\] net1050 net1049 vssd1 vssd1 vccd1
+ vccd1 _05049_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout680_X net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout778_X net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10081_ _01400_ _04996_ _01391_ vssd1 vssd1 vccd1 vccd1 _04997_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_7_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12772__3 clknet_leaf_25_clk vssd1 vssd1 vccd1 vccd1 net1313 sky130_fd_sc_hd__inv_2
XANTENNA__09406__A _01493_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11655__B net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout945_X net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10342__B2 final_design.data_from_mem\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_2502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11147__S net245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13840_ clknet_leaf_33_clk _01071_ net1238 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[828\]
+ sky130_fd_sc_hd__dfrtp_1
X_13771_ clknet_leaf_53_clk _01002_ net1187 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[759\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10983_ _05690_ _05694_ _05709_ vssd1 vssd1 vccd1 vccd1 _05710_ sky130_fd_sc_hd__nand3_1
XANTENNA__08394__S0 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12722_ _06354_ _06362_ vssd1 vssd1 vccd1 vccd1 _06363_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_6_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06765__A net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12653_ final_design.VGA_data_control.ready_data\[14\] net1021 net976 final_design.data_from_mem\[14\]
+ vssd1 vssd1 vccd1 vccd1 _06314_ sky130_fd_sc_hd__a22o_1
XFILLER_0_2_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10287__A net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12398__A2 net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11604_ net671 _05848_ _06158_ vssd1 vssd1 vccd1 vccd1 _06159_ sky130_fd_sc_hd__or3_4
X_12584_ net2377 net998 net984 final_design.data_from_mem\[2\] vssd1 vssd1 vccd1 vccd1
+ _01277_ sky130_fd_sc_hd__a22o_1
XFILLER_0_19_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11535_ net1745 net176 net524 vssd1 vssd1 vccd1 vccd1 _00402_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_22_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13814__CLK clknet_leaf_59_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14254_ net1308 vssd1 vssd1 vccd1 vccd1 gpio_out[32] sky130_fd_sc_hd__buf_2
XANTENNA__08615__A_N _02211_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11466_ net215 net2460 net307 vssd1 vssd1 vccd1 vccd1 _00350_ sky130_fd_sc_hd__mux2_1
XANTENNA__11358__B1 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13205_ clknet_leaf_7_clk _00436_ net1134 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[193\]
+ sky130_fd_sc_hd__dfrtp_1
X_10417_ _03257_ _05190_ vssd1 vssd1 vccd1 vccd1 _05192_ sky130_fd_sc_hd__nor2_1
X_14185_ clknet_leaf_20_clk final_design.VGA_data_control.next_state\[1\] net1159
+ vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.state\[1\] sky130_fd_sc_hd__dfrtp_4
X_11397_ net649 net178 vssd1 vssd1 vccd1 vccd1 _06082_ sky130_fd_sc_hd__and2_1
XANTENNA__09566__A3 net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07121__S1 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13136_ clknet_leaf_34_clk _00367_ net1245 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[124\]
+ sky130_fd_sc_hd__dfrtp_1
X_10348_ wb_manage.curr_state\[1\] net1 vssd1 vssd1 vccd1 vccd1 _05169_ sky130_fd_sc_hd__nand2_1
XANTENNA__13964__CLK clknet_leaf_46_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08698__Y _03649_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08765__A_N final_design.CPU_instr_adr\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07982__C1 net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12441__S net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13067_ clknet_leaf_53_clk _00298_ net1188 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[55\]
+ sky130_fd_sc_hd__dfrtp_1
X_10279_ final_design.uart.BAUD_counter\[29\] final_design.uart.BAUD_counter\[28\]
+ _05134_ vssd1 vssd1 vccd1 vccd1 _05138_ sky130_fd_sc_hd__and3_1
XANTENNA__09723__A0 net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07535__S net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12018_ _06220_ net291 net403 net2257 vssd1 vssd1 vccd1 vccd1 _00749_ sky130_fd_sc_hd__a22o_1
XFILLER_0_40_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10333__B2 final_design.data_from_mem\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07107__Y _02058_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12086__A1 net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13969_ clknet_leaf_34_clk _01200_ net1242 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[957\]
+ sky130_fd_sc_hd__dfrtp_1
X_06510_ _01393_ net993 net990 final_design.reqhand.instruction\[6\] vssd1 vssd1 vccd1
+ vccd1 _01461_ sky130_fd_sc_hd__a31o_1
XFILLER_0_18_1566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07490_ _02439_ _02440_ vssd1 vssd1 vccd1 vccd1 _02441_ sky130_fd_sc_hd__nor2_1
XFILLER_0_53_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12396__B net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10909__B net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13344__CLK clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06441_ wb_manage.BUSY_O final_design.reqhand.current_client\[0\] net34 vssd1 vssd1
+ vccd1 vccd1 _01395_ sky130_fd_sc_hd__or3b_2
XFILLER_0_5_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1891 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09160_ net614 net525 _03523_ _01627_ vssd1 vssd1 vccd1 vccd1 _04079_ sky130_fd_sc_hd__a211o_1
XFILLER_0_1_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08111_ final_design.cpu.reg_window\[524\] final_design.cpu.reg_window\[556\] net812
+ vssd1 vssd1 vccd1 vccd1 _03062_ sky130_fd_sc_hd__mux2_1
XANTENNA__11597__B1 net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09091_ final_design.CPU_instr_adr\[3\] net1018 final_design.CPU_instr_adr\[4\] vssd1
+ vssd1 vccd1 vccd1 _04015_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12616__S _05080_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13494__CLK clknet_leaf_59_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11520__S net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08042_ net602 _02991_ _02966_ vssd1 vssd1 vccd1 vccd1 _02993_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_47_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11349__B1 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold901 final_design.cpu.reg_window\[575\] vssd1 vssd1 vccd1 vccd1 net2243 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkload43_A clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold912 final_design.cpu.reg_window\[1000\] vssd1 vssd1 vccd1 vccd1 net2254 sky130_fd_sc_hd__dlygate4sd3_1
Xhold923 final_design.cpu.reg_window\[1023\] vssd1 vssd1 vccd1 vccd1 net2265 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold934 final_design.cpu.reg_window\[547\] vssd1 vssd1 vccd1 vccd1 net2276 sky130_fd_sc_hd__dlygate4sd3_1
Xhold945 final_design.cpu.reg_window\[817\] vssd1 vssd1 vccd1 vccd1 net2287 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_874 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold956 final_design.cpu.reg_window\[431\] vssd1 vssd1 vccd1 vccd1 net2298 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap664 _01851_ vssd1 vssd1 vccd1 vccd1 net664 sky130_fd_sc_hd__buf_4
XANTENNA__12561__A2 net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold967 final_design.cpu.reg_window\[840\] vssd1 vssd1 vccd1 vccd1 net2309 sky130_fd_sc_hd__dlygate4sd3_1
Xhold978 final_design.cpu.reg_window\[892\] vssd1 vssd1 vccd1 vccd1 net2320 sky130_fd_sc_hd__dlygate4sd3_1
Xhold989 final_design.cpu.reg_window\[539\] vssd1 vssd1 vccd1 vccd1 net2331 sky130_fd_sc_hd__dlygate4sd3_1
X_09993_ net474 _04401_ vssd1 vssd1 vccd1 vccd1 _04912_ sky130_fd_sc_hd__or2_1
XFILLER_0_50_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08944_ _03882_ _03884_ net625 vssd1 vssd1 vccd1 vccd1 _03885_ sky130_fd_sc_hd__mux2_1
XANTENNA__07953__B net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1013_A net1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07445__S net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11475__B net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08875_ _01571_ _01601_ _02473_ net621 vssd1 vssd1 vccd1 vccd1 _03823_ sky130_fd_sc_hd__a31o_1
XANTENNA__10324__B2 final_design.data_from_mem\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout473_A net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07826_ final_design.cpu.reg_window\[21\] final_design.cpu.reg_window\[53\] net859
+ vssd1 vssd1 vccd1 vccd1 _02777_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout640_A _06093_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07757_ final_design.cpu.reg_window\[344\] final_design.cpu.reg_window\[376\] net864
+ vssd1 vssd1 vccd1 vccd1 _02708_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout261_X net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout738_A net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout359_X net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06708_ final_design.reqhand.instruction\[25\] final_design.data_from_mem\[25\] _01415_
+ vssd1 vssd1 vccd1 vccd1 _01659_ sky130_fd_sc_hd__mux2_4
X_07688_ net606 _02635_ _02611_ _01452_ vssd1 vssd1 vccd1 vccd1 _02639_ sky130_fd_sc_hd__o211a_1
X_09427_ _02900_ _04088_ _04344_ _04345_ vssd1 vssd1 vccd1 vccd1 _04346_ sky130_fd_sc_hd__o211a_1
X_06639_ final_design.cpu.reg_window\[731\] final_design.cpu.reg_window\[763\] net941
+ vssd1 vssd1 vccd1 vccd1 _01590_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout905_A net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_207 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13837__CLK clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09358_ _03484_ _04065_ vssd1 vssd1 vccd1 vccd1 _04277_ sky130_fd_sc_hd__nor2_1
XFILLER_0_75_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08309_ net610 _03257_ _03258_ net536 vssd1 vssd1 vccd1 vccd1 _03260_ sky130_fd_sc_hd__a211oi_2
X_09289_ _01566_ _01596_ net458 vssd1 vssd1 vccd1 vccd1 _04208_ sky130_fd_sc_hd__mux2_1
XANTENNA__11430__S net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11320_ final_design.data_from_mem\[21\] net235 net233 vssd1 vssd1 vccd1 vccd1 _06014_
+ sky130_fd_sc_hd__a21o_2
XFILLER_0_16_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12861__CLK clknet_leaf_17_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09564__A2_N net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13987__CLK clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11251_ final_design.data_from_mem\[13\] _05914_ _05917_ vssd1 vssd1 vccd1 vccd1
+ _05953_ sky130_fd_sc_hd__a21o_1
XFILLER_0_31_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10202_ final_design.uart.BAUD_counter_state _05078_ vssd1 vssd1 vccd1 vccd1 _05090_
+ sky130_fd_sc_hd__and2_1
XANTENNA__12552__A2 net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11182_ net660 _04006_ net732 vssd1 vssd1 vccd1 vccd1 _05892_ sky130_fd_sc_hd__o21a_1
X_10133_ final_design.VGA_data_control.h_count\[3\] net1048 final_design.VGA_data_control.h_count\[5\]
+ _05013_ vssd1 vssd1 vccd1 vccd1 _05037_ sky130_fd_sc_hd__nand4_1
XANTENNA__13217__CLK clknet_leaf_49_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06862__S0 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07355__S net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10064_ _04962_ _04963_ _04980_ _04982_ vssd1 vssd1 vccd1 vccd1 _04983_ sky130_fd_sc_hd__and4_1
XANTENNA_input34_A en vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10866__A2 net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13367__CLK clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09423__X _04342_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12068__A1 net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13823_ clknet_leaf_7_clk _01054_ net1134 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[811\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_8_1818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12497__A net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11605__S net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13754_ clknet_leaf_64_clk _00985_ net1074 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[742\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08186__S net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10966_ _05673_ _05692_ vssd1 vssd1 vccd1 vccd1 _05694_ sky130_fd_sc_hd__nand2_1
XFILLER_0_70_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12705_ net1051 _06344_ vssd1 vssd1 vccd1 vccd1 _06346_ sky130_fd_sc_hd__or2_1
XFILLER_0_70_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_14_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13685_ clknet_leaf_58_clk _00916_ net1144 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[673\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11291__A2 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10897_ _04356_ net252 vssd1 vssd1 vccd1 vccd1 _05627_ sky130_fd_sc_hd__nor2_1
XFILLER_0_35_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_974 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12636_ _06305_ net2421 net980 vssd1 vssd1 vccd1 vccd1 _01320_ sky130_fd_sc_hd__mux2_1
XANTENNA__11579__B1 net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12240__A1 net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12436__S net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12567_ net2013 _06288_ _06286_ vssd1 vssd1 vccd1 vccd1 _01268_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11518_ net576 _05980_ _06116_ vssd1 vssd1 vccd1 vccd1 _06121_ sky130_fd_sc_hd__and3_1
XANTENNA__10540__A_N net250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10464__B net250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12498_ net555 net631 _06268_ net327 net1561 vssd1 vssd1 vccd1 vccd1 _01203_ sky130_fd_sc_hd__a32o_1
Xhold208 final_design.cpu.reg_window\[731\] vssd1 vssd1 vccd1 vccd1 net1550 sky130_fd_sc_hd__dlygate4sd3_1
Xhold219 final_design.cpu.reg_window\[960\] vssd1 vssd1 vccd1 vccd1 net1561 sky130_fd_sc_hd__dlygate4sd3_1
X_14237_ net1291 vssd1 vssd1 vccd1 vccd1 gpio_out[15] sky130_fd_sc_hd__buf_2
X_11449_ net242 net2382 net307 vssd1 vssd1 vccd1 vccd1 _00341_ sky130_fd_sc_hd__mux2_1
XANTENNA__09539__A3 _01784_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1873 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_1715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12543__A2 net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14168_ clknet_leaf_18_clk _01342_ net1108 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.data_to_VGA\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10554__A1 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11751__A0 net206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10554__B2 net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13119_ clknet_leaf_8_clk _00350_ net1154 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[107\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14142__CLK clknet_leaf_19_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12171__S net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14099_ clknet_leaf_14_clk _01296_ net1111 vssd1 vssd1 vccd1 vccd1 final_design.reqhand.instruction\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_06990_ _01937_ _01939_ vssd1 vssd1 vccd1 vccd1 _01941_ sky130_fd_sc_hd__nand2_1
XANTENNA__07265__S net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14246__1300 vssd1 vssd1 vccd1 vccd1 _14246__1300/HI net1300 sky130_fd_sc_hd__conb_1
XFILLER_0_56_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_1988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13759__RESET_B net1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08660_ _02542_ _03610_ vssd1 vssd1 vccd1 vccd1 _03611_ sky130_fd_sc_hd__and2b_1
XANTENNA__06957__X _01908_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07611_ final_design.cpu.reg_window\[669\] final_design.cpu.reg_window\[701\] net870
+ vssd1 vssd1 vccd1 vccd1 _02562_ sky130_fd_sc_hd__mux2_1
X_08591_ net709 _03541_ vssd1 vssd1 vccd1 vccd1 _03542_ sky130_fd_sc_hd__or2_1
XANTENNA__06930__B1 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1833 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11515__S net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07542_ final_design.cpu.reg_window\[927\] final_design.cpu.reg_window\[959\] net947
+ vssd1 vssd1 vccd1 vccd1 _02493_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_1877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07473_ net741 _01497_ _02420_ _02421_ vssd1 vssd1 vccd1 vccd1 _02424_ sky130_fd_sc_hd__a211oi_4
XTAP_TAPCELL_ROW_27_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_46_Left_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09212_ _04130_ vssd1 vssd1 vccd1 vccd1 _04131_ sky130_fd_sc_hd__inv_2
XANTENNA__10490__B1 net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06424_ final_design.data_from_mem\[5\] vssd1 vssd1 vccd1 vccd1 _01379_ sky130_fd_sc_hd__inv_2
XANTENNA__07581__S1 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12884__CLK clknet_leaf_15_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12786__17 clknet_leaf_27_clk vssd1 vssd1 vccd1 vccd1 net1327 sky130_fd_sc_hd__inv_2
X_09143_ net460 _03553_ _04061_ vssd1 vssd1 vccd1 vccd1 _04062_ sky130_fd_sc_hd__or3_1
XFILLER_0_16_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout221_A _05921_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09074_ _03702_ _03722_ vssd1 vssd1 vccd1 vccd1 _04000_ sky130_fd_sc_hd__or2_1
XFILLER_0_60_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08025_ final_design.cpu.reg_window\[147\] final_design.cpu.reg_window\[179\] net830
+ vssd1 vssd1 vccd1 vccd1 _02976_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_9_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_1913 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1350 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold720 final_design.cpu.reg_window\[926\] vssd1 vssd1 vccd1 vccd1 net2062 sky130_fd_sc_hd__dlygate4sd3_1
Xhold731 final_design.cpu.reg_window\[849\] vssd1 vssd1 vccd1 vccd1 net2073 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold742 final_design.cpu.reg_window\[425\] vssd1 vssd1 vccd1 vccd1 net2084 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1228_A net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold753 final_design.cpu.reg_window\[967\] vssd1 vssd1 vccd1 vccd1 net2095 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12534__A2 net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold764 final_design.cpu.reg_window\[687\] vssd1 vssd1 vccd1 vccd1 net2106 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout590_A net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold775 final_design.cpu.reg_window\[693\] vssd1 vssd1 vccd1 vccd1 net2117 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_55_Left_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout688_A net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold786 final_design.cpu.reg_window\[901\] vssd1 vssd1 vccd1 vccd1 net2128 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07946__C1 _01750_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold797 final_design.cpu.reg_window\[653\] vssd1 vssd1 vccd1 vccd1 net2139 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07410__A1 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06844__S0 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09976_ _03358_ _04720_ _03565_ vssd1 vssd1 vccd1 vccd1 _04895_ sky130_fd_sc_hd__a21o_1
X_08927_ _03869_ vssd1 vssd1 vccd1 vccd1 _03870_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout855_A net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09163__A1 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout476_X net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08858_ net624 _03807_ vssd1 vssd1 vccd1 vccd1 _03808_ sky130_fd_sc_hd__nor2_1
XANTENNA__08910__A1 net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07809_ final_design.cpu.reg_window\[537\] final_design.cpu.reg_window\[569\] net851
+ vssd1 vssd1 vccd1 vccd1 _02760_ sky130_fd_sc_hd__mux2_1
XANTENNA__13429__RESET_B net1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08789_ _03683_ _03686_ _03736_ _03739_ vssd1 vssd1 vccd1 vccd1 _03740_ sky130_fd_sc_hd__and4_1
XANTENNA_fanout643_X net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11425__S net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10820_ _01362_ _03909_ net1060 vssd1 vssd1 vccd1 vccd1 _05554_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_64_Left_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_1917 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10751_ net74 _05466_ _05487_ vssd1 vssd1 vccd1 vccd1 _05488_ sky130_fd_sc_hd__a21o_1
XFILLER_0_7_1873 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10481__B1 net1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13470_ clknet_leaf_9_clk _00701_ net1099 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[458\]
+ sky130_fd_sc_hd__dfrtp_1
X_10682_ _05421_ _05422_ vssd1 vssd1 vccd1 vccd1 _05423_ sky130_fd_sc_hd__xnor2_1
XANTENNA__14015__CLK clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12421_ _06244_ net501 net340 net2149 vssd1 vssd1 vccd1 vccd1 _01130_ sky130_fd_sc_hd__a22o_1
XANTENNA__12222__A1 net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07324__S1 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12352_ net2502 net362 net354 _06018_ vssd1 vssd1 vccd1 vccd1 _01064_ sky130_fd_sc_hd__a22o_1
XANTENNA__06988__B1 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11981__B1 net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11303_ net660 _03896_ net733 vssd1 vssd1 vccd1 vccd1 _05999_ sky130_fd_sc_hd__o21ai_1
XANTENNA__14165__CLK clknet_leaf_18_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12283_ net567 _06213_ net506 net369 net1799 vssd1 vssd1 vccd1 vccd1 _00998_ sky130_fd_sc_hd__a32o_1
XPHY_EDGE_ROW_73_Left_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_660 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14022_ clknet_leaf_51_clk _01253_ net1173 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[1010\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12525__A2 net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11234_ net732 _03965_ vssd1 vssd1 vccd1 vccd1 _05938_ sky130_fd_sc_hd__or2_1
X_11165_ net804 _05846_ vssd1 vssd1 vccd1 vccd1 _05877_ sky130_fd_sc_hd__nor2_4
XANTENNA__07085__S net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10116_ _05026_ vssd1 vssd1 vccd1 vccd1 _05027_ sky130_fd_sc_hd__inv_2
X_11096_ net1585 net1034 _05816_ _05817_ vssd1 vssd1 vccd1 vccd1 _00203_ sky130_fd_sc_hd__a22o_1
XANTENNA__12289__A1 net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1191 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10047_ _04577_ _04598_ _04925_ _04965_ vssd1 vssd1 vccd1 vccd1 _04966_ sky130_fd_sc_hd__a211oi_1
Xhold80 net164 vssd1 vssd1 vccd1 vccd1 net1422 sky130_fd_sc_hd__dlygate4sd3_1
Xhold91 net119 vssd1 vssd1 vccd1 vccd1 net1433 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11843__B net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_82_Left_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_19_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13806_ clknet_leaf_45_clk _01037_ net1216 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[794\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_19_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12801__32_A clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11998_ _06200_ net280 net401 net2501 vssd1 vssd1 vccd1 vccd1 _00729_ sky130_fd_sc_hd__a22o_1
XFILLER_0_19_1683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07114__A _02059_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13737_ clknet_leaf_36_clk _00968_ net1229 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[725\]
+ sky130_fd_sc_hd__dfrtp_1
X_10949_ net84 net1046 vssd1 vssd1 vccd1 vccd1 _05677_ sky130_fd_sc_hd__nand2_1
XANTENNA__11264__A2 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07468__B2 net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10472__B1 _04990_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13668_ clknet_leaf_54_clk _00899_ net1180 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[656\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_41_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12213__A1 net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12619_ final_design.uart.working_data\[6\] net2547 _05080_ vssd1 vssd1 vccd1 vccd1
+ _01312_ sky130_fd_sc_hd__mux2_1
XANTENNA__12166__S net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13599_ clknet_leaf_4_clk _00830_ net1084 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[587\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11972__B1 net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12516__A2 net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07784__A net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_39_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13532__CLK clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11724__B1 net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09830_ _04182_ _04745_ _04746_ vssd1 vssd1 vccd1 vccd1 _04749_ sky130_fd_sc_hd__and3_1
Xfanout507 net516 vssd1 vssd1 vccd1 vccd1 net507 sky130_fd_sc_hd__buf_4
Xfanout518 net520 vssd1 vssd1 vccd1 vccd1 net518 sky130_fd_sc_hd__buf_4
Xfanout529 _02294_ vssd1 vssd1 vccd1 vccd1 net529 sky130_fd_sc_hd__clkbuf_2
X_09761_ _04143_ _04157_ _03590_ vssd1 vssd1 vccd1 vccd1 _04680_ sky130_fd_sc_hd__o21ai_1
X_06973_ net756 _01917_ net747 vssd1 vssd1 vccd1 vccd1 _01924_ sky130_fd_sc_hd__o21a_1
XFILLER_0_20_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08712_ final_design.CPU_instr_adr\[26\] _01630_ vssd1 vssd1 vccd1 vccd1 _03663_
+ sky130_fd_sc_hd__or2_1
XANTENNA__13682__CLK clknet_leaf_38_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09692_ _03071_ _03102_ _04496_ _03581_ _03165_ vssd1 vssd1 vccd1 vccd1 _04611_ sky130_fd_sc_hd__a311o_1
XFILLER_0_59_1463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08643_ _02903_ net260 _03592_ _03040_ vssd1 vssd1 vccd1 vccd1 _03594_ sky130_fd_sc_hd__o31ai_4
XTAP_TAPCELL_ROW_1_236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout269_A net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08574_ final_design.cpu.reg_window\[320\] final_design.cpu.reg_window\[352\] net827
+ vssd1 vssd1 vccd1 vccd1 _03525_ sky130_fd_sc_hd__mux2_1
XANTENNA__14038__CLK clknet_leaf_15_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07525_ _01540_ _02475_ _01541_ vssd1 vssd1 vccd1 vccd1 _02476_ sky130_fd_sc_hd__a21bo_1
XANTENNA__12452__A1 net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11255__A2 _05953_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1080_A net1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_61_clk clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_61_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout436_A net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1178_A net1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07456_ net750 _02400_ net745 vssd1 vssd1 vccd1 vccd1 _02407_ sky130_fd_sc_hd__o21a_1
XFILLER_0_8_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06407_ final_design.CPU_instr_adr\[18\] vssd1 vssd1 vccd1 vccd1 _01362_ sky130_fd_sc_hd__inv_2
XANTENNA__13062__CLK clknet_leaf_51_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07387_ final_design.cpu.reg_window\[66\] final_design.cpu.reg_window\[98\] net918
+ vssd1 vssd1 vccd1 vccd1 _02338_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout224_X net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout603_A net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09126_ _03631_ _03647_ vssd1 vssd1 vccd1 vccd1 _04045_ sky130_fd_sc_hd__nor2_2
XFILLER_0_44_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11963__B1 net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09057_ _02441_ net620 _03984_ vssd1 vssd1 vccd1 vccd1 _03985_ sky130_fd_sc_hd__or3_1
XANTENNA__12507__A2 net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08008_ _02955_ _02956_ _02957_ _02958_ net682 net693 vssd1 vssd1 vccd1 vccd1 _02959_
+ sky130_fd_sc_hd__mux4_1
Xhold550 final_design.cpu.reg_window\[798\] vssd1 vssd1 vccd1 vccd1 net1892 sky130_fd_sc_hd__dlygate4sd3_1
Xhold561 final_design.cpu.reg_window\[883\] vssd1 vssd1 vccd1 vccd1 net1903 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout593_X net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout972_A _01415_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold572 final_design.cpu.reg_window\[671\] vssd1 vssd1 vccd1 vccd1 net1914 sky130_fd_sc_hd__dlygate4sd3_1
Xhold583 final_design.cpu.reg_window\[520\] vssd1 vssd1 vccd1 vccd1 net1925 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09384__A1 net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11647__C net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold594 final_design.cpu.reg_window\[64\] vssd1 vssd1 vccd1 vccd1 net1936 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11191__A1 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_1817 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_2586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout760_X net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_2597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09959_ net447 _04877_ vssd1 vssd1 vccd1 vccd1 _04878_ sky130_fd_sc_hd__nor2_1
X_12970_ clknet_leaf_15_clk _00208_ net1092 vssd1 vssd1 vccd1 vccd1 final_design.uart.bits_received\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_77_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09687__A2 net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07633__S net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11921_ net673 _06118_ _06124_ vssd1 vssd1 vccd1 vccd1 _06252_ sky130_fd_sc_hd__or3_1
XANTENNA__11663__B net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07793__S1 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11852_ _06102_ net277 net517 net2034 vssd1 vssd1 vccd1 vccd1 _00602_ sky130_fd_sc_hd__a22o_1
XFILLER_0_79_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10803_ net802 _05535_ _05537_ net962 vssd1 vssd1 vccd1 vccd1 _05538_ sky130_fd_sc_hd__o22a_1
XFILLER_0_55_1894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_64_2379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11246__A2 _05943_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11783_ net2412 net412 net278 _05935_ vssd1 vssd1 vccd1 vccd1 _00541_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_52_clk clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_52_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_55_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13405__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1889 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13522_ clknet_leaf_39_clk _00753_ net1205 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[510\]
+ sky130_fd_sc_hd__dfrtp_1
X_10734_ _01364_ _03940_ net1060 vssd1 vssd1 vccd1 vccd1 _05472_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_1534 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13453_ clknet_leaf_44_clk _00684_ net1201 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[441\]
+ sky130_fd_sc_hd__dfrtp_1
X_10665_ _04677_ net253 _04990_ vssd1 vssd1 vccd1 vccd1 _05406_ sky130_fd_sc_hd__o21ai_1
XANTENNA__12781__12_A clknet_leaf_28_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12404_ _06102_ net343 net338 net2269 vssd1 vssd1 vccd1 vccd1 _01114_ sky130_fd_sc_hd__a22o_1
XFILLER_0_63_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13384_ clknet_leaf_41_clk _00615_ net1225 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[372\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_63_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10596_ final_design.CPU_instr_adr\[7\] net1001 _05338_ net1042 vssd1 vssd1 vccd1
+ vccd1 _05341_ sky130_fd_sc_hd__o22a_1
XANTENNA__13555__CLK clknet_leaf_38_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10757__B2 net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11954__B1 net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12335_ net2338 net360 net343 _05891_ vssd1 vssd1 vccd1 vccd1 _01047_ sky130_fd_sc_hd__a22o_1
XANTENNA__11001__A1_N net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_1821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06712__S net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12266_ _06196_ net506 net369 net2026 vssd1 vssd1 vccd1 vccd1 _00981_ sky130_fd_sc_hd__a22o_1
XANTENNA__11706__B1 net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14005_ clknet_leaf_57_clk _01236_ net1144 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[993\]
+ sky130_fd_sc_hd__dfrtp_1
X_11217_ net662 _03976_ net735 vssd1 vssd1 vccd1 vccd1 _05923_ sky130_fd_sc_hd__a21o_1
X_12197_ net231 net2428 net376 vssd1 vssd1 vccd1 vccd1 _00915_ sky130_fd_sc_hd__mux2_1
XANTENNA__11182__A1 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07109__A final_design.data_from_mem\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11148_ _05855_ _05861_ vssd1 vssd1 vccd1 vccd1 _05862_ sky130_fd_sc_hd__nand2_1
XFILLER_0_78_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11079_ _05765_ _05779_ _05800_ vssd1 vssd1 vccd1 vccd1 _05801_ sky130_fd_sc_hd__a21o_1
XANTENNA__12131__A0 net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11065__S net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09395__A2_N _04087_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1311 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13085__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12986__RESET_B net1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09835__C1 net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_43_clk clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_43_clk sky130_fd_sc_hd__clkbuf_8
X_07310_ final_design.cpu.reg_window\[517\] final_design.cpu.reg_window\[549\] net923
+ vssd1 vssd1 vccd1 vccd1 _02261_ sky130_fd_sc_hd__mux2_1
XANTENNA__07536__S1 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08290_ final_design.cpu.reg_window\[201\] final_design.cpu.reg_window\[233\] net808
+ vssd1 vssd1 vccd1 vccd1 _03241_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_9_clk_A clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14139__RESET_B net1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07241_ _02188_ _02189_ _02190_ _02191_ net764 net780 vssd1 vssd1 vccd1 vccd1 _02192_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__12198__B1 net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07172_ final_design.cpu.reg_window\[522\] final_design.cpu.reg_window\[554\] net895
+ vssd1 vssd1 vccd1 vccd1 _02123_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11945__B1 net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12922__CLK clknet_leaf_61_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06622__S net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1039 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout304 net305 vssd1 vssd1 vccd1 vccd1 net304 sky130_fd_sc_hd__buf_4
Xfanout315 _05851_ vssd1 vssd1 vccd1 vccd1 net315 sky130_fd_sc_hd__buf_4
Xfanout326 net327 vssd1 vssd1 vccd1 vccd1 net326 sky130_fd_sc_hd__buf_4
X_09813_ net539 net538 net537 net535 net452 net461 vssd1 vssd1 vccd1 vccd1 _04732_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__07916__A2 _02863_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout337 _06282_ vssd1 vssd1 vccd1 vccd1 net337 sky130_fd_sc_hd__buf_8
XANTENNA__07019__A net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout348 net350 vssd1 vssd1 vccd1 vccd1 net348 sky130_fd_sc_hd__clkbuf_4
Xfanout359 _06277_ vssd1 vssd1 vccd1 vccd1 net359 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout386_A net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09744_ net541 net540 net539 _02091_ net455 net464 vssd1 vssd1 vccd1 vccd1 _04663_
+ sky130_fd_sc_hd__mux4_1
X_06956_ _01901_ _01906_ net756 vssd1 vssd1 vccd1 vccd1 _01907_ sky130_fd_sc_hd__mux2_1
XANTENNA__11483__B net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09675_ _04592_ _04593_ _04590_ vssd1 vssd1 vccd1 vccd1 _04594_ sky130_fd_sc_hd__o21ai_2
XANTENNA__12673__B2 final_design.data_from_mem\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06887_ final_design.cpu.reg_window\[851\] final_design.cpu.reg_window\[883\] net911
+ vssd1 vssd1 vccd1 vccd1 _01838_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout553_A _06238_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13428__CLK clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08341__A2 _03287_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08626_ _03231_ _03576_ vssd1 vssd1 vccd1 vccd1 _03577_ sky130_fd_sc_hd__nand2_1
XFILLER_0_33_1411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11770__Y _06228_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09888__B net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11228__A2 _05930_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08557_ final_design.cpu.reg_window\[641\] final_design.cpu.reg_window\[673\] net834
+ vssd1 vssd1 vccd1 vccd1 _03508_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout720_A net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout341_X net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_7_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout818_A net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout439_X net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_34_clk clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_34_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_82_2991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_1821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07508_ _01884_ _02457_ _01882_ vssd1 vssd1 vccd1 vccd1 _02459_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11930__C net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08488_ final_design.cpu.reg_window\[835\] final_design.cpu.reg_window\[867\] net831
+ vssd1 vssd1 vccd1 vccd1 _03439_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13578__CLK clknet_leaf_60_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07439_ net883 _02382_ _02388_ _02375_ _02376_ vssd1 vssd1 vccd1 vccd1 _02390_ sky130_fd_sc_hd__a32o_1
XFILLER_0_80_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10450_ _02763_ net592 vssd1 vssd1 vccd1 vccd1 _05209_ sky130_fd_sc_hd__or2_1
XFILLER_0_66_1220 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11936__B1 net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09109_ net619 _04028_ _04029_ _02428_ vssd1 vssd1 vccd1 vccd1 _04030_ sky130_fd_sc_hd__a22o_1
X_10381_ net25 net1026 net1008 final_design.data_from_mem\[30\] vssd1 vssd1 vccd1
+ vccd1 _00134_ sky130_fd_sc_hd__a22o_1
XFILLER_0_81_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_57_2150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_76_2784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12120_ net1915 net188 net390 vssd1 vssd1 vccd1 vccd1 _00844_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_57_2161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_76_2795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_2003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_2014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_2025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12051_ net1949 net190 net399 vssd1 vssd1 vccd1 vccd1 _00779_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold380 final_design.cpu.reg_window\[63\] vssd1 vssd1 vccd1 vccd1 net1722 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09128__B _04045_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold391 final_design.cpu.reg_window\[603\] vssd1 vssd1 vccd1 vccd1 net1733 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11164__B2 net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12361__B1 net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11002_ net670 _05714_ _05727_ net966 _05726_ vssd1 vssd1 vccd1 vccd1 _05728_ sky130_fd_sc_hd__o221a_1
XFILLER_0_79_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08600__X _03551_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10989__S net1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout860 net872 vssd1 vssd1 vccd1 vccd1 net860 sky130_fd_sc_hd__clkbuf_4
Xfanout871 net872 vssd1 vssd1 vccd1 vccd1 net871 sky130_fd_sc_hd__buf_2
XANTENNA__09415__Y _04334_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout882 net883 vssd1 vssd1 vccd1 vccd1 net882 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_5_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout893 net894 vssd1 vssd1 vccd1 vccd1 net893 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_5_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07363__S net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12953_ clknet_leaf_29_clk _00191_ net1195 vssd1 vssd1 vccd1 vccd1 net110 sky130_fd_sc_hd__dfrtp_1
Xhold1080 final_design.cpu.reg_window\[864\] vssd1 vssd1 vccd1 vccd1 net2422 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1091 final_design.cpu.reg_window\[437\] vssd1 vssd1 vccd1 vccd1 net2433 sky130_fd_sc_hd__dlygate4sd3_1
X_11904_ net200 net2129 net273 vssd1 vssd1 vccd1 vccd1 _00646_ sky130_fd_sc_hd__mux2_1
XANTENNA__07766__S1 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12884_ clknet_leaf_15_clk _00122_ net1094 vssd1 vssd1 vccd1 vccd1 final_design.data_from_mem\[18\]
+ sky130_fd_sc_hd__dfrtp_4
X_11835_ net191 net1981 net266 vssd1 vssd1 vccd1 vccd1 _00587_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_25_clk clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_25_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__09150__Y _04069_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11766_ net178 net2177 net418 vssd1 vssd1 vccd1 vccd1 _00529_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_1528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13505_ clknet_leaf_49_clk _00736_ net1186 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[493\]
+ sky130_fd_sc_hd__dfrtp_1
X_10717_ net669 _05444_ _05455_ vssd1 vssd1 vccd1 vccd1 _05456_ sky130_fd_sc_hd__o21a_1
X_11697_ net209 net628 vssd1 vssd1 vccd1 vccd1 _06207_ sky130_fd_sc_hd__and2_1
XANTENNA__12945__CLK clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13436_ clknet_leaf_5_clk _00667_ net1077 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[424\]
+ sky130_fd_sc_hd__dfrtp_1
X_10648_ net69 final_design.VGA_adr\[8\] vssd1 vssd1 vccd1 vccd1 _05390_ sky130_fd_sc_hd__xor2_1
XFILLER_0_67_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13367_ clknet_leaf_6_clk _00598_ net1132 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[355\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12444__S net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10579_ net64 _05324_ vssd1 vssd1 vccd1 vccd1 _05325_ sky130_fd_sc_hd__and2_1
XANTENNA__14225__A final_design.cpu.Error vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12318_ net2258 net196 net366 vssd1 vssd1 vccd1 vccd1 _01032_ sky130_fd_sc_hd__mux2_1
XANTENNA__11568__B net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13298_ clknet_leaf_38_clk _00529_ net1190 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[286\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_1782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12249_ net572 _06178_ net508 net375 net1536 vssd1 vssd1 vccd1 vccd1 _00965_ sky130_fd_sc_hd__a32o_1
XFILLER_0_43_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12352__B1 net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07454__S0 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06810_ final_design.cpu.reg_window\[149\] final_design.cpu.reg_window\[181\] net937
+ vssd1 vssd1 vccd1 vccd1 _01761_ sky130_fd_sc_hd__mux2_1
XANTENNA__08369__S net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07790_ final_design.cpu.reg_window\[281\] final_design.cpu.reg_window\[313\] net856
+ vssd1 vssd1 vccd1 vccd1 _02741_ sky130_fd_sc_hd__mux2_1
XANTENNA__08308__C1 net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06678__A net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06741_ _01686_ _01690_ vssd1 vssd1 vccd1 vccd1 _01692_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_79_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12655__B2 final_design.data_from_mem\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09460_ net320 _04373_ _04378_ _04117_ _04375_ vssd1 vssd1 vccd1 vccd1 _04379_ sky130_fd_sc_hd__a221o_1
X_06672_ final_design.cpu.reg_window\[666\] final_design.cpu.reg_window\[698\] net941
+ vssd1 vssd1 vccd1 vccd1 _01623_ sky130_fd_sc_hd__mux2_1
X_08411_ final_design.cpu.reg_window\[261\] final_design.cpu.reg_window\[293\] net840
+ vssd1 vssd1 vccd1 vccd1 _03362_ sky130_fd_sc_hd__mux2_1
XANTENNA__13720__CLK clknet_leaf_65_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09391_ net485 _04309_ _04306_ vssd1 vssd1 vccd1 vccd1 _04310_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_73_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12619__S _05080_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_16_clk clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_16_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__11523__S net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08342_ _03290_ _03292_ vssd1 vssd1 vccd1 vccd1 _03293_ sky130_fd_sc_hd__nor2_1
XANTENNA__06617__S net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1805 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07834__A1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08273_ net874 _03223_ _03212_ _03206_ vssd1 vssd1 vccd1 vccd1 _03224_ sky130_fd_sc_hd__o2bb2a_4
XFILLER_0_69_1849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13870__CLK clknet_leaf_45_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07224_ final_design.cpu.reg_window\[520\] final_design.cpu.reg_window\[552\] net888
+ vssd1 vssd1 vccd1 vccd1 _02175_ sky130_fd_sc_hd__mux2_1
X_07155_ _02102_ _02103_ _02104_ _02105_ net765 net780 vssd1 vssd1 vccd1 vccd1 _02106_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout301_A _06159_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1043_A final_design.VGA_adr\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11394__A1 _01507_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11394__B2 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12591__B1 net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13100__CLK clknet_leaf_46_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11478__B net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07086_ final_design.cpu.reg_window\[396\] final_design.cpu.reg_window\[428\] net906
+ vssd1 vssd1 vccd1 vccd1 _02037_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1210_A net1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11146__A1 final_design.CPU_instr_adr\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12343__B1 net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09516__X _04435_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout291_X net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout768_A net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout389_X net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07996__S1 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13250__CLK clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout178 _06081_ vssd1 vssd1 vccd1 vccd1 net178 sky130_fd_sc_hd__buf_2
X_07988_ final_design.cpu.reg_window\[272\] final_design.cpu.reg_window\[304\] net846
+ vssd1 vssd1 vccd1 vccd1 _02939_ sky130_fd_sc_hd__mux2_1
Xfanout189 _06045_ vssd1 vssd1 vccd1 vccd1 net189 sky130_fd_sc_hd__clkbuf_2
X_09727_ _04644_ _04645_ net477 vssd1 vssd1 vccd1 vccd1 _04646_ sky130_fd_sc_hd__mux2_2
X_06939_ final_design.cpu.reg_window\[81\] final_design.cpu.reg_window\[113\] net928
+ vssd1 vssd1 vccd1 vccd1 _01890_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout935_A net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09899__A net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09658_ _04576_ vssd1 vssd1 vccd1 vccd1 _04577_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_65_2430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_2441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_54_clk_X clknet_leaf_54_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07911__S net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08609_ _03559_ vssd1 vssd1 vccd1 vccd1 _03560_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_80_2928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_2305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout723_X net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10397__X _05181_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09589_ _03134_ _04506_ _04507_ vssd1 vssd1 vccd1 vccd1 _04508_ sky130_fd_sc_hd__a21o_2
XANTENNA__11433__S net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12968__CLK clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11620_ net558 net420 _06167_ net298 net1446 vssd1 vssd1 vccd1 vccd1 _00442_ sky130_fd_sc_hd__a32o_1
XFILLER_0_4_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11551_ net564 net421 _06131_ net303 net1772 vssd1 vssd1 vccd1 vccd1 _00409_ sky130_fd_sc_hd__a32o_1
XFILLER_0_64_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10502_ net93 final_design.VGA_adr\[1\] vssd1 vssd1 vccd1 vccd1 _05251_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_59_2212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11482_ net192 net2355 net309 vssd1 vssd1 vccd1 vccd1 _00362_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_59_2223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_2857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_2234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_2868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13221_ clknet_leaf_49_clk _00452_ net1181 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[209\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_78_2879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10433_ net1927 net1034 _05200_ net248 vssd1 vssd1 vccd1 vccd1 _00157_ sky130_fd_sc_hd__a22o_1
XANTENNA__11669__A net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12264__S net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11385__A1 final_design.data_from_mem\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12582__B1 net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input64_A mem_adr_start[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13152_ clknet_leaf_12_clk _00383_ net1090 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[140\]
+ sky130_fd_sc_hd__dfrtp_1
X_10364_ net6 net1024 net1007 final_design.data_from_mem\[13\] vssd1 vssd1 vccd1 vccd1
+ _00117_ sky130_fd_sc_hd__o22a_1
X_12103_ net1579 net220 net388 vssd1 vssd1 vccd1 vccd1 _00827_ sky130_fd_sc_hd__mux2_1
XANTENNA__11956__X _06255_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13083_ clknet_leaf_0_clk _00314_ net1061 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[71\]
+ sky130_fd_sc_hd__dfrtp_1
X_10295_ final_design.VGA_data_control.h_count\[2\] _05148_ vssd1 vssd1 vccd1 vccd1
+ _05149_ sky130_fd_sc_hd__and2b_1
XANTENNA__11137__A1 final_design.CPU_instr_adr\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12334__B1 net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1212 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12034_ net1893 net243 net396 vssd1 vssd1 vccd1 vccd1 _00762_ sky130_fd_sc_hd__mux2_1
XANTENNA__07436__S0 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_1466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10360__A2 net1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout690 _01787_ vssd1 vssd1 vccd1 vccd1 net690 sky130_fd_sc_hd__buf_4
XANTENNA__13743__CLK clknet_leaf_43_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13985_ clknet_leaf_47_clk _01216_ net1198 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[973\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12637__B2 final_design.data_from_mem\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12936_ clknet_leaf_22_clk _00174_ net1165 vssd1 vssd1 vccd1 vccd1 net112 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12439__S net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12867_ clknet_leaf_25_clk _00105_ net1151 vssd1 vssd1 vccd1 vccd1 final_design.data_from_mem\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__11860__A2 net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13893__CLK clknet_leaf_52_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11818_ net244 net2041 net264 vssd1 vssd1 vccd1 vccd1 _00570_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08164__S1 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11749_ net209 net2050 net418 vssd1 vssd1 vccd1 vccd1 _00512_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_1347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11612__A2 net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09281__A3 net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13123__CLK clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06961__A _01908_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13419_ clknet_leaf_38_clk _00650_ net1190 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[407\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12174__S net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11376__A1 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06680__B _01630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_1708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08241__B2 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13273__CLK clknet_leaf_55_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08960_ net625 _03898_ vssd1 vssd1 vccd1 vccd1 _03899_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_5_clk clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_5_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_45_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07911_ _02856_ _02861_ net714 vssd1 vssd1 vccd1 vccd1 _02862_ sky130_fd_sc_hd__mux2_1
X_08891_ net257 _03837_ net1015 vssd1 vssd1 vccd1 vccd1 _03838_ sky130_fd_sc_hd__a21oi_1
X_07842_ final_design.cpu.reg_window\[597\] final_design.cpu.reg_window\[629\] net857
+ vssd1 vssd1 vccd1 vccd1 _02793_ sky130_fd_sc_hd__mux2_1
XANTENNA__10351__A2 net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07773_ _02720_ _02721_ _02722_ _02723_ net686 net704 vssd1 vssd1 vccd1 vccd1 _02724_
+ sky130_fd_sc_hd__mux4_1
X_09512_ _02965_ _03028_ _04351_ vssd1 vssd1 vccd1 vccd1 _04431_ sky130_fd_sc_hd__and3_1
X_06724_ final_design.cpu.reg_window\[984\] final_design.cpu.reg_window\[1016\] net944
+ vssd1 vssd1 vccd1 vccd1 _01675_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_758 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1717 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07731__S net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09443_ net463 _04079_ _04081_ vssd1 vssd1 vccd1 vccd1 _04362_ sky130_fd_sc_hd__and3_1
X_06655_ _01602_ _01603_ _01604_ _01605_ net775 net793 vssd1 vssd1 vccd1 vccd1 _01606_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout251_A _04961_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11851__A2 net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_920 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout349_A net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09374_ net462 _04103_ _04257_ vssd1 vssd1 vccd1 vccd1 _04293_ sky130_fd_sc_hd__and3_1
X_06586_ final_design.reqhand.instruction\[29\] final_design.data_from_mem\[29\] net973
+ vssd1 vssd1 vccd1 vccd1 _01537_ sky130_fd_sc_hd__mux2_4
XFILLER_0_30_1403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08325_ final_design.cpu.reg_window\[840\] final_design.cpu.reg_window\[872\] net817
+ vssd1 vssd1 vccd1 vccd1 _03276_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout1160_A net1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10811__B1 net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08256_ final_design.cpu.reg_window\[74\] final_design.cpu.reg_window\[106\] net817
+ vssd1 vssd1 vccd1 vccd1 _03207_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07207_ net535 _02157_ vssd1 vssd1 vccd1 vccd1 _02158_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout304_X net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08187_ final_design.cpu.reg_window\[462\] final_design.cpu.reg_window\[494\] net816
+ vssd1 vssd1 vccd1 vccd1 _03138_ sky130_fd_sc_hd__mux2_1
XANTENNA__11367__A1 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06590__B _01539_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13616__CLK clknet_leaf_36_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_2710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07138_ _02085_ _02086_ _02087_ _02088_ net768 net781 vssd1 vssd1 vccd1 vccd1 _02089_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_30_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout885_A net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07069_ final_design.cpu.reg_window\[845\] final_design.cpu.reg_window\[877\] net935
+ vssd1 vssd1 vccd1 vccd1 _02020_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_7_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10080_ final_design.VGA_data_control.v_count\[2\] final_design.VGA_data_control.v_count\[1\]
+ final_design.VGA_data_control.v_count\[3\] vssd1 vssd1 vccd1 vccd1 _04996_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_7_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13766__CLK clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07418__S0 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06810__S net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11428__S net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09732__A1 net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08535__A2 _03481_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09732__B2 _04341_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_2503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07207__A net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13770_ clknet_leaf_60_clk _01001_ net1141 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[758\]
+ sky130_fd_sc_hd__dfrtp_1
X_10982_ net53 _05708_ vssd1 vssd1 vccd1 vccd1 _05709_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_35_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07641__S net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12721_ final_design.VGA_data_control.v_count\[2\] _06359_ vssd1 vssd1 vccd1 vccd1
+ _06362_ sky130_fd_sc_hd__and2b_1
XANTENNA__09422__A net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08394__S1 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12652_ _06313_ net1530 net979 vssd1 vssd1 vccd1 vccd1 _01328_ sky130_fd_sc_hd__mux2_1
XANTENNA__13146__CLK clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_34_clk_A clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1634 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11055__B1 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11603_ net805 _02359_ net803 vssd1 vssd1 vccd1 vccd1 _06158_ sky130_fd_sc_hd__or3b_2
X_12583_ net1565 net996 net982 final_design.data_from_mem\[1\] vssd1 vssd1 vccd1 vccd1
+ _01276_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09568__S net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11534_ net1604 net179 net524 vssd1 vssd1 vccd1 vccd1 _00401_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14253_ net1307 vssd1 vssd1 vccd1 vccd1 gpio_out[31] sky130_fd_sc_hd__buf_2
XFILLER_0_64_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_49_clk_A clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11465_ net216 net2396 net306 vssd1 vssd1 vccd1 vccd1 _00349_ sky130_fd_sc_hd__mux2_1
XANTENNA__13296__CLK clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11358__A1 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12555__B1 net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_917 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13204_ clknet_leaf_12_clk _00435_ net1090 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[192\]
+ sky130_fd_sc_hd__dfrtp_1
X_10416_ net1422 net1027 _05191_ net245 vssd1 vssd1 vccd1 vccd1 _00149_ sky130_fd_sc_hd__a22o_1
X_14184_ clknet_leaf_20_clk final_design.VGA_data_control.next_state\[0\] net1159
+ vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.state\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_0_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11396_ _04248_ net657 _06080_ vssd1 vssd1 vccd1 vccd1 _06081_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_81_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13135_ clknet_leaf_42_clk _00366_ net1222 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[123\]
+ sky130_fd_sc_hd__dfrtp_1
X_10347_ wb_manage.curr_state\[1\] net1 vssd1 vssd1 vccd1 vccd1 _05168_ sky130_fd_sc_hd__and2_1
XFILLER_0_0_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06720__S net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13066_ clknet_leaf_60_clk _00297_ net1141 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[54\]
+ sky130_fd_sc_hd__dfrtp_1
X_10278_ final_design.uart.BAUD_counter\[27\] final_design.uart.BAUD_counter\[28\]
+ _05133_ final_design.uart.BAUD_counter\[29\] vssd1 vssd1 vccd1 vccd1 _05137_ sky130_fd_sc_hd__a31o_1
XANTENNA__09184__C1 _02423_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12017_ _06219_ net290 net403 net2249 vssd1 vssd1 vccd1 vccd1 _00748_ sky130_fd_sc_hd__a22o_1
XANTENNA__09723__A1 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11530__A1 net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13968_ clknet_leaf_34_clk _01199_ net1238 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[956\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11294__B1 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12919_ clknet_leaf_31_clk _00157_ net1233 vssd1 vssd1 vccd1 vccd1 net141 sky130_fd_sc_hd__dfrtp_1
XANTENNA__12169__S net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13899_ clknet_leaf_53_clk _01130_ net1190 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[887\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06440_ wb_manage.BUSY_O net34 vssd1 vssd1 vccd1 vccd1 _01394_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_29_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_17_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14071__CLK clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13639__CLK clknet_leaf_62_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11597__A1 net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08110_ final_design.cpu.reg_window\[588\] final_design.cpu.reg_window\[620\] net812
+ vssd1 vssd1 vccd1 vccd1 _03061_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_25_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09090_ _03708_ _03720_ vssd1 vssd1 vccd1 vccd1 _04014_ sky130_fd_sc_hd__xor2_1
XFILLER_0_66_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08041_ _01853_ net618 vssd1 vssd1 vccd1 vccd1 _02992_ sky130_fd_sc_hd__nor2_1
XANTENNA__11349__A1 net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold902 final_design.reqhand.instruction\[13\] vssd1 vssd1 vccd1 vccd1 net2244 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12546__B1 net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold913 final_design.cpu.reg_window\[100\] vssd1 vssd1 vccd1 vccd1 net2255 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13789__CLK clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12010__A2 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold924 final_design.cpu.reg_window\[407\] vssd1 vssd1 vccd1 vccd1 net2266 sky130_fd_sc_hd__dlygate4sd3_1
Xhold935 final_design.cpu.reg_window\[943\] vssd1 vssd1 vccd1 vccd1 net2277 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkload36_A clknet_leaf_48_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold946 final_design.cpu.reg_window\[940\] vssd1 vssd1 vccd1 vccd1 net2288 sky130_fd_sc_hd__dlygate4sd3_1
Xhold957 final_design.cpu.reg_window\[224\] vssd1 vssd1 vccd1 vccd1 net2299 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold968 final_design.cpu.reg_window\[404\] vssd1 vssd1 vccd1 vccd1 net2310 sky130_fd_sc_hd__dlygate4sd3_1
X_09992_ net262 _04908_ _04910_ vssd1 vssd1 vccd1 vccd1 _04911_ sky130_fd_sc_hd__and3_1
XFILLER_0_42_1830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold979 final_design.cpu.reg_window\[413\] vssd1 vssd1 vccd1 vccd1 net2321 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_wire739_X net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08943_ _02462_ _03883_ vssd1 vssd1 vccd1 vccd1 _03884_ sky130_fd_sc_hd__xnor2_1
XANTENNA__13019__CLK clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout299_A _06159_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08874_ final_design.CPU_instr_adr\[29\] net1015 _03819_ _03822_ vssd1 vssd1 vccd1
+ vccd1 _00240_ sky130_fd_sc_hd__a22o_1
X_07825_ final_design.cpu.reg_window\[85\] final_design.cpu.reg_window\[117\] net867
+ vssd1 vssd1 vccd1 vccd1 _02776_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout466_A _03518_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11772__A _05849_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07756_ _01690_ net615 vssd1 vssd1 vccd1 vccd1 _02707_ sky130_fd_sc_hd__or2_1
XFILLER_0_75_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08557__S net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13169__CLK clknet_leaf_34_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1060 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06707_ net885 _01650_ _01656_ _01643_ _01644_ vssd1 vssd1 vccd1 vccd1 _01658_ sky130_fd_sc_hd__a32o_2
XFILLER_0_71_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07687_ _02637_ vssd1 vssd1 vccd1 vccd1 _02638_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout633_A _06157_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout254_X net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09426_ _02899_ net442 net439 _02898_ vssd1 vssd1 vccd1 vccd1 _04345_ sky130_fd_sc_hd__o22a_1
X_06638_ net753 _01588_ vssd1 vssd1 vccd1 vccd1 _01589_ sky130_fd_sc_hd__or2_1
XFILLER_0_66_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_964 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09357_ net489 _04275_ vssd1 vssd1 vccd1 vccd1 _04276_ sky130_fd_sc_hd__nor2_1
XFILLER_0_81_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout421_X net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_997 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06569_ _01516_ _01517_ _01518_ _01519_ net776 net794 vssd1 vssd1 vccd1 vccd1 _01520_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_69_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout519_X net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08989__C1 _03655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08308_ net597 _03257_ _03232_ net536 vssd1 vssd1 vccd1 vccd1 _03259_ sky130_fd_sc_hd__o211a_1
XANTENNA__08145__X _03096_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09288_ net606 _03550_ _03524_ _01535_ vssd1 vssd1 vccd1 vccd1 _04207_ sky130_fd_sc_hd__o211a_1
X_08239_ _03186_ _03187_ _03188_ _03189_ net678 net691 vssd1 vssd1 vccd1 vccd1 _03190_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__12537__B1 net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11250_ net425 net560 _05952_ net314 net1888 vssd1 vssd1 vccd1 vccd1 _00287_ sky130_fd_sc_hd__a32o_1
XFILLER_0_15_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12001__A2 net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1020 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout790_X net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10201_ _05088_ _05089_ _00039_ vssd1 vssd1 vccd1 vccd1 _00038_ sky130_fd_sc_hd__o21a_1
X_11181_ net427 net564 _05891_ net314 net1808 vssd1 vssd1 vccd1 vccd1 _00279_ sky130_fd_sc_hd__a32o_1
XANTENNA__06767__A1 net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07636__S net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10132_ final_design.vga.v_current_state\[1\] _04997_ _05036_ _01404_ vssd1 vssd1
+ vccd1 vccd1 final_design.vga.v_next_state\[1\] sky130_fd_sc_hd__a211o_1
XFILLER_0_21_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06862__S1 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10063_ _04290_ _04328_ _04389_ _04981_ vssd1 vssd1 vccd1 vccd1 _04982_ sky130_fd_sc_hd__and4_1
XANTENNA__09136__B _04053_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08064__S0 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07716__B1 net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input27_A DAT_I[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11369__A1_N _01599_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13822_ clknet_leaf_14_clk _01053_ net1100 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[810\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14094__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10079__A1 net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07371__S net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08694__C _03593_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13753_ clknet_leaf_56_clk _00984_ net1147 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[741\]
+ sky130_fd_sc_hd__dfrtp_1
X_10965_ _05692_ vssd1 vssd1 vccd1 vccd1 _05693_ sky130_fd_sc_hd__inv_2
X_12704_ _06340_ _06344_ vssd1 vssd1 vccd1 vccd1 _06345_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_14_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13684_ clknet_leaf_10_clk _00915_ net1102 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[672\]
+ sky130_fd_sc_hd__dfrtp_1
X_10896_ net1423 net1033 _05624_ _05626_ vssd1 vssd1 vccd1 vccd1 _00194_ sky130_fd_sc_hd__a22o_1
XFILLER_0_6_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12635_ final_design.VGA_data_control.ready_data\[5\] net1022 net976 final_design.data_from_mem\[5\]
+ vssd1 vssd1 vccd1 vccd1 _06305_ sky130_fd_sc_hd__a22o_1
XANTENNA__11579__A1 net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06715__S net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12566_ final_design.uart.receiving final_design.uart.working_data\[3\] vssd1 vssd1
+ vccd1 vccd1 _06288_ sky130_fd_sc_hd__and2_1
XFILLER_0_31_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11517_ net2126 net205 net521 vssd1 vssd1 vccd1 vccd1 _00386_ sky130_fd_sc_hd__mux2_1
XANTENNA__13931__CLK clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12497_ net568 _06158_ _06260_ vssd1 vssd1 vccd1 vccd1 _06284_ sky130_fd_sc_hd__or3_4
XANTENNA__12528__B1 net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14236_ net1290 vssd1 vssd1 vccd1 vccd1 gpio_out[14] sky130_fd_sc_hd__buf_2
XFILLER_0_65_1841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold209 final_design.cpu.reg_window\[724\] vssd1 vssd1 vccd1 vccd1 net1551 sky130_fd_sc_hd__dlygate4sd3_1
X_11448_ net241 net639 vssd1 vssd1 vccd1 vccd1 _06097_ sky130_fd_sc_hd__and2_1
XFILLER_0_46_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_1885 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08747__A2 _01598_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14167_ clknet_leaf_18_clk _01341_ net1108 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.data_to_VGA\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12452__S net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11379_ _04420_ net656 vssd1 vssd1 vccd1 vccd1 _06066_ sky130_fd_sc_hd__nand2_1
XFILLER_0_81_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08502__Y _03453_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07546__S net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13118_ clknet_leaf_13_clk _00349_ net1089 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[106\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11576__B net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14098_ clknet_leaf_22_clk _01295_ net1164 vssd1 vssd1 vccd1 vccd1 final_design.reqhand.instruction\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_37_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13049_ clknet_leaf_56_clk _00280_ net1146 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[37\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_33_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11503__A1 net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13311__CLK clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07610_ final_design.cpu.reg_window\[733\] final_design.cpu.reg_window\[765\] net870
+ vssd1 vssd1 vccd1 vccd1 _02561_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_1801 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08590_ _03537_ _03538_ _03539_ _03540_ net678 net698 vssd1 vssd1 vccd1 vccd1 _03541_
+ sky130_fd_sc_hd__mux4_1
Xclkbuf_3_4_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_3_4_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_53_1200 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06930__B2 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07541_ final_design.cpu.reg_window\[991\] final_design.cpu.reg_window\[1023\] net939
+ vssd1 vssd1 vccd1 vccd1 _02492_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_1845 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11806__A2 net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13461__CLK clknet_leaf_57_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_1889 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07472_ _02420_ _02421_ vssd1 vssd1 vccd1 vccd1 _02423_ sky130_fd_sc_hd__or2_4
XTAP_TAPCELL_ROW_27_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09211_ _02800_ _02834_ _02802_ vssd1 vssd1 vccd1 vccd1 _04130_ sky130_fd_sc_hd__o21ai_1
X_06423_ final_design.reqhand.instruction\[5\] vssd1 vssd1 vccd1 vccd1 _01378_ sky130_fd_sc_hd__inv_2
XANTENNA__10490__B2 net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11531__S net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09142_ net595 _03549_ _02389_ _02422_ vssd1 vssd1 vccd1 vccd1 _04061_ sky130_fd_sc_hd__o211a_1
XANTENNA__12231__A2 net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09073_ _02242_ _02436_ _03998_ vssd1 vssd1 vccd1 vccd1 _03999_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_31_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout214_A net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12519__B1 net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08024_ final_design.cpu.reg_window\[211\] final_design.cpu.reg_window\[243\] net830
+ vssd1 vssd1 vccd1 vccd1 _02975_ sky130_fd_sc_hd__mux2_1
Xhold710 final_design.cpu.reg_window\[85\] vssd1 vssd1 vccd1 vccd1 net2052 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold721 final_design.cpu.reg_window\[1016\] vssd1 vssd1 vccd1 vccd1 net2063 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold732 final_design.cpu.reg_window\[444\] vssd1 vssd1 vccd1 vccd1 net2074 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_9_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold743 final_design.cpu.reg_window\[78\] vssd1 vssd1 vccd1 vccd1 net2085 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold754 final_design.cpu.reg_window\[33\] vssd1 vssd1 vccd1 vccd1 net2096 sky130_fd_sc_hd__dlygate4sd3_1
Xhold765 final_design.cpu.reg_window\[888\] vssd1 vssd1 vccd1 vccd1 net2107 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1123_A net1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold776 final_design.cpu.reg_window\[281\] vssd1 vssd1 vccd1 vccd1 net2118 sky130_fd_sc_hd__dlygate4sd3_1
Xhold787 final_design.cpu.reg_window\[403\] vssd1 vssd1 vccd1 vccd1 net2129 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11486__B net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold798 final_design.cpu.reg_window\[952\] vssd1 vssd1 vccd1 vccd1 net2140 sky130_fd_sc_hd__dlygate4sd3_1
X_09975_ _04221_ _04533_ _04539_ _04728_ _04893_ vssd1 vssd1 vccd1 vccd1 _04894_ sky130_fd_sc_hd__a221o_1
XANTENNA__06844__S1 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout583_A net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08926_ _03797_ _03868_ vssd1 vssd1 vccd1 vccd1 _03869_ sky130_fd_sc_hd__or2_1
XANTENNA__09699__A0 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08857_ _03658_ _03778_ vssd1 vssd1 vccd1 vccd1 _03807_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout371_X net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout750_A net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06867__Y _01818_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout469_X net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07808_ final_design.cpu.reg_window\[601\] final_design.cpu.reg_window\[633\] net850
+ vssd1 vssd1 vccd1 vccd1 _02759_ sky130_fd_sc_hd__mux2_1
X_08788_ _03679_ _03680_ vssd1 vssd1 vccd1 vccd1 _03739_ sky130_fd_sc_hd__nor2_1
XANTENNA__13804__CLK clknet_leaf_46_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06596__A net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11258__B1 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07739_ final_design.cpu.reg_window\[922\] final_design.cpu.reg_window\[954\] net863
+ vssd1 vssd1 vccd1 vccd1 _02690_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout636_X net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10750_ _05485_ _05486_ _05466_ vssd1 vssd1 vccd1 vccd1 _05487_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_3_1705 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12470__A2 net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1885 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09409_ _04325_ _04326_ vssd1 vssd1 vccd1 vccd1 _04328_ sky130_fd_sc_hd__nand2_1
XFILLER_0_36_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13954__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10681_ _05402_ _05404_ _05400_ vssd1 vssd1 vccd1 vccd1 _05422_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_36_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07882__C1 net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1749 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11441__S net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12758__B1 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12420_ net194 net553 net501 net339 net1724 vssd1 vssd1 vccd1 vccd1 _01129_ sky130_fd_sc_hd__a32o_1
XFILLER_0_8_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10565__B final_design.VGA_adr\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12351_ _06235_ _06264_ net362 net2517 vssd1 vssd1 vccd1 vccd1 _01063_ sky130_fd_sc_hd__a22o_1
XANTENNA__06988__A1 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06988__B2 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11302_ final_design.data_from_mem\[19\] net235 net233 vssd1 vssd1 vccd1 vccd1 _05998_
+ sky130_fd_sc_hd__a21o_1
X_12282_ net572 _06212_ net508 net371 net1747 vssd1 vssd1 vccd1 vccd1 _00997_ sky130_fd_sc_hd__a32o_1
X_14021_ clknet_leaf_49_clk _01252_ net1182 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[1009\]
+ sky130_fd_sc_hd__dfrtp_1
X_11233_ net662 _03962_ net736 vssd1 vssd1 vccd1 vccd1 _05937_ sky130_fd_sc_hd__a21o_1
XFILLER_0_43_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11164_ net2486 net315 _05876_ net430 vssd1 vssd1 vccd1 vccd1 _00277_ sky130_fd_sc_hd__a22o_1
XANTENNA__13334__CLK clknet_leaf_59_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10115_ final_design.VGA_data_control.v_count\[5\] net1051 _05023_ vssd1 vssd1 vccd1
+ vccd1 _05026_ sky130_fd_sc_hd__and3_1
XFILLER_0_25_1891 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11095_ _05798_ _05815_ net1003 vssd1 vssd1 vccd1 vccd1 _05817_ sky130_fd_sc_hd__o21a_1
X_10046_ net730 _04576_ _04597_ _04421_ _04423_ vssd1 vssd1 vccd1 vccd1 _04965_ sky130_fd_sc_hd__a32o_1
Xhold70 final_design.reqhand.data_from_UART\[0\] vssd1 vssd1 vccd1 vccd1 net1412 sky130_fd_sc_hd__dlygate4sd3_1
Xhold81 net114 vssd1 vssd1 vccd1 vccd1 net1423 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13484__CLK clknet_leaf_46_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold92 final_design.cpu.reg_window\[710\] vssd1 vssd1 vccd1 vccd1 net1434 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09153__Y _04072_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08197__S net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13805_ clknet_leaf_53_clk _01036_ net1190 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[793\]
+ sky130_fd_sc_hd__dfrtp_1
X_11997_ _06199_ net283 net401 net2125 vssd1 vssd1 vccd1 vccd1 _00728_ sky130_fd_sc_hd__a22o_1
X_10948_ _05634_ _05653_ _05675_ vssd1 vssd1 vccd1 vccd1 _05676_ sky130_fd_sc_hd__a21o_1
X_13736_ clknet_leaf_40_clk _00967_ net1220 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[724\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_50_1439 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10472__A1 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09610__A net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10879_ net81 net1046 vssd1 vssd1 vccd1 vccd1 _05610_ sky130_fd_sc_hd__nor2_1
X_13667_ clknet_leaf_0_clk _00898_ net1061 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[655\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12447__S net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12618_ net1806 final_design.reqhand.data_from_UART\[4\] _05080_ vssd1 vssd1 vccd1
+ vccd1 _01311_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13598_ clknet_leaf_12_clk _00829_ net1086 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[586\]
+ sky130_fd_sc_hd__dfrtp_1
X_12549_ _06212_ net351 net325 net2181 vssd1 vssd1 vccd1 vccd1 _01253_ sky130_fd_sc_hd__a22o_1
XFILLER_0_13_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_1 _01752_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14219_ net1277 vssd1 vssd1 vccd1 vccd1 gpio_oeb[31] sky130_fd_sc_hd__buf_2
XANTENNA__12182__S net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout508 net515 vssd1 vssd1 vccd1 vccd1 net508 sky130_fd_sc_hd__clkbuf_4
Xfanout519 net520 vssd1 vssd1 vccd1 vccd1 net519 sky130_fd_sc_hd__buf_4
X_09760_ _04659_ _04677_ vssd1 vssd1 vccd1 vccd1 _04679_ sky130_fd_sc_hd__nand2_1
X_06972_ net763 _01922_ vssd1 vssd1 vccd1 vccd1 _01923_ sky130_fd_sc_hd__or2_1
XANTENNA__13827__CLK clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08628__A_N _02026_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08711_ final_design.CPU_instr_adr\[26\] _01630_ vssd1 vssd1 vccd1 vccd1 _03662_
+ sky130_fd_sc_hd__nand2_1
X_09691_ _04340_ _04608_ _04609_ _04604_ _04605_ vssd1 vssd1 vccd1 vccd1 _04610_ sky130_fd_sc_hd__a311o_1
XFILLER_0_59_1431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11526__S net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1090 net1117 vssd1 vssd1 vccd1 vccd1 net1090 sky130_fd_sc_hd__clkbuf_4
X_08642_ _02838_ _02901_ _03030_ _03591_ vssd1 vssd1 vccd1 vccd1 _03593_ sky130_fd_sc_hd__and4_1
XPHY_EDGE_ROW_16_Left_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_1_237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12851__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13977__CLK clknet_leaf_56_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08573_ _02424_ net596 vssd1 vssd1 vccd1 vccd1 _03524_ sky130_fd_sc_hd__nand2_4
XFILLER_0_77_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07524_ _01567_ _01570_ _02474_ vssd1 vssd1 vccd1 vccd1 _02475_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_77_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08656__A1 _01535_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09853__B1 net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10463__B2 net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11660__B1 net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07455_ net758 _02405_ vssd1 vssd1 vccd1 vccd1 _02406_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout331_A _06283_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13207__CLK clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout429_A net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06406_ final_design.CPU_instr_adr\[24\] vssd1 vssd1 vccd1 vccd1 _01361_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07386_ _02333_ _02334_ _02335_ _02336_ net770 net789 vssd1 vssd1 vccd1 vccd1 _02337_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__12204__A2 net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09125_ net958 net955 net961 vssd1 vssd1 vccd1 vccd1 _04044_ sky130_fd_sc_hd__a21o_1
XFILLER_0_66_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout217_X net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1240_A net1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_1446 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09056_ _02439_ _02440_ vssd1 vssd1 vccd1 vccd1 _03984_ sky130_fd_sc_hd__and2_1
XANTENNA__13357__CLK clknet_leaf_44_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08007_ final_design.cpu.reg_window\[528\] final_design.cpu.reg_window\[560\] net843
+ vssd1 vssd1 vccd1 vccd1 _02958_ sky130_fd_sc_hd__mux2_1
Xhold540 final_design.cpu.reg_window\[833\] vssd1 vssd1 vccd1 vccd1 net1882 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09238__Y _04157_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold551 final_design.cpu.reg_window\[519\] vssd1 vssd1 vccd1 vccd1 net1893 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10518__A2 net1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold562 final_design.cpu.reg_window\[250\] vssd1 vssd1 vccd1 vccd1 net1904 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_3_3_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold573 final_design.cpu.reg_window\[601\] vssd1 vssd1 vccd1 vccd1 net1915 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09384__A2 _02091_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold584 final_design.cpu.reg_window\[655\] vssd1 vssd1 vccd1 vccd1 net1926 sky130_fd_sc_hd__dlygate4sd3_1
Xhold595 final_design.cpu.reg_window\[568\] vssd1 vssd1 vccd1 vccd1 net1937 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout965_A net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout586_X net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_1829 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_2587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09958_ _03488_ _04145_ vssd1 vssd1 vccd1 vccd1 _04877_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_70_2598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11479__A0 net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08909_ _03853_ vssd1 vssd1 vccd1 vccd1 _03854_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout753_X net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09889_ net90 net93 vssd1 vssd1 vccd1 vccd1 _04808_ sky130_fd_sc_hd__xor2_1
XANTENNA__11436__S net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09687__A3 net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11920_ net177 net2221 net275 vssd1 vssd1 vccd1 vccd1 _00658_ sky130_fd_sc_hd__mux2_1
XANTENNA__12691__A2 _05039_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11851_ _06101_ net281 net518 net2292 vssd1 vssd1 vccd1 vccd1 _00601_ sky130_fd_sc_hd__a22o_1
X_10802_ net959 _05534_ _05536_ net956 vssd1 vssd1 vccd1 vccd1 _05537_ sky130_fd_sc_hd__o22a_1
XFILLER_0_79_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11782_ net2322 net412 net277 _05929_ vssd1 vssd1 vccd1 vccd1 _00540_ sky130_fd_sc_hd__a22o_1
XFILLER_0_36_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10733_ _05469_ _05470_ vssd1 vssd1 vccd1 vccd1 _05471_ sky130_fd_sc_hd__or2_1
X_13521_ clknet_leaf_35_clk _00752_ net1240 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[509\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14132__CLK clknet_leaf_17_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1546 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13452_ clknet_leaf_45_clk _00683_ net1215 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[440\]
+ sky130_fd_sc_hd__dfrtp_1
X_10664_ net1449 net1031 net1003 _05405_ vssd1 vssd1 vccd1 vccd1 _00183_ sky130_fd_sc_hd__a22o_1
XANTENNA_input94_A memory_size[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12403_ _06101_ net347 net338 net2414 vssd1 vssd1 vccd1 vccd1 _01113_ sky130_fd_sc_hd__a22o_1
XFILLER_0_63_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13383_ clknet_leaf_58_clk _00614_ net1125 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[371\]
+ sky130_fd_sc_hd__dfrtp_1
X_10595_ net958 _05338_ _05339_ net955 vssd1 vssd1 vccd1 vccd1 _05340_ sky130_fd_sc_hd__o22a_1
XFILLER_0_10_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_11_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12334_ _06230_ net500 net360 net2311 vssd1 vssd1 vccd1 vccd1 _01046_ sky130_fd_sc_hd__a22o_1
XANTENNA__09429__X _04348_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07622__A2 _02570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12265_ net566 _06195_ net506 net369 net1682 vssd1 vssd1 vccd1 vccd1 _00980_ sky130_fd_sc_hd__a32o_1
XFILLER_0_62_1833 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11706__A1 net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14004_ clknet_leaf_8_clk _01235_ net1154 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[992\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14091__RESET_B net1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11216_ net2403 net314 _05922_ net425 vssd1 vssd1 vccd1 vccd1 _00283_ sky130_fd_sc_hd__a22o_1
XFILLER_0_62_1877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12196_ net671 _06124_ _06262_ vssd1 vssd1 vccd1 vccd1 _06271_ sky130_fd_sc_hd__or3_4
XFILLER_0_43_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11147_ final_design.reqhand.data_from_UART\[1\] final_design.data_from_mem\[1\]
+ net245 vssd1 vssd1 vccd1 vccd1 _05861_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12874__CLK clknet_leaf_15_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11078_ _05763_ _05779_ _05782_ vssd1 vssd1 vccd1 vccd1 _05800_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_21_1585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10029_ net494 _04836_ _04838_ _04231_ vssd1 vssd1 vccd1 vccd1 _04948_ sky130_fd_sc_hd__a31o_1
XFILLER_0_76_1063 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11890__A0 net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09611__Y _04530_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10445__B2 net245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11642__B1 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13719_ clknet_leaf_6_clk _00950_ net1130 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[707\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12177__S net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07240_ final_design.cpu.reg_window\[7\] final_design.cpu.reg_window\[39\] net887
+ vssd1 vssd1 vccd1 vccd1 _02191_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12198__A1 net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07171_ final_design.cpu.reg_window\[586\] final_design.cpu.reg_window\[618\] net895
+ vssd1 vssd1 vccd1 vccd1 _02122_ sky130_fd_sc_hd__mux2_1
XANTENNA__08497__S0 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12955__RESET_B net1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11110__A net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1917 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout305 _06125_ vssd1 vssd1 vccd1 vccd1 net305 sky130_fd_sc_hd__buf_4
XFILLER_0_1_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11173__A2 net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout316 net317 vssd1 vssd1 vccd1 vccd1 net316 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_22_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09812_ net489 _04368_ _04727_ _04730_ net263 vssd1 vssd1 vccd1 vccd1 _04731_ sky130_fd_sc_hd__o311a_1
Xfanout327 _06284_ vssd1 vssd1 vccd1 vccd1 net327 sky130_fd_sc_hd__buf_4
Xfanout338 net339 vssd1 vssd1 vccd1 vccd1 net338 sky130_fd_sc_hd__buf_4
XANTENNA__10381__B1 net1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout349 net350 vssd1 vssd1 vccd1 vccd1 net349 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10920__A2 net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14005__CLK clknet_leaf_57_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06955_ _01902_ _01903_ _01904_ _01905_ net772 net784 vssd1 vssd1 vccd1 vccd1 _01906_
+ sky130_fd_sc_hd__mux4_1
X_09743_ net318 _04278_ vssd1 vssd1 vccd1 vccd1 _04662_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout281_A net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout379_A _06271_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09674_ _02838_ _04352_ net321 _03035_ vssd1 vssd1 vccd1 vccd1 _04593_ sky130_fd_sc_hd__a211o_1
X_06886_ net759 _01836_ vssd1 vssd1 vccd1 vccd1 _01837_ sky130_fd_sc_hd__nor2_1
X_08625_ _03262_ _03574_ _03573_ vssd1 vssd1 vccd1 vccd1 _03576_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_39_1879 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11881__B1 net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1190_A net1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14155__CLK clknet_leaf_18_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11780__A net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout546_A _01880_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08556_ final_design.cpu.reg_window\[705\] final_design.cpu.reg_window\[737\] net833
+ vssd1 vssd1 vccd1 vccd1 _03507_ sky130_fd_sc_hd__mux2_1
XANTENNA__08629__A1 net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12425__A2 net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09888__C _04805_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06874__A net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07507_ _01884_ _02457_ vssd1 vssd1 vccd1 vccd1 _02458_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_82_2992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_1833 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08487_ net709 _03431_ net722 vssd1 vssd1 vccd1 vccd1 _03438_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout334_X net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout713_A net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07438_ net883 _02382_ _02388_ _02375_ _02376_ vssd1 vssd1 vccd1 vccd1 _02389_ sky130_fd_sc_hd__a32oi_4
XANTENNA__12189__A1 net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwire739 _01490_ vssd1 vssd1 vccd1 vccd1 net739 sky130_fd_sc_hd__buf_2
XANTENNA_fanout501_X net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07369_ final_design.cpu.reg_window\[643\] final_design.cpu.reg_window\[675\] net908
+ vssd1 vssd1 vccd1 vccd1 _02320_ sky130_fd_sc_hd__mux2_1
XANTENNA__09054__B2 net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09108_ _02426_ _02427_ net619 vssd1 vssd1 vccd1 vccd1 _04029_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_60_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10380_ net23 net1023 net1007 final_design.data_from_mem\[29\] vssd1 vssd1 vccd1
+ vccd1 _00133_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_57_2140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_2151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_2785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_57_2162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09039_ _02159_ _02443_ _02130_ vssd1 vssd1 vccd1 vccd1 _03969_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_53_2004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_2796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_2015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_2026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12050_ net1700 net192 net399 vssd1 vssd1 vccd1 vccd1 _00778_ sky130_fd_sc_hd__mux2_1
XANTENNA__12897__CLK clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold370 final_design.cpu.reg_window\[94\] vssd1 vssd1 vccd1 vccd1 net1712 sky130_fd_sc_hd__dlygate4sd3_1
Xhold381 final_design.cpu.reg_window\[553\] vssd1 vssd1 vccd1 vccd1 net1723 sky130_fd_sc_hd__dlygate4sd3_1
X_11001_ net1055 _05724_ _05239_ final_design.CPU_instr_adr\[26\] vssd1 vssd1 vccd1
+ vccd1 _05727_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__11164__A2 net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold392 final_design.cpu.reg_window\[67\] vssd1 vssd1 vccd1 vccd1 net1734 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10372__B1 net1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout850 net851 vssd1 vssd1 vccd1 vccd1 net850 sky130_fd_sc_hd__clkbuf_4
Xfanout861 net862 vssd1 vssd1 vccd1 vccd1 net861 sky130_fd_sc_hd__clkbuf_4
Xfanout872 net873 vssd1 vssd1 vccd1 vccd1 net872 sky130_fd_sc_hd__clkbuf_4
Xfanout883 _01437_ vssd1 vssd1 vccd1 vccd1 net883 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_5_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout894 net896 vssd1 vssd1 vccd1 vccd1 net894 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_5_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12952_ clknet_leaf_29_clk _00190_ net1195 vssd1 vssd1 vccd1 vccd1 net109 sky130_fd_sc_hd__dfrtp_1
Xhold1070 final_design.cpu.reg_window\[298\] vssd1 vssd1 vccd1 vccd1 net2412 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_73_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1081 final_design.uart.working_data\[7\] vssd1 vssd1 vccd1 vccd1 net2423 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10675__A1 net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11903_ net201 net1962 net273 vssd1 vssd1 vccd1 vccd1 _00645_ sky130_fd_sc_hd__mux2_1
Xhold1092 final_design.cpu.reg_window\[357\] vssd1 vssd1 vccd1 vccd1 net2434 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10675__B2 net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12883_ clknet_leaf_18_clk _00121_ net1111 vssd1 vssd1 vccd1 vccd1 final_design.data_from_mem\[17\]
+ sky130_fd_sc_hd__dfrtp_4
X_11834_ net193 net2069 net266 vssd1 vssd1 vccd1 vccd1 _00586_ sky130_fd_sc_hd__mux2_1
XANTENNA__12416__A2 net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09817__B1 net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13522__CLK clknet_leaf_39_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11624__B1 net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11765_ net181 net2345 net418 vssd1 vssd1 vccd1 vccd1 _00528_ sky130_fd_sc_hd__mux2_1
X_10716_ net802 _05452_ _05454_ _04036_ vssd1 vssd1 vccd1 vccd1 _05455_ sky130_fd_sc_hd__o22a_1
X_13504_ clknet_leaf_11_clk _00735_ net1097 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[492\]
+ sky130_fd_sc_hd__dfrtp_1
X_11696_ net426 net560 _06206_ net294 net1940 vssd1 vssd1 vccd1 vccd1 _00479_ sky130_fd_sc_hd__a32o_1
X_10647_ _05354_ _05374_ _05373_ _05371_ vssd1 vssd1 vccd1 vccd1 _05389_ sky130_fd_sc_hd__o211a_1
X_13435_ clknet_leaf_0_clk _00666_ net1071 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[423\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13672__CLK clknet_leaf_40_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11927__B2 net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13366_ clknet_leaf_58_clk _00597_ net1125 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[354\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09596__A2 _04240_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10578_ net668 _05310_ _05323_ vssd1 vssd1 vccd1 vccd1 _05324_ sky130_fd_sc_hd__o21a_1
XFILLER_0_24_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08504__A _02325_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_929 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12317_ net2262 net197 net366 vssd1 vssd1 vccd1 vccd1 _01031_ sky130_fd_sc_hd__mux2_1
X_13297_ clknet_leaf_35_clk _00528_ net1241 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[285\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_1761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09348__A2 net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12248_ net574 _06177_ net509 net375 net1569 vssd1 vssd1 vccd1 vccd1 _00964_ sky130_fd_sc_hd__a32o_1
XANTENNA__14028__CLK clknet_leaf_46_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12460__S net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12179_ net1926 net205 net380 vssd1 vssd1 vccd1 vccd1 _00898_ sky130_fd_sc_hd__mux2_1
XANTENNA__10363__B1 net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07454__S1 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11584__B net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14178__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13052__CLK clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06740_ _01499_ net665 _01689_ vssd1 vssd1 vccd1 vccd1 _01691_ sky130_fd_sc_hd__or3b_2
XFILLER_0_3_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09520__A2 _04435_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06671_ final_design.cpu.reg_window\[730\] final_design.cpu.reg_window\[762\] net941
+ vssd1 vssd1 vccd1 vccd1 _01622_ sky130_fd_sc_hd__mux2_1
X_08410_ final_design.cpu.reg_window\[325\] final_design.cpu.reg_window\[357\] net842
+ vssd1 vssd1 vccd1 vccd1 _03361_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09390_ _04307_ _04308_ net475 vssd1 vssd1 vccd1 vccd1 _04309_ sky130_fd_sc_hd__mux2_2
XANTENNA__12407__A2 net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08341_ net598 _03287_ _03263_ _02184_ vssd1 vssd1 vccd1 vccd1 _03292_ sky130_fd_sc_hd__o211a_1
XANTENNA__10418__B2 net246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10969__A2 net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_1817 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08272_ _03217_ _03222_ net708 vssd1 vssd1 vccd1 vccd1 _03223_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07223_ final_design.cpu.reg_window\[584\] final_design.cpu.reg_window\[616\] net888
+ vssd1 vssd1 vccd1 vccd1 _02174_ sky130_fd_sc_hd__mux2_1
XANTENNA__07729__S net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07154_ final_design.cpu.reg_window\[266\] final_design.cpu.reg_window\[298\] net898
+ vssd1 vssd1 vccd1 vccd1 _02105_ sky130_fd_sc_hd__mux2_1
XANTENNA__08244__C1 net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11394__A2 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12591__B2 final_design.data_from_mem\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07085_ final_design.cpu.reg_window\[460\] final_design.cpu.reg_window\[492\] net898
+ vssd1 vssd1 vccd1 vccd1 _02036_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_1861 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11146__A2 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout496_A net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12343__B2 _05952_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12370__S net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10354__B1 net1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1203_A net1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07464__S net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input1_A ACK_I vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11494__B net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07987_ final_design.cpu.reg_window\[336\] final_design.cpu.reg_window\[368\] net847
+ vssd1 vssd1 vccd1 vccd1 _02938_ sky130_fd_sc_hd__mux2_1
Xfanout179 _06081_ vssd1 vssd1 vccd1 vccd1 net179 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout284_X net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06938_ _01885_ _01886_ _01887_ _01888_ net772 net784 vssd1 vssd1 vccd1 vccd1 _01889_
+ sky130_fd_sc_hd__mux4_1
X_09726_ _01596_ _01626_ _01657_ net552 net453 net463 vssd1 vssd1 vccd1 vccd1 _04645_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_9_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10657__A1 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13545__CLK clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_2420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09657_ _04190_ _04575_ vssd1 vssd1 vccd1 vccd1 _04576_ sky130_fd_sc_hd__and2_1
XANTENNA__10657__B2 net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06869_ _01464_ _01468_ _01475_ _01483_ vssd1 vssd1 vccd1 vccd1 _01820_ sky130_fd_sc_hd__or4_2
XANTENNA__11854__B1 net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout830_A net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_2431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_2442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout928_A net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout549_X net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08608_ net528 net475 vssd1 vssd1 vccd1 vccd1 _03559_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_80_2929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09588_ _03134_ _04506_ net450 vssd1 vssd1 vccd1 vccd1 _04507_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_61_2306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10409__B2 net246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08539_ final_design.cpu.reg_window\[257\] final_design.cpu.reg_window\[289\] net838
+ vssd1 vssd1 vccd1 vccd1 _03490_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout716_X net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13695__CLK clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11550_ net237 net635 vssd1 vssd1 vccd1 vccd1 _06131_ sky130_fd_sc_hd__and2_1
XFILLER_0_65_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10501_ net725 _04825_ net250 _04990_ vssd1 vssd1 vccd1 vccd1 _05250_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_11_1551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11481_ net194 net2302 net307 vssd1 vssd1 vccd1 vccd1 _00361_ sky130_fd_sc_hd__mux2_1
Xwire525 _03549_ vssd1 vssd1 vccd1 vccd1 net525 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_59_2213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire536 _02155_ vssd1 vssd1 vccd1 vccd1 net536 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_59_2224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_78_2858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13220_ clknet_leaf_54_clk _00451_ net1179 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[208\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_59_2235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_2869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10432_ net592 _02961_ vssd1 vssd1 vccd1 vccd1 _05200_ sky130_fd_sc_hd__and2b_1
X_14190__1249 vssd1 vssd1 vccd1 vccd1 _14190__1249/HI net1249 sky130_fd_sc_hd__conb_1
XANTENNA__07589__A1 net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07133__S0 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13151_ clknet_leaf_8_clk _00382_ net1154 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[139\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_61_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10363_ net5 net1024 net1006 final_design.data_from_mem\[12\] vssd1 vssd1 vccd1 vccd1
+ _00116_ sky130_fd_sc_hd__o22a_1
XFILLER_0_66_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12102_ net1640 net243 net388 vssd1 vssd1 vccd1 vccd1 _00826_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_1901 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13082_ clknet_leaf_6_clk _00313_ net1128 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[70\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input57_A mem_adr_start[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10294_ final_design.VGA_data_control.data_to_VGA\[7\] final_design.VGA_data_control.data_to_VGA\[6\]
+ net1050 vssd1 vssd1 vccd1 vccd1 _05148_ sky130_fd_sc_hd__mux2_1
XFILLER_0_40_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12033_ net1571 net237 net397 vssd1 vssd1 vccd1 vccd1 _00761_ sky130_fd_sc_hd__mux2_1
XANTENNA__13075__CLK clknet_leaf_40_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10345__B1 net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07436__S1 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09750__A2 net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_8_clk_A clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout680 net681 vssd1 vssd1 vccd1 vccd1 net680 sky130_fd_sc_hd__buf_4
Xfanout691 net692 vssd1 vssd1 vccd1 vccd1 net691 sky130_fd_sc_hd__clkbuf_8
X_13984_ clknet_leaf_11_clk _01215_ net1097 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[972\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11845__A0 net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12935_ clknet_leaf_22_clk _00173_ net1165 vssd1 vssd1 vccd1 vccd1 net101 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12912__CLK clknet_leaf_61_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06718__S net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12866_ clknet_leaf_25_clk _00104_ net1156 vssd1 vssd1 vccd1 vccd1 final_design.data_from_mem\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_69_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1331 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11817_ net238 net2209 net265 vssd1 vssd1 vccd1 vccd1 _00569_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12270__B1 net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07816__A2 _02763_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11748_ net213 net2246 net416 vssd1 vssd1 vccd1 vccd1 _00511_ sky130_fd_sc_hd__mux2_1
XANTENNA__07372__S0 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_12_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12455__S net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11679_ net239 net626 vssd1 vssd1 vccd1 vccd1 _06198_ sky130_fd_sc_hd__and2_1
X_13418_ clknet_leaf_59_clk _00649_ net1143 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[406\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12022__B1 net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13349_ clknet_leaf_52_clk _00580_ net1182 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[337\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13418__CLK clknet_leaf_59_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07910_ _02857_ _02858_ _02859_ _02860_ net683 net693 vssd1 vssd1 vccd1 vccd1 _02861_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__12190__S net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08890_ final_design.CPU_instr_adr\[27\] _03799_ vssd1 vssd1 vccd1 vccd1 _03837_
+ sky130_fd_sc_hd__xnor2_1
XANTENNA__13568__CLK clknet_leaf_11_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07841_ final_design.cpu.reg_window\[661\] final_design.cpu.reg_window\[693\] net858
+ vssd1 vssd1 vccd1 vccd1 _02792_ sky130_fd_sc_hd__mux2_1
X_07772_ final_design.cpu.reg_window\[920\] final_design.cpu.reg_window\[952\] net864
+ vssd1 vssd1 vccd1 vccd1 _02723_ sky130_fd_sc_hd__mux2_1
XANTENNA__12089__B1 net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10004__A _04918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10639__A1 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12797__28_A clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06723_ net753 _01673_ net748 vssd1 vssd1 vccd1 vccd1 _01674_ sky130_fd_sc_hd__o21a_1
X_09511_ _02965_ _04351_ _03028_ vssd1 vssd1 vccd1 vccd1 _04430_ sky130_fd_sc_hd__a21oi_1
XANTENNA__06938__S0 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11534__S net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09442_ _02769_ _03597_ _04046_ vssd1 vssd1 vccd1 vccd1 _04361_ sky130_fd_sc_hd__o21a_1
X_06654_ final_design.cpu.reg_window\[410\] final_design.cpu.reg_window\[442\] net944
+ vssd1 vssd1 vccd1 vccd1 _01605_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06628__S net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09373_ _03606_ _04046_ vssd1 vssd1 vccd1 vccd1 _04292_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06585_ net884 _01528_ _01534_ _01521_ _01522_ vssd1 vssd1 vccd1 vccd1 _01536_ sky130_fd_sc_hd__a32o_2
XANTENNA_fanout244_A _05910_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11064__A1 net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08324_ net707 _03268_ net722 vssd1 vssd1 vccd1 vccd1 _03275_ sky130_fd_sc_hd__o21a_1
XFILLER_0_34_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12261__B1 net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08255_ net708 _03205_ vssd1 vssd1 vccd1 vccd1 _03206_ sky130_fd_sc_hd__nor2_1
XANTENNA__09009__A1 net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12365__S net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout509_A net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1153_A net1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07459__S net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07206_ net666 _01537_ vssd1 vssd1 vccd1 vccd1 _02157_ sky130_fd_sc_hd__nand2_1
XANTENNA__12013__B1 net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08186_ final_design.cpu.reg_window\[270\] final_design.cpu.reg_window\[302\] net825
+ vssd1 vssd1 vccd1 vccd1 _03137_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_73_2700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_73_2711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13098__CLK clknet_leaf_61_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07137_ final_design.cpu.reg_window\[523\] final_design.cpu.reg_window\[555\] net908
+ vssd1 vssd1 vccd1 vccd1 _02088_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1246 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07068_ _02015_ _02016_ _02017_ _02018_ net774 net792 vssd1 vssd1 vccd1 vccd1 _02019_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__07440__B1 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout780_A net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout878_A net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout499_X net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10613__S net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07418__S1 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12935__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_2504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07922__S net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09709_ _03068_ _04627_ _03101_ vssd1 vssd1 vccd1 vccd1 _04628_ sky130_fd_sc_hd__a21oi_1
X_10981_ net802 _05704_ _05707_ _05696_ vssd1 vssd1 vccd1 vccd1 _05708_ sky130_fd_sc_hd__o211a_1
XFILLER_0_69_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12720_ _06355_ _06356_ _06360_ vssd1 vssd1 vccd1 vccd1 _06361_ sky130_fd_sc_hd__a21o_1
XFILLER_0_74_1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12651_ final_design.VGA_data_control.ready_data\[13\] net1020 net975 final_design.data_from_mem\[13\]
+ vssd1 vssd1 vccd1 vccd1 _06313_ sky130_fd_sc_hd__a22o_1
XANTENNA__09248__A1 _04158_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_4_Left_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11602_ _02095_ _02358_ net803 vssd1 vssd1 vccd1 vccd1 _06157_ sky130_fd_sc_hd__and3b_2
XFILLER_0_13_1646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12252__B1 net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12582_ net1510 net997 net983 final_design.data_from_mem\[0\] vssd1 vssd1 vccd1 vccd1
+ _01275_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07354__S0 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10802__A1 net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10802__B2 net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11533_ net2230 net180 net523 vssd1 vssd1 vccd1 vccd1 _00400_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_22_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08471__A2 _03415_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14252_ net1306 vssd1 vssd1 vccd1 vccd1 gpio_out[30] sky130_fd_sc_hd__buf_2
XFILLER_0_29_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12004__B1 net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11464_ net217 net638 vssd1 vssd1 vccd1 vccd1 _06105_ sky130_fd_sc_hd__and2_1
X_10415_ _03287_ _05190_ vssd1 vssd1 vccd1 vccd1 _05191_ sky130_fd_sc_hd__nor2_1
X_13203_ clknet_leaf_40_clk _00434_ net1206 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[191\]
+ sky130_fd_sc_hd__dfrtp_1
X_14183_ clknet_leaf_29_clk _01357_ net1194 vssd1 vssd1 vccd1 vccd1 final_design.VGA_adr\[10\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_1_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11395_ net657 _06077_ _06079_ net590 vssd1 vssd1 vccd1 vccd1 _06080_ sky130_fd_sc_hd__o31a_1
XFILLER_0_60_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10346_ net1468 net1012 net989 final_design.data_from_mem\[31\] vssd1 vssd1 vccd1
+ vccd1 _00103_ sky130_fd_sc_hd__a22o_1
X_13134_ clknet_leaf_45_clk _00365_ net1213 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[122\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_46_1488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12307__A1 net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13710__CLK clknet_leaf_43_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07982__A1 net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13065_ clknet_leaf_36_clk _00296_ net1229 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[53\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10318__B1 net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10277_ net1911 _05134_ _05136_ vssd1 vssd1 vccd1 vccd1 _00026_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_29_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12016_ _06218_ net291 net402 net2058 vssd1 vssd1 vccd1 vccd1 _00747_ sky130_fd_sc_hd__a22o_1
XANTENNA__09184__B1 _01536_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09723__A2 net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1827 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_1849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13860__CLK clknet_leaf_52_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11818__A0 net244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13967_ clknet_leaf_42_clk _01198_ net1222 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[955\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12086__A3 net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11294__A1 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12918_ clknet_leaf_62_clk _00156_ net1123 vssd1 vssd1 vccd1 vccd1 net140 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12491__B1 net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13898_ clknet_leaf_59_clk _01129_ net1142 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[886\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_75_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12849_ clknet_leaf_17_clk _00087_ net1113 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.ready_data\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_8_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11046__A1 net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11046__B2 net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12243__B1 net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06972__A net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_1779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10494__A net58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13240__CLK clknet_leaf_62_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08040_ net875 _02972_ _02978_ _02984_ _02990_ vssd1 vssd1 vccd1 vccd1 _02991_ sky130_fd_sc_hd__o32a_4
XFILLER_0_9_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11349__A2 net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold903 final_design.cpu.reg_window\[156\] vssd1 vssd1 vccd1 vccd1 net2245 sky130_fd_sc_hd__dlygate4sd3_1
Xhold914 final_design.cpu.reg_window\[875\] vssd1 vssd1 vccd1 vccd1 net2256 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09411__A1 _04158_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold925 final_design.reqhand.data_from_UART\[2\] vssd1 vssd1 vccd1 vccd1 net2267
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold936 final_design.cpu.reg_window\[813\] vssd1 vssd1 vccd1 vccd1 net2278 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_53_clk_X clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold947 final_design.cpu.reg_window\[323\] vssd1 vssd1 vccd1 vccd1 net2289 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13390__CLK clknet_leaf_42_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold958 final_design.cpu.reg_window\[680\] vssd1 vssd1 vccd1 vccd1 net2300 sky130_fd_sc_hd__dlygate4sd3_1
Xhold969 final_design.cpu.reg_window\[803\] vssd1 vssd1 vccd1 vccd1 net2311 sky130_fd_sc_hd__dlygate4sd3_1
X_09991_ _02738_ net445 net439 _02735_ _04909_ vssd1 vssd1 vccd1 vccd1 _04910_ sky130_fd_sc_hd__o221a_1
XANTENNA_clkload29_A clknet_leaf_51_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11529__S net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12958__CLK clknet_leaf_30_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08942_ _01789_ _01790_ vssd1 vssd1 vccd1 vccd1 _03883_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_77_1905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08873_ net257 _03821_ net1015 vssd1 vssd1 vccd1 vccd1 _03822_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout194_A net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07824_ final_design.cpu.reg_window\[149\] final_design.cpu.reg_window\[181\] net857
+ vssd1 vssd1 vccd1 vccd1 _02775_ sky130_fd_sc_hd__mux2_1
XANTENNA__11772__B net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11809__B1 net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07755_ _02670_ _02671_ _02701_ _02703_ vssd1 vssd1 vccd1 vccd1 _02706_ sky130_fd_sc_hd__o22a_1
XANTENNA__12077__A3 net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout361_A net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout459_A _03551_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06706_ net885 _01650_ _01656_ _01643_ _01644_ vssd1 vssd1 vccd1 vccd1 _01657_ sky130_fd_sc_hd__a32oi_4
XANTENNA__11285__A1 final_design.data_from_mem\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12482__B1 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07686_ net614 _02635_ _02636_ _01452_ vssd1 vssd1 vccd1 vccd1 _02637_ sky130_fd_sc_hd__a211oi_2
XANTENNA__10021__X _04940_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1072 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07043__A net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06637_ _01584_ _01585_ _01586_ _01587_ net777 net793 vssd1 vssd1 vccd1 vccd1 _01588_
+ sky130_fd_sc_hd__mux4_1
X_09425_ _04342_ _04343_ _04339_ vssd1 vssd1 vccd1 vccd1 _04344_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_19_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout247_X net247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout626_A net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12234__B1 net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09356_ _04058_ _04060_ net476 vssd1 vssd1 vccd1 vccd1 _04275_ sky130_fd_sc_hd__mux2_1
X_06568_ final_design.cpu.reg_window\[157\] final_design.cpu.reg_window\[189\] net949
+ vssd1 vssd1 vccd1 vccd1 _01519_ sky130_fd_sc_hd__mux2_1
XANTENNA__07336__S0 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_1819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08307_ _02157_ net598 vssd1 vssd1 vccd1 vccd1 _03258_ sky130_fd_sc_hd__and2_1
X_09287_ net496 _04097_ _04205_ vssd1 vssd1 vccd1 vccd1 _04206_ sky130_fd_sc_hd__or3_1
XANTENNA__12095__S net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout414_X net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06499_ _01446_ _01447_ _01448_ _01449_ net772 net783 vssd1 vssd1 vccd1 vccd1 _01450_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_7_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08238_ final_design.cpu.reg_window\[523\] final_design.cpu.reg_window\[555\] net826
+ vssd1 vssd1 vccd1 vccd1 _03189_ sky130_fd_sc_hd__mux2_1
X_12800__31 clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 net1341 sky130_fd_sc_hd__inv_2
XANTENNA__13733__CLK clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08169_ final_design.cpu.reg_window\[975\] final_design.cpu.reg_window\[1007\] net811
+ vssd1 vssd1 vccd1 vccd1 _03120_ sky130_fd_sc_hd__mux2_1
X_10200_ net1052 net35 vssd1 vssd1 vccd1 vccd1 _05089_ sky130_fd_sc_hd__nor2_1
XFILLER_0_82_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11180_ net647 net239 vssd1 vssd1 vccd1 vccd1 _05891_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout783_X net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10131_ final_design.VGA_data_control.v_count\[0\] _01399_ _05000_ _01401_ vssd1
+ vssd1 vccd1 vccd1 _05036_ sky130_fd_sc_hd__o31a_1
XFILLER_0_30_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11439__S net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08684__A_N _03617_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10062_ _04249_ _04252_ _04356_ _04358_ vssd1 vssd1 vccd1 vccd1 _04981_ sky130_fd_sc_hd__o22a_1
XANTENNA__09705__A2 net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout950_X net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08064__S1 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07716__A1 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13113__CLK clknet_leaf_52_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13821_ clknet_leaf_1_clk _01052_ net1078 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[809\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12068__A3 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13752_ clknet_leaf_65_clk _00983_ net1076 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[740\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12473__B1 net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10964_ _05689_ _05691_ vssd1 vssd1 vccd1 vccd1 _05692_ sky130_fd_sc_hd__nor2_1
XANTENNA__07575__S0 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12703_ _06341_ _06343_ _06338_ vssd1 vssd1 vccd1 vccd1 _06344_ sky130_fd_sc_hd__a21oi_2
XTAP_TAPCELL_ROW_14_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13683_ clknet_leaf_38_clk _00914_ net1206 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[671\]
+ sky130_fd_sc_hd__dfrtp_1
X_10895_ _05606_ _05623_ _05625_ net1005 vssd1 vssd1 vccd1 vccd1 _05626_ sky130_fd_sc_hd__a211oi_1
XANTENNA__13263__CLK clknet_leaf_43_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11902__S net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07888__A _01722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12634_ _06304_ net1555 net980 vssd1 vssd1 vccd1 vccd1 _01319_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12225__B1 net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06792__A net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11579__A2 net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12565_ net1398 _06287_ _06286_ vssd1 vssd1 vccd1 vccd1 _01267_ sky130_fd_sc_hd__mux2_1
XANTENNA__12240__A3 net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11203__A net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11516_ net2143 net208 net521 vssd1 vssd1 vccd1 vccd1 _00385_ sky130_fd_sc_hd__mux2_1
X_12496_ _06156_ net354 net332 net2099 vssd1 vssd1 vccd1 vccd1 _01202_ sky130_fd_sc_hd__a22o_1
X_14235_ net1289 vssd1 vssd1 vccd1 vccd1 gpio_out[13] sky130_fd_sc_hd__buf_2
XFILLER_0_80_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11447_ net229 net2251 net307 vssd1 vssd1 vccd1 vccd1 _00340_ sky130_fd_sc_hd__mux2_1
XANTENNA__10539__B1 net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14166_ clknet_leaf_18_clk _01340_ net1108 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.data_to_VGA\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_65_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06731__S net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08071__X _03022_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11378_ _01570_ net641 _06064_ net643 net658 vssd1 vssd1 vccd1 vccd1 _06065_ sky130_fd_sc_hd__a221o_1
XFILLER_0_61_1739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10329_ net1522 net1011 net988 final_design.data_from_mem\[14\] vssd1 vssd1 vccd1
+ vccd1 _00086_ sky130_fd_sc_hd__a22o_1
X_13117_ clknet_leaf_2_clk _00348_ net1068 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[105\]
+ sky130_fd_sc_hd__dfrtp_1
X_14097_ clknet_leaf_9_clk _01294_ net1104 vssd1 vssd1 vccd1 vccd1 final_design.reqhand.instruction\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09157__A0 net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13048_ clknet_leaf_62_clk _00279_ net1119 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[36\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_33_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11592__B net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10489__A net1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06930__A2 _01498_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13606__CLK clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07540_ final_design.cpu.reg_window\[799\] final_design.cpu.reg_window\[831\] net939
+ vssd1 vssd1 vccd1 vccd1 _02491_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11267__A1 final_design.data_from_mem\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_1857 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07471_ _02420_ _02421_ vssd1 vssd1 vccd1 vccd1 _02422_ sky130_fd_sc_hd__nor2_4
XFILLER_0_53_1267 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_27_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11812__S net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06422_ final_design.data_from_mem\[4\] vssd1 vssd1 vccd1 vccd1 _01377_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09210_ _02867_ _02897_ vssd1 vssd1 vccd1 vccd1 _04129_ sky130_fd_sc_hd__nor2_1
XANTENNA__12216__B1 net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08393__S net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13756__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09141_ net533 net532 net530 net529 net456 net466 vssd1 vssd1 vccd1 vccd1 _04060_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_44_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09072_ _02242_ _02436_ net619 vssd1 vssd1 vccd1 vccd1 _03998_ sky130_fd_sc_hd__a21o_1
XFILLER_0_47_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08023_ final_design.cpu.reg_window\[19\] final_design.cpu.reg_window\[51\] net830
+ vssd1 vssd1 vccd1 vccd1 _02974_ sky130_fd_sc_hd__mux2_1
Xhold700 final_design.cpu.reg_window\[398\] vssd1 vssd1 vccd1 vccd1 net2042 sky130_fd_sc_hd__dlygate4sd3_1
Xhold711 final_design.cpu.reg_window\[1005\] vssd1 vssd1 vccd1 vccd1 net2053 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout207_A net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold722 final_design.cpu.reg_window\[577\] vssd1 vssd1 vccd1 vccd1 net2064 sky130_fd_sc_hd__dlygate4sd3_1
Xhold733 final_design.cpu.reg_window\[466\] vssd1 vssd1 vccd1 vccd1 net2075 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09935__A2 _04619_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold744 final_design.cpu.reg_window\[949\] vssd1 vssd1 vccd1 vccd1 net2086 sky130_fd_sc_hd__dlygate4sd3_1
Xhold755 final_design.cpu.reg_window\[877\] vssd1 vssd1 vccd1 vccd1 net2097 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold766 final_design.cpu.reg_window\[481\] vssd1 vssd1 vccd1 vccd1 net2108 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07946__A1 net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold777 final_design.cpu.reg_window\[882\] vssd1 vssd1 vccd1 vccd1 net2119 sky130_fd_sc_hd__dlygate4sd3_1
Xhold788 final_design.cpu.reg_window\[189\] vssd1 vssd1 vccd1 vccd1 net2130 sky130_fd_sc_hd__dlygate4sd3_1
Xhold799 final_design.cpu.reg_window\[353\] vssd1 vssd1 vccd1 vccd1 net2141 sky130_fd_sc_hd__dlygate4sd3_1
X_09974_ net491 _04487_ _04892_ vssd1 vssd1 vccd1 vccd1 _04893_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout1116_A net1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13136__CLK clknet_leaf_34_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_33_clk_A clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08925_ final_design.CPU_instr_adr\[23\] _03796_ vssd1 vssd1 vccd1 vccd1 _03868_
+ sky130_fd_sc_hd__nor2_1
XANTENNA__09699__A1 net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout197_X net197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout576_A _05868_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07980__B net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08856_ _01510_ _02476_ vssd1 vssd1 vccd1 vccd1 _03806_ sky130_fd_sc_hd__xnor2_1
X_07807_ final_design.cpu.reg_window\[665\] final_design.cpu.reg_window\[697\] net850
+ vssd1 vssd1 vccd1 vccd1 _02758_ sky130_fd_sc_hd__mux2_1
X_08787_ _03684_ _03737_ _03681_ vssd1 vssd1 vccd1 vccd1 _03738_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout364_X net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout743_A _01476_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13286__CLK clknet_leaf_51_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_48_clk_A clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11258__A1 net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07044__Y _01995_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08087__A_N _01750_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07738_ final_design.cpu.reg_window\[986\] final_design.cpu.reg_window\[1018\] net863
+ vssd1 vssd1 vccd1 vccd1 _02689_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout910_A net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07669_ final_design.cpu.reg_window\[158\] final_design.cpu.reg_window\[190\] net853
+ vssd1 vssd1 vccd1 vccd1 _02620_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout629_X net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09408_ _04325_ _04326_ vssd1 vssd1 vccd1 vccd1 _04327_ sky130_fd_sc_hd__or2_1
XFILLER_0_3_1717 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10680_ _05418_ _05420_ vssd1 vssd1 vccd1 vccd1 _05421_ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_1897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12207__B1 net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12758__B2 final_design.VGA_adr\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09339_ _04103_ _04257_ net462 vssd1 vssd1 vccd1 vccd1 _04258_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12222__A3 net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12350_ _06234_ net500 net361 net2200 vssd1 vssd1 vccd1 vccd1 _01062_ sky130_fd_sc_hd__a22o_1
XFILLER_0_23_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11430__A1 net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_938 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout998_X net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06988__A2 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11301_ net432 net573 _05997_ net317 net1576 vssd1 vssd1 vccd1 vccd1 _00293_ sky130_fd_sc_hd__a32o_1
XANTENNA__11981__A2 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12281_ net574 _06211_ net509 net371 net1782 vssd1 vssd1 vccd1 vccd1 _00996_ sky130_fd_sc_hd__a32o_1
X_14020_ clknet_leaf_54_clk _01251_ net1179 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[1008\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07647__S net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11232_ final_design.data_from_mem\[11\] _05914_ _05917_ vssd1 vssd1 vccd1 vccd1
+ _05936_ sky130_fd_sc_hd__a21o_1
XANTENNA__11677__B net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13091__RESET_B net1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09482__S0 net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11163_ net648 net569 net242 vssd1 vssd1 vccd1 vccd1 _05876_ sky130_fd_sc_hd__and3_1
XFILLER_0_30_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09139__A0 net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10114_ net1051 _05023_ _05025_ vssd1 vssd1 vccd1 vccd1 final_design.vga.v_next_count\[4\]
+ sky130_fd_sc_hd__a21oi_1
X_11094_ _05798_ _05815_ vssd1 vssd1 vccd1 vccd1 _05816_ sky130_fd_sc_hd__nand2_1
XANTENNA__14061__CLK clknet_leaf_15_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12289__A3 net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10045_ _04632_ _04634_ _04421_ _04423_ vssd1 vssd1 vccd1 vccd1 _04964_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__13629__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10801__S net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08478__S net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold60 net128 vssd1 vssd1 vccd1 vccd1 net1402 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07382__S net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold71 final_design.VGA_data_control.data_to_VGA\[7\] vssd1 vssd1 vccd1 vccd1 net1413
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold82 final_design.reqhand.instruction\[26\] vssd1 vssd1 vccd1 vccd1 net1424 sky130_fd_sc_hd__dlygate4sd3_1
Xhold93 net140 vssd1 vssd1 vccd1 vccd1 net1435 sky130_fd_sc_hd__dlygate4sd3_1
X_13804_ clknet_leaf_46_clk _01035_ net1217 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[792\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_19_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11996_ _06198_ net280 net400 net2151 vssd1 vssd1 vccd1 vccd1 _00727_ sky130_fd_sc_hd__a22o_1
XANTENNA__08114__B2 net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13779__CLK clknet_leaf_39_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13735_ clknet_leaf_63_clk _00966_ net1120 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[723\]
+ sky130_fd_sc_hd__dfrtp_1
X_10947_ _05632_ _05653_ _05652_ vssd1 vssd1 vccd1 vccd1 _05675_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_50_1407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09862__A1 net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06676__A1 net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10472__A2 _04805_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06726__S net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13666_ clknet_leaf_11_clk _00897_ net1067 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[654\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_45_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10878_ net81 net1046 vssd1 vssd1 vccd1 vccd1 _05609_ sky130_fd_sc_hd__and2_1
XFILLER_0_6_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_45_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_41_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12617_ net2528 final_design.reqhand.data_from_UART\[3\] _05080_ vssd1 vssd1 vccd1
+ vccd1 _01310_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_41_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13597_ clknet_leaf_2_clk _00828_ net1068 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[585\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12213__A3 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_7_Left_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11421__A1 net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12548_ _06211_ net351 net325 net2183 vssd1 vssd1 vccd1 vccd1 _01252_ sky130_fd_sc_hd__a22o_1
XANTENNA__12463__S net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_2 _01752_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12479_ _06139_ net344 net330 net2523 vssd1 vssd1 vccd1 vccd1 _01185_ sky130_fd_sc_hd__a22o_1
XFILLER_0_65_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12791__22 clknet_leaf_30_clk vssd1 vssd1 vccd1 vccd1 net1332 sky130_fd_sc_hd__inv_2
XANTENNA__09378__B1 _04223_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14218_ net1276 vssd1 vssd1 vccd1 vccd1 gpio_oeb[30] sky130_fd_sc_hd__buf_2
XANTENNA__13159__CLK clknet_leaf_62_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_1683 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08242__A _02097_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11724__A2 net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14149_ clknet_leaf_15_clk _01323_ net1107 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.data_to_VGA\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09057__B net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout509 net515 vssd1 vssd1 vccd1 vccd1 net509 sky130_fd_sc_hd__buf_2
XFILLER_0_67_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06971_ _01918_ _01919_ _01920_ _01921_ net773 net791 vssd1 vssd1 vccd1 vccd1 _01922_
+ sky130_fd_sc_hd__mux4_1
X_08710_ _01359_ _01599_ vssd1 vssd1 vccd1 vccd1 _03661_ sky130_fd_sc_hd__nand2_1
XFILLER_0_59_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09690_ net493 _04338_ vssd1 vssd1 vccd1 vccd1 _04609_ sky130_fd_sc_hd__nand2_1
Xfanout1080 net1085 vssd1 vssd1 vccd1 vccd1 net1080 sky130_fd_sc_hd__clkbuf_2
X_08641_ _03030_ _03591_ vssd1 vssd1 vccd1 vccd1 _03592_ sky130_fd_sc_hd__nand2_1
Xfanout1091 net1092 vssd1 vssd1 vccd1 vccd1 net1091 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_1_238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_1_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10012__A net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08572_ _02425_ net612 vssd1 vssd1 vccd1 vccd1 _03523_ sky130_fd_sc_hd__nor2_4
XANTENNA__09527__B1_N _04223_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07523_ _01601_ _02473_ _01571_ vssd1 vssd1 vccd1 vccd1 _02474_ sky130_fd_sc_hd__a21o_1
XFILLER_0_72_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07454_ _02401_ _02402_ _02403_ _02404_ net765 net786 vssd1 vssd1 vccd1 vccd1 _02405_
+ sky130_fd_sc_hd__mux4_2
XANTENNA__10463__A2 net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11660__A1 net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06405_ final_design.CPU_instr_adr\[26\] vssd1 vssd1 vccd1 vccd1 _01360_ sky130_fd_sc_hd__inv_2
XFILLER_0_57_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07385_ final_design.cpu.reg_window\[386\] final_design.cpu.reg_window\[418\] net918
+ vssd1 vssd1 vccd1 vccd1 _02336_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout324_A net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1066_A net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09124_ _01409_ net992 vssd1 vssd1 vccd1 vccd1 _04043_ sky130_fd_sc_hd__nand2_1
XANTENNA__11412__A1 net242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_1436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09055_ _03725_ _03727_ vssd1 vssd1 vccd1 vccd1 _03983_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_5_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11963__A2 net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12373__S net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1233_A net1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07467__S net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08006_ final_design.cpu.reg_window\[592\] final_design.cpu.reg_window\[624\] net843
+ vssd1 vssd1 vccd1 vccd1 _02957_ sky130_fd_sc_hd__mux2_1
Xhold530 final_design.cpu.reg_window\[642\] vssd1 vssd1 vccd1 vccd1 net1872 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14084__CLK clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold541 final_design.cpu.reg_window\[487\] vssd1 vssd1 vccd1 vccd1 net1883 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout693_A net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold552 final_design.cpu.reg_window\[360\] vssd1 vssd1 vccd1 vccd1 net1894 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap260 _03585_ vssd1 vssd1 vccd1 vccd1 net260 sky130_fd_sc_hd__buf_2
Xhold563 final_design.cpu.reg_window\[432\] vssd1 vssd1 vccd1 vccd1 net1905 sky130_fd_sc_hd__dlygate4sd3_1
Xhold574 final_design.cpu.reg_window\[685\] vssd1 vssd1 vccd1 vccd1 net1916 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09384__A3 net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold585 net141 vssd1 vssd1 vccd1 vccd1 net1927 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_55_2090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold596 final_design.cpu.reg_window\[938\] vssd1 vssd1 vccd1 vccd1 net1938 sky130_fd_sc_hd__dlygate4sd3_1
X_09957_ _03557_ _04875_ _04874_ _03652_ vssd1 vssd1 vccd1 vccd1 _04876_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_70_2588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout860_A net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout958_A _04041_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_2599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout579_X net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08908_ _03798_ _03852_ vssd1 vssd1 vccd1 vccd1 _03853_ sky130_fd_sc_hd__or2_1
XFILLER_0_77_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_1532 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09888_ net79 net725 _04805_ vssd1 vssd1 vccd1 vccd1 _04807_ sky130_fd_sc_hd__or3_1
XANTENNA__07778__S0 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08839_ final_design.CPU_instr_adr\[13\] final_design.CPU_instr_adr\[12\] _03789_
+ vssd1 vssd1 vccd1 vccd1 _03790_ sky130_fd_sc_hd__and3_1
XANTENNA__13921__CLK clknet_leaf_47_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout746_X net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12428__B1 net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11850_ _06100_ net284 net518 net2434 vssd1 vssd1 vccd1 vccd1 _00600_ sky130_fd_sc_hd__a22o_1
XFILLER_0_68_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10801_ final_design.CPU_instr_adr\[17\] _03919_ net1060 vssd1 vssd1 vccd1 vccd1
+ _05536_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout913_X net913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11781_ net2315 net412 _06231_ net431 vssd1 vssd1 vccd1 vccd1 _00539_ sky130_fd_sc_hd__a22o_1
XANTENNA__11305__X _06001_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13520_ clknet_leaf_33_clk _00751_ net1238 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[508\]
+ sky130_fd_sc_hd__dfrtp_1
X_10732_ _05464_ _05468_ vssd1 vssd1 vccd1 vccd1 _05470_ sky130_fd_sc_hd__nor2_1
XFILLER_0_3_1558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13451_ clknet_leaf_38_clk _00682_ net1190 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[439\]
+ sky130_fd_sc_hd__dfrtp_1
X_10663_ _05402_ _05404_ vssd1 vssd1 vccd1 vccd1 _05405_ sky130_fd_sc_hd__xor2_1
XFILLER_0_14_1582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12402_ _06100_ net348 net339 net2203 vssd1 vssd1 vccd1 vccd1 _01112_ sky130_fd_sc_hd__a22o_1
XFILLER_0_49_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07607__B1 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input87_A memory_size[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10594_ final_design.CPU_instr_adr\[7\] _03995_ net1058 vssd1 vssd1 vccd1 vccd1 _05339_
+ sky130_fd_sc_hd__mux2_1
X_13382_ clknet_leaf_52_clk _00613_ net1174 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[370\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13301__CLK clknet_leaf_56_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11954__A2 net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12333_ _06229_ net500 net361 net1975 vssd1 vssd1 vccd1 vccd1 _01045_ sky130_fd_sc_hd__a22o_1
Xclkbuf_3_3_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_3_3_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_10_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12264_ net231 net2398 net368 vssd1 vssd1 vccd1 vccd1 _00979_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_1845 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11706__A2 net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14003_ clknet_leaf_40_clk _01234_ net1210 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[991\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11215_ net646 net559 net220 vssd1 vssd1 vccd1 vccd1 _05922_ sky130_fd_sc_hd__and3_1
XANTENNA__13451__CLK clknet_leaf_38_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12195_ net1914 net176 net383 vssd1 vssd1 vccd1 vccd1 _00914_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_1889 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11146_ final_design.CPU_instr_adr\[1\] net731 _05859_ vssd1 vssd1 vccd1 vccd1 _05860_
+ sky130_fd_sc_hd__o21ai_1
X_11077_ _04249_ net252 _04990_ vssd1 vssd1 vccd1 vccd1 _05799_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_37_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10028_ _04342_ _04836_ _04946_ net261 vssd1 vssd1 vccd1 vccd1 _04947_ sky130_fd_sc_hd__o211a_1
XFILLER_0_56_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10142__A1 net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_47_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1903 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12458__S net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11979_ _06181_ net288 net407 net2170 vssd1 vssd1 vccd1 vccd1 _00712_ sky130_fd_sc_hd__a22o_1
XFILLER_0_15_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13718_ clknet_leaf_59_clk _00949_ net1138 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[706\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11642__A1 net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07941__S0 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13649_ clknet_leaf_35_clk _00880_ net1237 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[637\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07170_ final_design.cpu.reg_window\[650\] final_design.cpu.reg_window\[682\] net896
+ vssd1 vssd1 vccd1 vccd1 _02121_ sky130_fd_sc_hd__mux2_1
XANTENNA__08497__S1 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11945__A2 net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12193__S net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1901 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07287__S net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout306 net307 vssd1 vssd1 vccd1 vccd1 net306 sky130_fd_sc_hd__clkbuf_8
Xfanout317 _05851_ vssd1 vssd1 vccd1 vccd1 net317 sky130_fd_sc_hd__buf_4
X_09811_ _03259_ net441 net438 _03261_ _04729_ vssd1 vssd1 vccd1 vccd1 _04730_ sky130_fd_sc_hd__o221a_1
Xfanout328 net329 vssd1 vssd1 vccd1 vccd1 net328 sky130_fd_sc_hd__buf_4
Xfanout339 net341 vssd1 vssd1 vccd1 vccd1 net339 sky130_fd_sc_hd__buf_4
XANTENNA__10381__A1 net25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload11_A clknet_leaf_63_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09742_ _03198_ _03571_ _04495_ _03231_ net321 vssd1 vssd1 vccd1 vccd1 _04661_ sky130_fd_sc_hd__a221oi_1
X_06954_ final_design.cpu.reg_window\[529\] final_design.cpu.reg_window\[561\] net925
+ vssd1 vssd1 vccd1 vccd1 _01905_ sky130_fd_sc_hd__mux2_1
XANTENNA__09523__A0 _04233_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09673_ _02837_ _04352_ _04591_ vssd1 vssd1 vccd1 vccd1 _04592_ sky130_fd_sc_hd__a21oi_1
X_06885_ _01832_ _01833_ _01834_ _01835_ net769 net790 vssd1 vssd1 vccd1 vccd1 _01836_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout274_A net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11330__B1 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08624_ _03262_ _03574_ vssd1 vssd1 vccd1 vccd1 _03575_ sky130_fd_sc_hd__nor2_1
XANTENNA__11780__B net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08555_ net710 _03505_ vssd1 vssd1 vccd1 vccd1 _03506_ sky130_fd_sc_hd__or2_1
XANTENNA__12368__S net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout441_A net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08629__A2 _03065_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_1801 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1183_A net1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout539_A _02058_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07506_ _01911_ _02456_ _01912_ vssd1 vssd1 vccd1 vccd1 _02457_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_82_2993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_2370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08486_ net717 _03436_ vssd1 vssd1 vccd1 vccd1 _03437_ sky130_fd_sc_hd__or2_1
XANTENNA__13324__CLK clknet_leaf_46_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1845 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10396__B net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07051__A _01996_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07437_ net760 _02387_ vssd1 vssd1 vccd1 vccd1 _02388_ sky130_fd_sc_hd__or2_2
XFILLER_0_0_1709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1889 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout327_X net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout706_A _01752_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1069_X net1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07368_ final_design.cpu.reg_window\[707\] final_design.cpu.reg_window\[739\] net908
+ vssd1 vssd1 vccd1 vccd1 _02319_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09107_ _03715_ _03717_ vssd1 vssd1 vccd1 vccd1 _04028_ sky130_fd_sc_hd__xor2_1
XANTENNA__06499__S0 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07299_ final_design.cpu.reg_window\[261\] final_design.cpu.reg_window\[293\] net919
+ vssd1 vssd1 vccd1 vccd1 _02250_ sky130_fd_sc_hd__mux2_1
XANTENNA__13474__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_2141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09038_ _03788_ _03967_ vssd1 vssd1 vccd1 vccd1 _03968_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_57_2152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_2786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_2163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_2797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_2005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout696_X net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_2016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_2027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold360 final_design.cpu.reg_window\[978\] vssd1 vssd1 vccd1 vccd1 net1702 sky130_fd_sc_hd__dlygate4sd3_1
Xhold371 final_design.cpu.reg_window\[963\] vssd1 vssd1 vccd1 vccd1 net1713 sky130_fd_sc_hd__dlygate4sd3_1
Xhold382 final_design.cpu.reg_window\[886\] vssd1 vssd1 vccd1 vccd1 net1724 sky130_fd_sc_hd__dlygate4sd3_1
X_11000_ net967 _05725_ vssd1 vssd1 vccd1 vccd1 _05726_ sky130_fd_sc_hd__nand2_1
Xhold393 final_design.cpu.reg_window\[879\] vssd1 vssd1 vccd1 vccd1 net1735 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12361__A2 net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09762__B1 net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10372__B2 final_design.data_from_mem\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout840 net841 vssd1 vssd1 vccd1 vccd1 net840 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11447__S net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout851 net852 vssd1 vssd1 vccd1 vccd1 net851 sky130_fd_sc_hd__clkbuf_4
Xfanout862 net865 vssd1 vssd1 vccd1 vccd1 net862 sky130_fd_sc_hd__buf_4
XANTENNA__09425__B _04343_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout873 _01818_ vssd1 vssd1 vccd1 vccd1 net873 sky130_fd_sc_hd__clkbuf_4
Xfanout884 net885 vssd1 vssd1 vccd1 vccd1 net884 sky130_fd_sc_hd__buf_6
XANTENNA__09514__B1 net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_5_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07226__A net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout895 net896 vssd1 vssd1 vccd1 vccd1 net895 sky130_fd_sc_hd__clkbuf_4
X_12951_ clknet_leaf_29_clk _00189_ net1195 vssd1 vssd1 vccd1 vccd1 net108 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_5_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1060 final_design.cpu.reg_window\[252\] vssd1 vssd1 vccd1 vccd1 net2402 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11321__B1 _06014_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1071 final_design.cpu.reg_window\[609\] vssd1 vssd1 vccd1 vccd1 net2413 sky130_fd_sc_hd__dlygate4sd3_1
X_11902_ net204 net2381 net274 vssd1 vssd1 vccd1 vccd1 _00644_ sky130_fd_sc_hd__mux2_1
Xhold1082 final_design.cpu.reg_window\[226\] vssd1 vssd1 vccd1 vccd1 net2424 sky130_fd_sc_hd__dlygate4sd3_1
X_12882_ clknet_leaf_17_clk _00120_ net1114 vssd1 vssd1 vccd1 vccd1 final_design.data_from_mem\[16\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_38_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1093 final_design.cpu.reg_window\[108\] vssd1 vssd1 vccd1 vccd1 net2435 sky130_fd_sc_hd__dlygate4sd3_1
X_11833_ net195 net2146 net265 vssd1 vssd1 vccd1 vccd1 _00585_ sky130_fd_sc_hd__mux2_1
XANTENNA__09817__A1 _04378_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12416__A3 net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08176__S0 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11764_ net182 net2511 net418 vssd1 vssd1 vccd1 vccd1 _00527_ sky130_fd_sc_hd__mux2_1
XANTENNA__09293__A2 net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07923__S0 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13503_ clknet_leaf_7_clk _00734_ net1135 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[491\]
+ sky130_fd_sc_hd__dfrtp_1
X_10715_ net958 _05451_ _05453_ net955 vssd1 vssd1 vccd1 vccd1 _05454_ sky130_fd_sc_hd__o22a_1
XFILLER_0_82_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11695_ net212 net626 vssd1 vssd1 vccd1 vccd1 _06206_ sky130_fd_sc_hd__and2_1
XFILLER_0_71_819 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13817__CLK clknet_leaf_54_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13434_ clknet_leaf_58_clk _00665_ net1128 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[422\]
+ sky130_fd_sc_hd__dfrtp_1
X_10646_ _04767_ net250 vssd1 vssd1 vccd1 vccd1 _05388_ sky130_fd_sc_hd__nor2_1
XFILLER_0_3_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08491__S net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11927__A2 net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13365_ clknet_leaf_55_clk _00596_ net1146 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[353\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10577_ net801 _05320_ _05322_ net961 vssd1 vssd1 vccd1 vccd1 _05323_ sky130_fd_sc_hd__o22a_1
XANTENNA__08504__B net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12316_ net1677 net199 net365 vssd1 vssd1 vccd1 vccd1 _01030_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12841__CLK clknet_leaf_19_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13296_ clknet_leaf_33_clk _00527_ net1232 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[284\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13967__CLK clknet_leaf_42_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12247_ net572 _06176_ net501 _06273_ vssd1 vssd1 vccd1 vccd1 _00963_ sky130_fd_sc_hd__a31o_1
XANTENNA__06799__X _01750_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08100__S0 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12352__A2 net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11865__B net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12178_ net2030 net208 net380 vssd1 vssd1 vccd1 vccd1 _00897_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_79_Left_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10363__B2 final_design.data_from_mem\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14140__1246 vssd1 vssd1 vccd1 vccd1 _14140__1246/HI net1246 sky130_fd_sc_hd__conb_1
XFILLER_0_78_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11129_ net804 _05839_ vssd1 vssd1 vccd1 vccd1 _05844_ sky130_fd_sc_hd__or2_1
XFILLER_0_3_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06670_ final_design.cpu.reg_window\[538\] final_design.cpu.reg_window\[570\] net941
+ vssd1 vssd1 vccd1 vccd1 _01621_ sky130_fd_sc_hd__mux2_1
XANTENNA__13347__CLK clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12188__S net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08340_ net534 _03289_ vssd1 vssd1 vccd1 vccd1 _03291_ sky130_fd_sc_hd__or2_1
XFILLER_0_58_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09284__A2 net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08271_ _03218_ _03219_ _03220_ _03221_ net675 net691 vssd1 vssd1 vccd1 vccd1 _03222_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_69_1829 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13497__CLK clknet_leaf_56_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11820__S net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07222_ final_design.cpu.reg_window\[648\] final_design.cpu.reg_window\[680\] net889
+ vssd1 vssd1 vccd1 vccd1 _02173_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07153_ final_design.cpu.reg_window\[330\] final_design.cpu.reg_window\[362\] net906
+ vssd1 vssd1 vccd1 vccd1 _02104_ sky130_fd_sc_hd__mux2_1
XANTENNA__07047__A1 final_design.data_from_mem\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12591__A2 net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07084_ final_design.cpu.reg_window\[268\] final_design.cpu.reg_window\[300\] net907
+ vssd1 vssd1 vccd1 vccd1 _02035_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_1873 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_1715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09744__A0 net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1029_A net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12343__A2 net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06502__X _01453_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout391_A _06265_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10354__A1 net27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10354__B2 final_design.data_from_mem\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06869__B _01468_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11551__B1 net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout489_A net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14122__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07986_ _01939_ net613 vssd1 vssd1 vccd1 vccd1 _02937_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_2_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09725_ _01717_ net551 net550 _01815_ net453 net463 vssd1 vssd1 vccd1 vccd1 _04644_
+ sky130_fd_sc_hd__mux4_1
X_06937_ final_design.cpu.reg_window\[273\] final_design.cpu.reg_window\[305\] net930
+ vssd1 vssd1 vccd1 vccd1 _01888_ sky130_fd_sc_hd__mux2_1
XANTENNA__11303__B1 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout277_X net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout656_A _05142_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09656_ net80 _04189_ net81 vssd1 vssd1 vccd1 vccd1 _04575_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_65_2410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_2421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06868_ net742 net873 vssd1 vssd1 vccd1 vccd1 _01819_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_65_2432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_2443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08607_ _03555_ _03556_ _03488_ vssd1 vssd1 vccd1 vccd1 _03558_ sky130_fd_sc_hd__a21o_1
XANTENNA__12098__S net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout823_A net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09587_ _03164_ _04505_ _03162_ vssd1 vssd1 vccd1 vccd1 _04506_ sky130_fd_sc_hd__a21oi_1
X_06799_ net883 _01731_ _01737_ _01743_ _01749_ vssd1 vssd1 vccd1 vccd1 _01750_ sky130_fd_sc_hd__o32a_4
XANTENNA_fanout444_X net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_2307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10409__A2 net1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08538_ final_design.cpu.reg_window\[321\] final_design.cpu.reg_window\[353\] net838
+ vssd1 vssd1 vccd1 vccd1 _03489_ sky130_fd_sc_hd__mux2_1
XANTENNA__10200__A net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07905__S0 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11176__A_N final_design.reqhand.data_from_UART\[4\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_4_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08469_ net609 _03415_ _03416_ _02294_ vssd1 vssd1 vccd1 vccd1 _03420_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_18_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout709_X net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10500_ _05233_ _05246_ _05244_ vssd1 vssd1 vccd1 vccd1 _05249_ sky130_fd_sc_hd__o21bai_2
XANTENNA__09027__A2 net1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwire526 _03129_ vssd1 vssd1 vccd1 vccd1 net526 sky130_fd_sc_hd__buf_4
X_11480_ _06017_ net2504 net308 vssd1 vssd1 vccd1 vccd1 _00360_ sky130_fd_sc_hd__mux2_1
XANTENNA__06824__S net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12864__CLK clknet_leaf_19_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_2214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_59_2225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_2859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_2236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12031__A1 net240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10431_ _03613_ _05180_ vssd1 vssd1 vccd1 vccd1 _05199_ sky130_fd_sc_hd__or2_2
XANTENNA__07133__S1 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12582__A2 net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13150_ clknet_leaf_13_clk _00381_ net1088 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[138\]
+ sky130_fd_sc_hd__dfrtp_1
X_10362_ net4 net1024 net1006 final_design.data_from_mem\[11\] vssd1 vssd1 vccd1 vccd1
+ _00115_ sky130_fd_sc_hd__o22a_1
X_12101_ net2169 net237 net389 vssd1 vssd1 vccd1 vccd1 _00825_ sky130_fd_sc_hd__mux2_1
XANTENNA__11790__B1 net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10293_ net1048 _05146_ vssd1 vssd1 vccd1 vccd1 _05147_ sky130_fd_sc_hd__nand2_1
X_13081_ clknet_leaf_59_clk _00312_ net1143 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[69\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_1913 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12334__A2 net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12032_ net1804 net225 net399 vssd1 vssd1 vccd1 vccd1 _00760_ sky130_fd_sc_hd__mux2_1
XANTENNA__11685__B net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold190 final_design.cpu.reg_window\[990\] vssd1 vssd1 vccd1 vccd1 net1532 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09155__B net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10896__A2 net1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout670 _04989_ vssd1 vssd1 vccd1 vccd1 net670 sky130_fd_sc_hd__clkbuf_4
Xfanout681 net690 vssd1 vssd1 vccd1 vccd1 net681 sky130_fd_sc_hd__buf_4
Xfanout692 _01753_ vssd1 vssd1 vccd1 vccd1 net692 sky130_fd_sc_hd__clkbuf_8
X_13983_ clknet_leaf_7_clk _01214_ net1131 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[971\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11905__S net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12934_ clknet_leaf_29_clk _00172_ net1195 vssd1 vssd1 vccd1 vccd1 net158 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_1023 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_16_Right_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12865_ clknet_leaf_20_clk _00103_ net1158 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.ready_data\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11206__A net245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11816_ net224 net2226 net265 vssd1 vssd1 vccd1 vccd1 _00568_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_1917 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12270__A1 net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11747_ net215 net2124 net417 vssd1 vssd1 vccd1 vccd1 _00510_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_1376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07372__S1 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06734__S net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11678_ net564 net421 _06197_ net295 net2016 vssd1 vssd1 vccd1 vccd1 _00470_ sky130_fd_sc_hd__a32o_1
X_13417_ clknet_leaf_37_clk _00648_ net1229 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[405\]
+ sky130_fd_sc_hd__dfrtp_1
X_10629_ net98 final_design.VGA_adr\[6\] _05370_ vssd1 vssd1 vccd1 vccd1 _05372_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_25_Right_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10033__B1 net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13348_ clknet_leaf_52_clk _00579_ net1174 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[336\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14145__CLK clknet_leaf_18_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13279_ clknet_leaf_7_clk _00510_ net1135 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[267\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09726__A0 _01596_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10336__B2 final_design.data_from_mem\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07840_ final_design.cpu.reg_window\[725\] final_design.cpu.reg_window\[757\] net858
+ vssd1 vssd1 vccd1 vccd1 _02791_ sky130_fd_sc_hd__mux2_1
XANTENNA__07752__A2 _02698_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07771_ final_design.cpu.reg_window\[984\] final_design.cpu.reg_window\[1016\] net864
+ vssd1 vssd1 vccd1 vccd1 _02722_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_34_Right_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11815__S net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09510_ _04427_ _04428_ net448 vssd1 vssd1 vccd1 vccd1 _04429_ sky130_fd_sc_hd__a21o_1
X_06722_ _01669_ _01670_ _01671_ _01672_ net775 net793 vssd1 vssd1 vccd1 vccd1 _01673_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__08396__S net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06938__S1 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09441_ _02738_ _03594_ _04359_ vssd1 vssd1 vccd1 vccd1 _04360_ sky130_fd_sc_hd__a21o_1
X_06653_ final_design.cpu.reg_window\[474\] final_design.cpu.reg_window\[506\] net943
+ vssd1 vssd1 vccd1 vccd1 _01604_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_1298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09372_ _02609_ _04050_ _03605_ _02573_ _02575_ vssd1 vssd1 vccd1 vccd1 _04291_ sky130_fd_sc_hd__a2111oi_1
X_06584_ net884 _01528_ _01534_ _01521_ _01522_ vssd1 vssd1 vccd1 vccd1 _01535_ sky130_fd_sc_hd__a32oi_4
XANTENNA__12887__CLK clknet_leaf_18_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08323_ net716 _03273_ vssd1 vssd1 vccd1 vccd1 _03274_ sky130_fd_sc_hd__or2_1
XANTENNA__12261__A1 net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08560__S0 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08254_ _03201_ _03202_ _03203_ _03204_ net676 net697 vssd1 vssd1 vccd1 vccd1 _03205_
+ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_43_Right_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07205_ net881 _02148_ _02154_ _02141_ _02142_ vssd1 vssd1 vccd1 vccd1 _02156_ sky130_fd_sc_hd__a32o_2
X_08185_ final_design.cpu.reg_window\[334\] final_design.cpu.reg_window\[366\] net825
+ vssd1 vssd1 vccd1 vccd1 _03136_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout404_A net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10024__B1 net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_2701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07136_ final_design.cpu.reg_window\[587\] final_design.cpu.reg_window\[619\] net908
+ vssd1 vssd1 vccd1 vccd1 _02087_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_73_2712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07067_ final_design.cpu.reg_window\[653\] final_design.cpu.reg_window\[685\] net934
+ vssd1 vssd1 vccd1 vccd1 _02018_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12381__S net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13512__CLK clknet_leaf_41_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10327__B2 final_design.data_from_mem\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout394_X net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout773_A net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_52_Right_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_67_2505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07969_ final_design.cpu.reg_window\[849\] final_design.cpu.reg_window\[881\] net845
+ vssd1 vssd1 vccd1 vccd1 _02920_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout561_X net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout940_A net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout659_X net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09708_ _03070_ _04504_ vssd1 vssd1 vccd1 vccd1 _04627_ sky130_fd_sc_hd__nand2_1
XFILLER_0_69_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13662__CLK clknet_leaf_11_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10980_ net962 _05706_ vssd1 vssd1 vccd1 vccd1 _05707_ sky130_fd_sc_hd__or2_1
XANTENNA__09496__A2 _04086_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09639_ _02997_ net445 net442 _02994_ _04557_ vssd1 vssd1 vccd1 vccd1 _04558_ sky130_fd_sc_hd__o221a_1
XFILLER_0_70_1229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_1737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12650_ _06312_ net1471 net979 vssd1 vssd1 vccd1 vccd1 _01327_ sky130_fd_sc_hd__mux2_1
XANTENNA__14018__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11601_ net580 net423 _06156_ net304 net2087 vssd1 vssd1 vccd1 vccd1 _00434_ sky130_fd_sc_hd__a32o_1
XANTENNA__11055__A2 net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12581_ _01395_ net1001 vssd1 vssd1 vccd1 vccd1 _06296_ sky130_fd_sc_hd__nor2_1
XFILLER_0_66_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10865__A net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_61_Right_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07354__S1 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11532_ net2245 net182 net523 vssd1 vssd1 vccd1 vccd1 _00399_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_22_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14251_ net1305 vssd1 vssd1 vccd1 vccd1 gpio_out[29] sky130_fd_sc_hd__buf_2
XFILLER_0_11_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08208__B1 net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11463_ net218 net2474 net306 vssd1 vssd1 vccd1 vccd1 _00348_ sky130_fd_sc_hd__mux2_1
XANTENNA__13042__CLK clknet_leaf_39_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14168__CLK clknet_leaf_18_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13202_ clknet_leaf_39_clk _00433_ net1206 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[190\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12555__A2 net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09956__B1 _04124_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10414_ _05176_ _05180_ vssd1 vssd1 vccd1 vccd1 _05190_ sky130_fd_sc_hd__or2_4
X_14182_ clknet_leaf_29_clk _01356_ net1193 vssd1 vssd1 vccd1 vccd1 final_design.VGA_adr\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_11394_ _01507_ net641 _06078_ net644 vssd1 vssd1 vccd1 vccd1 _06079_ sky130_fd_sc_hd__a22o_1
X_13133_ clknet_leaf_45_clk _00364_ net1202 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[121\]
+ sky130_fd_sc_hd__dfrtp_1
X_10345_ net1508 net1011 net988 final_design.data_from_mem\[30\] vssd1 vssd1 vccd1
+ vccd1 _00102_ sky130_fd_sc_hd__a22o_1
XFILLER_0_24_1721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13192__CLK clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09166__A net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07982__A2 _02929_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13064_ clknet_leaf_35_clk _00295_ net1237 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[52\]
+ sky130_fd_sc_hd__dfrtp_1
X_10276_ final_design.uart.BAUD_counter\[28\] _05134_ net797 vssd1 vssd1 vccd1 vccd1
+ _05136_ sky130_fd_sc_hd__o21ai_1
XANTENNA__10318__B2 final_design.data_from_mem\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_70_Right_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07719__C1 _01596_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12015_ _06217_ net285 net402 net2133 vssd1 vssd1 vccd1 vccd1 _00746_ sky130_fd_sc_hd__a22o_1
XANTENNA__09723__A3 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_31_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11279__C1 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13966_ clknet_leaf_45_clk _01197_ net1215 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[954\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_31_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06729__S net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09105__S net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12917_ clknet_leaf_62_clk _00155_ net1123 vssd1 vssd1 vccd1 vccd1 net139 sky130_fd_sc_hd__dfrtp_1
XANTENNA__07042__S0 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13897_ clknet_leaf_33_clk _01128_ net1231 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[885\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12848_ clknet_leaf_18_clk _00086_ net1110 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.ready_data\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08944__S net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12243__A1 net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09644__C1 _04222_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08542__S0 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_25_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12546__A2 net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold904 final_design.cpu.reg_window\[268\] vssd1 vssd1 vccd1 vccd1 net2246 sky130_fd_sc_hd__dlygate4sd3_1
Xhold915 final_design.cpu.reg_window\[506\] vssd1 vssd1 vccd1 vccd1 net2257 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13535__CLK clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold926 final_design.cpu.reg_window\[493\] vssd1 vssd1 vccd1 vccd1 net2268 sky130_fd_sc_hd__dlygate4sd3_1
Xhold937 final_design.cpu.reg_window\[320\] vssd1 vssd1 vccd1 vccd1 net2279 sky130_fd_sc_hd__dlygate4sd3_1
Xhold948 final_design.cpu.reg_window\[623\] vssd1 vssd1 vccd1 vccd1 net2290 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10714__S net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold959 final_design.cpu.reg_window\[624\] vssd1 vssd1 vccd1 vccd1 net2301 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06856__S0 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09990_ _02736_ net443 vssd1 vssd1 vccd1 vccd1 _04909_ sky130_fd_sc_hd__or2_1
X_08941_ _03762_ _03881_ vssd1 vssd1 vccd1 vccd1 _03882_ sky130_fd_sc_hd__xor2_1
XFILLER_0_23_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09507__C _04157_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08872_ _03801_ _03820_ vssd1 vssd1 vccd1 vccd1 _03821_ sky130_fd_sc_hd__or2_1
XANTENNA__13685__CLK clknet_leaf_58_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1917 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07823_ final_design.cpu.reg_window\[213\] final_design.cpu.reg_window\[245\] net859
+ vssd1 vssd1 vccd1 vccd1 _02774_ sky130_fd_sc_hd__mux2_1
XANTENNA__07281__S0 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout187_A _06052_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07754_ _02704_ vssd1 vssd1 vccd1 vccd1 _02705_ sky130_fd_sc_hd__inv_2
XANTENNA__11809__B2 _06090_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06705_ net762 _01655_ vssd1 vssd1 vccd1 vccd1 _01656_ sky130_fd_sc_hd__or2_1
X_07685_ _01507_ net614 vssd1 vssd1 vccd1 vccd1 _02636_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout354_A net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1096_A net1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09424_ net493 _04205_ vssd1 vssd1 vccd1 vccd1 _04343_ sky130_fd_sc_hd__nand2_1
XFILLER_0_14_1901 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06636_ final_design.cpu.reg_window\[923\] final_design.cpu.reg_window\[955\] net943
+ vssd1 vssd1 vccd1 vccd1 _01587_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12234__A1 net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09355_ _04074_ _04264_ _04273_ _04263_ vssd1 vssd1 vccd1 vccd1 _04274_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout521_A net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13065__CLK clknet_leaf_36_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12376__S net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06567_ final_design.cpu.reg_window\[221\] final_design.cpu.reg_window\[253\] net949
+ vssd1 vssd1 vccd1 vccd1 _01518_ sky130_fd_sc_hd__mux2_1
XANTENNA__12229__X _06272_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout619_A net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_2910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08989__A1 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07336__S1 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08306_ net874 _03238_ _03244_ _03250_ _03256_ vssd1 vssd1 vccd1 vccd1 _03257_ sky130_fd_sc_hd__o32a_4
XFILLER_0_63_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09286_ net479 _04204_ vssd1 vssd1 vccd1 vccd1 _04205_ sky130_fd_sc_hd__or2_1
X_06498_ final_design.cpu.reg_window\[542\] final_design.cpu.reg_window\[574\] net931
+ vssd1 vssd1 vccd1 vccd1 _01449_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_7_clk_A clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08237_ final_design.cpu.reg_window\[587\] final_design.cpu.reg_window\[619\] net826
+ vssd1 vssd1 vccd1 vccd1 _03188_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout407_X net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12537__A2 net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1149_X net1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1612 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09938__B1 _04586_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08168_ final_design.cpu.reg_window\[783\] final_design.cpu.reg_window\[815\] net811
+ vssd1 vssd1 vccd1 vccd1 _03119_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11745__A0 net219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout890_A net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout988_A _05167_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07119_ final_design.cpu.reg_window\[459\] final_design.cpu.reg_window\[491\] net915
+ vssd1 vssd1 vccd1 vccd1 _02070_ sky130_fd_sc_hd__mux2_1
X_08099_ final_design.cpu.reg_window\[140\] final_design.cpu.reg_window\[172\] net814
+ vssd1 vssd1 vccd1 vccd1 _03050_ sky130_fd_sc_hd__mux2_1
XANTENNA__12902__CLK clknet_leaf_25_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10130_ _05002_ _05035_ final_design.v_out vssd1 vssd1 vccd1 vccd1 final_design.vga.v_next_state\[0\]
+ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout776_X net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10061_ _04325_ _04326_ _04964_ _04966_ _04979_ vssd1 vssd1 vccd1 vccd1 _04980_ sky130_fd_sc_hd__o2111a_1
XANTENNA__08374__C1 _02211_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11455__S net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13820_ clknet_leaf_5_clk _01051_ net1080 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[808\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_1861 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13751_ clknet_leaf_6_clk _00982_ net1130 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[739\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07024__S0 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10963_ net52 _05688_ vssd1 vssd1 vccd1 vccd1 _05691_ sky130_fd_sc_hd__nor2_1
XFILLER_0_15_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13408__CLK clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12702_ final_design.VGA_data_control.v_count\[5\] _06337_ _06342_ vssd1 vssd1 vccd1
+ vccd1 _06343_ sky130_fd_sc_hd__o21ai_2
XANTENNA__10484__B1 _04990_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07575__S1 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13682_ clknet_leaf_38_clk _00913_ net1189 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[670\]
+ sky130_fd_sc_hd__dfrtp_1
X_10894_ _05600_ _05621_ vssd1 vssd1 vccd1 vccd1 _05625_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_14_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12633_ final_design.VGA_data_control.ready_data\[4\] net1021 net976 final_design.data_from_mem\[4\]
+ vssd1 vssd1 vccd1 vccd1 _06304_ sky130_fd_sc_hd__a22o_1
XFILLER_0_52_1460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_1471 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08336__Y _03287_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12564_ net1052 final_design.uart.working_data\[2\] vssd1 vssd1 vccd1 vccd1 _06287_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_80_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13558__CLK clknet_leaf_61_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11984__B1 net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11515_ net1984 net209 net524 vssd1 vssd1 vccd1 vccd1 _00384_ sky130_fd_sc_hd__mux2_1
X_12495_ _06155_ net353 net332 net1929 vssd1 vssd1 vccd1 vccd1 _01201_ sky130_fd_sc_hd__a22o_1
XFILLER_0_53_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14234_ net1288 vssd1 vssd1 vccd1 vccd1 gpio_out[12] sky130_fd_sc_hd__buf_2
XANTENNA__12528__A2 net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11446_ net229 net639 vssd1 vssd1 vccd1 vccd1 _06096_ sky130_fd_sc_hd__and2_1
XFILLER_0_46_1220 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14165_ clknet_leaf_18_clk _01339_ net1116 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.data_to_VGA\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08601__B1 _02423_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09167__Y _04086_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11377_ final_design.data_from_mem\[28\] net236 net234 vssd1 vssd1 vccd1 vccd1 _06064_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_0_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13116_ clknet_leaf_3_clk _00347_ net1066 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[104\]
+ sky130_fd_sc_hd__dfrtp_1
X_10328_ net1524 net1010 net987 final_design.data_from_mem\[13\] vssd1 vssd1 vccd1
+ vccd1 _00085_ sky130_fd_sc_hd__a22o_1
X_14096_ clknet_leaf_9_clk _01293_ net1151 vssd1 vssd1 vccd1 vccd1 final_design.reqhand.instruction\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09157__A1 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13047_ clknet_leaf_5_clk _00278_ net1081 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[35\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_37_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10259_ _05124_ _05125_ vssd1 vssd1 vccd1 vccd1 _00019_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_33_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12161__A0 net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1240 net1244 vssd1 vssd1 vccd1 vccd1 net1240 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_52_1969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07843__S net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09624__A _04072_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11218__X _05924_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08117__C1 _02058_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13949_ clknet_leaf_1_clk _01180_ net1077 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[937\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10475__B1 net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07470_ _01480_ net728 net805 vssd1 vssd1 vccd1 vccd1 _02421_ sky130_fd_sc_hd__and3_2
XFILLER_0_5_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_27_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06421_ final_design.reqhand.instruction\[4\] vssd1 vssd1 vccd1 vccd1 _01376_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_27_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12216__A1 net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09140_ _04057_ _04058_ net477 vssd1 vssd1 vccd1 vccd1 _04059_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09093__B1 net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11975__B1 net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09071_ net2337 net1013 _03997_ vssd1 vssd1 vccd1 vccd1 _00218_ sky130_fd_sc_hd__a21o_1
XANTENNA__12925__CLK clknet_leaf_61_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08022_ final_design.cpu.reg_window\[83\] final_design.cpu.reg_window\[115\] net834
+ vssd1 vssd1 vccd1 vccd1 _02973_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12519__A2 net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold701 final_design.cpu.reg_window\[345\] vssd1 vssd1 vccd1 vccd1 net2043 sky130_fd_sc_hd__dlygate4sd3_1
Xhold712 final_design.cpu.reg_window\[372\] vssd1 vssd1 vccd1 vccd1 net2054 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold723 final_design.cpu.reg_window\[331\] vssd1 vssd1 vccd1 vccd1 net2065 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold734 final_design.cpu.reg_window\[263\] vssd1 vssd1 vccd1 vccd1 net2076 sky130_fd_sc_hd__dlygate4sd3_1
Xhold745 final_design.cpu.reg_window\[191\] vssd1 vssd1 vccd1 vccd1 net2087 sky130_fd_sc_hd__dlygate4sd3_1
Xhold756 final_design.cpu.reg_window\[922\] vssd1 vssd1 vccd1 vccd1 net2098 sky130_fd_sc_hd__dlygate4sd3_1
Xhold767 final_design.cpu.reg_window\[913\] vssd1 vssd1 vccd1 vccd1 net2109 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07946__A2 _02894_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold778 final_design.cpu.reg_window\[388\] vssd1 vssd1 vccd1 vccd1 net2120 sky130_fd_sc_hd__dlygate4sd3_1
X_09973_ net484 _04891_ _04341_ vssd1 vssd1 vccd1 vccd1 _04892_ sky130_fd_sc_hd__a21o_1
XFILLER_0_60_1239 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold789 final_design.cpu.reg_window\[92\] vssd1 vssd1 vccd1 vccd1 net2131 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09148__A1 _04066_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08924_ _02507_ _03864_ _03866_ net257 vssd1 vssd1 vccd1 vccd1 _03867_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout1011_A _05166_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12152__A0 net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09699__A2 net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1109_A net1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08855_ _03783_ _03805_ final_design.CPU_instr_adr\[31\] net1038 vssd1 vssd1 vccd1
+ vccd1 _00242_ sky130_fd_sc_hd__o2bb2a_1
XPHY_EDGE_ROW_24_Left_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout471_A _03485_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout569_A net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07806_ final_design.cpu.reg_window\[729\] final_design.cpu.reg_window\[761\] net850
+ vssd1 vssd1 vccd1 vccd1 _02757_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_2_Right_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08786_ _03734_ _03736_ _03686_ vssd1 vssd1 vccd1 vccd1 _03737_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_19_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11258__A2 net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07737_ final_design.cpu.reg_window\[794\] final_design.cpu.reg_window\[826\] net863
+ vssd1 vssd1 vccd1 vccd1 _02688_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout736_A _01490_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout357_X net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_64_clk clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_64_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_7_1821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10466__B1 net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07668_ final_design.cpu.reg_window\[222\] final_design.cpu.reg_window\[254\] net853
+ vssd1 vssd1 vccd1 vccd1 _02619_ sky130_fd_sc_hd__mux2_1
XANTENNA__07331__B1 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09407_ net89 _04195_ vssd1 vssd1 vccd1 vccd1 _04326_ sky130_fd_sc_hd__xor2_2
XANTENNA__13700__CLK clknet_leaf_54_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06619_ net741 _01497_ net665 _01569_ vssd1 vssd1 vccd1 vccd1 _01570_ sky130_fd_sc_hd__a211o_4
XFILLER_0_3_1729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout524_X net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07599_ final_design.cpu.reg_window\[285\] final_design.cpu.reg_window\[317\] net871
+ vssd1 vssd1 vccd1 vccd1 _02550_ sky130_fd_sc_hd__mux2_1
XANTENNA__11304__A net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09338_ net614 net525 _03523_ _01453_ vssd1 vssd1 vccd1 vccd1 _04257_ sky130_fd_sc_hd__a211o_1
XPHY_EDGE_ROW_33_Left_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_1431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11966__B1 net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09269_ net76 net77 _04187_ vssd1 vssd1 vccd1 vccd1 _04188_ sky130_fd_sc_hd__or3_1
XANTENNA__10604__A_N _04961_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13850__CLK clknet_leaf_58_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11300_ net650 net201 vssd1 vssd1 vccd1 vccd1 _05997_ sky130_fd_sc_hd__and2_1
X_12280_ net572 _06210_ net508 net371 net1740 vssd1 vssd1 vccd1 vccd1 _00995_ sky130_fd_sc_hd__a32o_1
XANTENNA__11718__B1 net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11231_ net560 net420 _05935_ net314 net1689 vssd1 vssd1 vccd1 vccd1 _00285_ sky130_fd_sc_hd__a32o_1
XANTENNA__09482__S1 net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11162_ _04879_ net651 net588 _05874_ vssd1 vssd1 vccd1 vccd1 _05875_ sky130_fd_sc_hd__o211a_1
XANTENNA__13407__RESET_B net1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09139__A1 net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10113_ net1051 _05023_ _05003_ vssd1 vssd1 vccd1 vccd1 _05025_ sky130_fd_sc_hd__o21ai_1
X_11093_ _05813_ _05814_ vssd1 vssd1 vccd1 vccd1 _05815_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_42_Left_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input32_A DAT_I[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10044_ _04249_ _04252_ _04289_ vssd1 vssd1 vccd1 vccd1 _04963_ sky130_fd_sc_hd__a21boi_1
XANTENNA__11693__B net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold50 final_design.cpu.reg_window\[0\] vssd1 vssd1 vccd1 vccd1 net1392 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13230__CLK clknet_leaf_43_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold61 final_design.reqhand.instruction\[17\] vssd1 vssd1 vccd1 vccd1 net1403 sky130_fd_sc_hd__dlygate4sd3_1
Xhold72 final_design.VGA_data_control.data_to_VGA\[10\] vssd1 vssd1 vccd1 vccd1 net1414
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold83 net108 vssd1 vssd1 vccd1 vccd1 net1425 sky130_fd_sc_hd__dlygate4sd3_1
Xhold94 net160 vssd1 vssd1 vccd1 vccd1 net1436 sky130_fd_sc_hd__dlygate4sd3_1
X_13803_ clknet_leaf_53_clk _01034_ net1185 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[791\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12446__A1 net207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11995_ _06197_ net281 net400 net2021 vssd1 vssd1 vccd1 vccd1 _00726_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_55_clk clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_55_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__11913__S net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09311__A1 _04222_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13734_ clknet_leaf_50_clk _00965_ net1173 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[722\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07899__A net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10946_ _04918_ net252 vssd1 vssd1 vccd1 vccd1 _05674_ sky130_fd_sc_hd__nor2_1
XFILLER_0_42_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_52_clk_X clknet_leaf_52_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13380__CLK clknet_leaf_52_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13665_ clknet_leaf_47_clk _00896_ net1199 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[653\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_32_1831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10472__A3 net250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10877_ _04598_ net252 vssd1 vssd1 vccd1 vccd1 _05608_ sky130_fd_sc_hd__nor2_1
XFILLER_0_32_1842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_51_Left_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_45_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12948__CLK clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11214__A net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12616_ net2259 net2267 _05080_ vssd1 vssd1 vccd1 vccd1 _01309_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_41_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13596_ clknet_leaf_3_clk _00827_ net1064 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[584\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_41_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_1905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_906 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12547_ _06210_ net351 net325 net2198 vssd1 vssd1 vccd1 vccd1 _01251_ sky130_fd_sc_hd__a22o_1
XANTENNA__09178__X _04097_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07838__S net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12478_ _06138_ net353 net332 net2264 vssd1 vssd1 vccd1 vccd1 _01184_ sky130_fd_sc_hd__a22o_1
XANTENNA__06742__S net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_3 _04589_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14217_ net1275 vssd1 vssd1 vccd1 vccd1 gpio_oeb[29] sky130_fd_sc_hd__buf_2
X_11429_ net1695 net199 net311 vssd1 vssd1 vccd1 vccd1 _00326_ sky130_fd_sc_hd__mux2_1
XANTENNA__09378__B2 net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_1695 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_39_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14148_ clknet_leaf_19_clk _01322_ net1112 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.data_to_VGA\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13148__RESET_B net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_60_Left_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06970_ final_design.cpu.reg_window\[144\] final_design.cpu.reg_window\[176\] net926
+ vssd1 vssd1 vccd1 vccd1 _01921_ sky130_fd_sc_hd__mux2_1
X_14079_ clknet_leaf_19_clk _01276_ net1111 vssd1 vssd1 vccd1 vccd1 final_design.reqhand.instruction\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12134__A0 net240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1070 net1072 vssd1 vssd1 vccd1 vccd1 net1070 sky130_fd_sc_hd__clkbuf_4
Xfanout1081 net1085 vssd1 vssd1 vccd1 vccd1 net1081 sky130_fd_sc_hd__clkbuf_4
X_08640_ _02932_ _02933_ _03586_ _03588_ vssd1 vssd1 vccd1 vccd1 _03591_ sky130_fd_sc_hd__o22a_1
Xfanout1092 net1093 vssd1 vssd1 vccd1 vccd1 net1092 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_59_1466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_1_239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08571_ _03520_ _03521_ vssd1 vssd1 vccd1 vccd1 _03522_ sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_46_clk clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_46_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_72_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11823__S net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07522_ _01631_ _02471_ _01600_ vssd1 vssd1 vccd1 vccd1 _02473_ sky130_fd_sc_hd__a21bo_1
XANTENNA__09360__Y _04279_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10999__A1 _04042_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10999__B2 _04040_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07453_ final_design.cpu.reg_window\[128\] final_design.cpu.reg_window\[160\] net895
+ vssd1 vssd1 vccd1 vccd1 _02404_ sky130_fd_sc_hd__mux2_1
XANTENNA__11660__A2 net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06404_ final_design.CPU_instr_adr\[27\] vssd1 vssd1 vccd1 vccd1 _01359_ sky130_fd_sc_hd__inv_2
XANTENNA__11124__A net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13873__CLK clknet_leaf_34_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07384_ final_design.cpu.reg_window\[450\] final_design.cpu.reg_window\[482\] net918
+ vssd1 vssd1 vccd1 vccd1 _02335_ sky130_fd_sc_hd__mux2_1
XANTENNA__11948__B1 net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09123_ net995 _01414_ vssd1 vssd1 vccd1 vccd1 _04042_ sky130_fd_sc_hd__nor2_8
XFILLER_0_33_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08704__Y _03655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout317_A _05851_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1059_A net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09054_ _03980_ _03982_ final_design.CPU_instr_adr\[9\] net1037 vssd1 vssd1 vccd1
+ vccd1 _00220_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__13103__CLK clknet_leaf_43_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08005_ final_design.cpu.reg_window\[656\] final_design.cpu.reg_window\[688\] net843
+ vssd1 vssd1 vccd1 vccd1 _02956_ sky130_fd_sc_hd__mux2_1
XANTENNA__11130__Y _05845_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold520 final_design.cpu.reg_window\[799\] vssd1 vssd1 vccd1 vccd1 net1862 sky130_fd_sc_hd__dlygate4sd3_1
Xhold531 final_design.cpu.reg_window\[980\] vssd1 vssd1 vccd1 vccd1 net1873 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1226_A net1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold542 final_design.cpu.reg_window\[200\] vssd1 vssd1 vccd1 vccd1 net1884 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold553 final_design.cpu.reg_window\[190\] vssd1 vssd1 vccd1 vccd1 net1895 sky130_fd_sc_hd__dlygate4sd3_1
Xhold564 final_design.cpu.reg_window\[768\] vssd1 vssd1 vccd1 vccd1 net1906 sky130_fd_sc_hd__dlygate4sd3_1
Xhold575 final_design.cpu.reg_window\[607\] vssd1 vssd1 vccd1 vccd1 net1917 sky130_fd_sc_hd__dlygate4sd3_1
Xhold586 final_design.cpu.reg_window\[507\] vssd1 vssd1 vccd1 vccd1 net1928 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_55_2080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold597 final_design.cpu.reg_window\[440\] vssd1 vssd1 vccd1 vccd1 net1939 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout686_A net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_2091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11794__A net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13253__CLK clknet_leaf_49_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09956_ _03488_ _03555_ _03556_ _04124_ vssd1 vssd1 vccd1 vccd1 _04875_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_70_2589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08907_ final_design.CPU_instr_adr\[24\] _03797_ final_design.CPU_instr_adr\[25\]
+ vssd1 vssd1 vccd1 vccd1 _03852_ sky130_fd_sc_hd__a21oi_1
X_09887_ net725 _04805_ net79 vssd1 vssd1 vccd1 vccd1 _04806_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout853_A net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout474_X net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08838_ final_design.CPU_instr_adr\[11\] _03788_ vssd1 vssd1 vccd1 vccd1 _03789_
+ sky130_fd_sc_hd__and2_1
XANTENNA__07778__S1 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout641_X net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08769_ _03710_ _03719_ _03709_ vssd1 vssd1 vccd1 vccd1 _03720_ sky130_fd_sc_hd__a21o_1
Xclkbuf_leaf_37_clk clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_37_clk sky130_fd_sc_hd__clkbuf_8
X_10800_ final_design.CPU_instr_adr\[17\] _05534_ net1055 vssd1 vssd1 vccd1 vccd1
+ _05535_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_836 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11780_ net646 net555 net221 vssd1 vssd1 vccd1 vccd1 _06231_ sky130_fd_sc_hd__and3_1
X_10731_ _05464_ _05468_ vssd1 vssd1 vccd1 vccd1 _05469_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout906_X net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11034__A _04421_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13450_ clknet_leaf_60_clk _00681_ net1143 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[438\]
+ sky130_fd_sc_hd__dfrtp_1
X_10662_ _05347_ _05385_ _05403_ vssd1 vssd1 vccd1 vccd1 _05404_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_12_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11939__B1 net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12401_ _06099_ net346 net338 net1987 vssd1 vssd1 vccd1 vccd1 _01111_ sky130_fd_sc_hd__a22o_1
XFILLER_0_36_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07607__A1 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13381_ clknet_leaf_52_clk _00612_ net1182 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[369\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_36_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10593_ _05336_ _05337_ vssd1 vssd1 vccd1 vccd1 _05338_ sky130_fd_sc_hd__nor2_1
XANTENNA__12600__B2 final_design.data_from_mem\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12332_ net2380 net361 net349 _05865_ vssd1 vssd1 vccd1 vccd1 _01044_ sky130_fd_sc_hd__a22o_1
XFILLER_0_23_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12263_ net672 _06193_ _06262_ vssd1 vssd1 vccd1 vccd1 _06274_ sky130_fd_sc_hd__or3_4
XANTENNA__11167__A1 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14002_ clknet_leaf_44_clk _01233_ net1207 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[990\]
+ sky130_fd_sc_hd__dfrtp_1
X_11214_ net588 _05919_ _05920_ vssd1 vssd1 vccd1 vccd1 _05921_ sky130_fd_sc_hd__and3_1
XFILLER_0_62_1857 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12194_ net1742 net178 net382 vssd1 vssd1 vccd1 vccd1 _00913_ sky130_fd_sc_hd__mux2_1
XANTENNA__07466__S0 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11145_ net662 _04028_ net734 vssd1 vssd1 vccd1 vccd1 _05859_ sky130_fd_sc_hd__a21o_1
XFILLER_0_43_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09174__A net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input35_X net35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07218__S0 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11076_ _05757_ _05775_ _05792_ _05797_ vssd1 vssd1 vccd1 vccd1 _05798_ sky130_fd_sc_hd__o31ai_2
XANTENNA__13746__CLK clknet_leaf_39_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12667__B2 final_design.data_from_mem\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10027_ _02837_ net445 _04943_ _04945_ vssd1 vssd1 vccd1 vccd1 _04946_ sky130_fd_sc_hd__o211a_1
XANTENNA__12419__A1 _06017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_28_clk clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_28_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_47_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13896__CLK clknet_leaf_41_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_1915 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11978_ _06180_ net292 net406 net1843 vssd1 vssd1 vccd1 vccd1 _00711_ sky130_fd_sc_hd__a22o_1
XFILLER_0_53_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10929_ net1055 _05656_ _05657_ vssd1 vssd1 vccd1 vccd1 _05658_ sky130_fd_sc_hd__a21oi_1
X_13717_ clknet_leaf_58_clk _00948_ net1133 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[705\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_1347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11642__A2 net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07141__B net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07941__S1 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_32_clk_A clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13126__CLK clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13648_ clknet_leaf_36_clk _00879_ net1236 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[636\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12198__A3 net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13579_ clknet_leaf_52_clk _00810_ net1183 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[567\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10602__B1 net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11598__B net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10387__B1_N _05174_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14239__1293 vssd1 vssd1 vccd1 vccd1 _14239__1293/HI net1293 sky130_fd_sc_hd__conb_1
XANTENNA_clkbuf_leaf_47_clk_A clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13276__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1913 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11158__A1 net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12355__B1 net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10007__B net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11818__S net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout307 _06095_ vssd1 vssd1 vccd1 vccd1 net307 sky130_fd_sc_hd__buf_4
X_09810_ _03262_ _04087_ vssd1 vssd1 vccd1 vccd1 _04729_ sky130_fd_sc_hd__nand2_1
Xfanout318 _04117_ vssd1 vssd1 vccd1 vccd1 net318 sky130_fd_sc_hd__clkbuf_4
Xfanout329 _06284_ vssd1 vssd1 vccd1 vccd1 net329 sky130_fd_sc_hd__clkbuf_8
XANTENNA__06585__A1 net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09741_ _03230_ _04495_ _03571_ _03198_ vssd1 vssd1 vccd1 vccd1 _04660_ sky130_fd_sc_hd__a211o_1
X_06953_ final_design.cpu.reg_window\[593\] final_design.cpu.reg_window\[625\] net925
+ vssd1 vssd1 vccd1 vccd1 _01904_ sky130_fd_sc_hd__mux2_1
XANTENNA__12964__RESET_B net1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09672_ _02803_ _03034_ vssd1 vssd1 vccd1 vccd1 _04591_ sky130_fd_sc_hd__nand2_1
XANTENNA__07316__B _01659_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10023__A net68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06884_ final_design.cpu.reg_window\[147\] final_design.cpu.reg_window\[179\] net911
+ vssd1 vssd1 vccd1 vccd1 _01835_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08623_ _02185_ _03289_ vssd1 vssd1 vccd1 vccd1 _03574_ sky130_fd_sc_hd__nand2_1
XANTENNA__10958__A net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_19_clk clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_19_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__11881__A2 net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11406__X _06090_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08554_ _03501_ _03502_ _03503_ _03504_ net680 net700 vssd1 vssd1 vccd1 vccd1 _03505_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__06647__S net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11780__C net221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07505_ _01941_ _02455_ _01940_ vssd1 vssd1 vccd1 vccd1 _02456_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_4_1813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08485_ _03432_ _03433_ _03434_ _03435_ net677 net701 vssd1 vssd1 vccd1 vccd1 _03436_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_63_2360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout434_A net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_2371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1176_A net1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10396__C net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1857 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07436_ _02383_ _02384_ _02385_ _02386_ net769 net782 vssd1 vssd1 vccd1 vccd1 _02387_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__14051__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07367_ net751 _02317_ vssd1 vssd1 vccd1 vccd1 _02318_ sky130_fd_sc_hd__or2_1
XANTENNA__12384__S net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout601_A _02514_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07986__B net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13619__CLK clknet_leaf_40_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12594__B1 net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09106_ net1018 _04027_ net1037 vssd1 vssd1 vccd1 vccd1 _00213_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06499__S1 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07298_ final_design.cpu.reg_window\[325\] final_design.cpu.reg_window\[357\] net921
+ vssd1 vssd1 vccd1 vccd1 _02249_ sky130_fd_sc_hd__mux2_1
X_09037_ final_design.CPU_instr_adr\[9\] _03787_ final_design.CPU_instr_adr\[10\]
+ vssd1 vssd1 vccd1 vccd1 _03967_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_57_2142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_2153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_2787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12775__6 clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 net1316 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_57_2164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_2798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12346__B1 net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_2006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_2017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08014__A1 _01908_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_2028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold350 final_design.cpu.reg_window\[221\] vssd1 vssd1 vccd1 vccd1 net1692 sky130_fd_sc_hd__dlygate4sd3_1
Xhold361 final_design.cpu.reg_window\[756\] vssd1 vssd1 vccd1 vccd1 net1703 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13769__CLK clknet_leaf_36_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout591_X net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout689_X net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold372 final_design.cpu.reg_window\[846\] vssd1 vssd1 vccd1 vccd1 net1714 sky130_fd_sc_hd__dlygate4sd3_1
Xhold383 final_design.cpu.reg_window\[855\] vssd1 vssd1 vccd1 vccd1 net1725 sky130_fd_sc_hd__dlygate4sd3_1
Xhold394 final_design.cpu.reg_window\[699\] vssd1 vssd1 vccd1 vccd1 net1736 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10372__A2 net1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout830 net834 vssd1 vssd1 vccd1 vccd1 net830 sky130_fd_sc_hd__clkbuf_4
Xfanout841 net842 vssd1 vssd1 vccd1 vccd1 net841 sky130_fd_sc_hd__buf_2
XANTENNA__08970__C1 net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout852 net873 vssd1 vssd1 vccd1 vccd1 net852 sky130_fd_sc_hd__buf_2
X_09939_ net263 _04854_ _04857_ vssd1 vssd1 vccd1 vccd1 _04858_ sky130_fd_sc_hd__and3_1
XANTENNA__12649__B2 final_design.data_from_mem\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout863 net864 vssd1 vssd1 vccd1 vccd1 net863 sky130_fd_sc_hd__clkbuf_4
Xfanout874 net876 vssd1 vssd1 vccd1 vccd1 net874 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_77_1330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout885 net886 vssd1 vssd1 vccd1 vccd1 net885 sky130_fd_sc_hd__clkbuf_8
X_12950_ clknet_leaf_29_clk _00188_ net1194 vssd1 vssd1 vccd1 vccd1 net107 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_5_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout896 net899 vssd1 vssd1 vccd1 vccd1 net896 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_5_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1050 final_design.cpu.reg_window\[122\] vssd1 vssd1 vccd1 vccd1 net2392 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11321__A1 _01788_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11321__B2 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11901_ net223 net2046 net274 vssd1 vssd1 vccd1 vccd1 _00643_ sky130_fd_sc_hd__mux2_1
Xhold1061 final_design.cpu.reg_window\[40\] vssd1 vssd1 vccd1 vccd1 net2403 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_73_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1072 final_design.cpu.reg_window\[870\] vssd1 vssd1 vccd1 vccd1 net2414 sky130_fd_sc_hd__dlygate4sd3_1
X_12881_ clknet_leaf_17_clk _00119_ net1114 vssd1 vssd1 vccd1 vccd1 final_design.data_from_mem\[15\]
+ sky130_fd_sc_hd__dfrtp_4
Xhold1083 final_design.cpu.reg_window\[368\] vssd1 vssd1 vccd1 vccd1 net2425 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1094 final_design.cpu.reg_window\[909\] vssd1 vssd1 vccd1 vccd1 net2436 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11463__S net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11832_ _06017_ net2323 net266 vssd1 vssd1 vccd1 vccd1 _00584_ sky130_fd_sc_hd__mux2_1
XANTENNA__13149__CLK clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07242__A net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08176__S1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11763_ net185 net2019 net419 vssd1 vssd1 vccd1 vccd1 _00526_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11624__A2 net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10714_ final_design.CPU_instr_adr\[13\] _03951_ net1058 vssd1 vssd1 vccd1 vccd1
+ _05453_ sky130_fd_sc_hd__mux2_1
XANTENNA__07923__S1 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13502_ clknet_leaf_13_clk _00733_ net1099 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[490\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11694_ net429 net568 _06205_ net295 net1696 vssd1 vssd1 vccd1 vccd1 _00478_ sky130_fd_sc_hd__a32o_1
X_13433_ clknet_leaf_56_clk _00664_ net1147 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[421\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11699__A net207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10645_ net1002 _05384_ _05387_ net1031 net1360 vssd1 vssd1 vccd1 vccd1 _00182_ sky130_fd_sc_hd__a32o_1
XFILLER_0_67_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13299__CLK clknet_leaf_40_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12585__B1 net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13364_ clknet_leaf_9_clk _00595_ net1151 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[352\]
+ sky130_fd_sc_hd__dfrtp_1
X_10576_ net958 _05319_ _05321_ net955 vssd1 vssd1 vccd1 vccd1 _05322_ sky130_fd_sc_hd__o22a_1
XANTENNA__09450__B1 net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12315_ net1941 net202 net366 vssd1 vssd1 vccd1 vccd1 _01029_ sky130_fd_sc_hd__mux2_1
X_13295_ clknet_leaf_41_clk _00526_ net1224 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[283\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12337__B1 net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12246_ final_design.cpu.reg_window\[720\] net375 vssd1 vssd1 vccd1 vccd1 _06273_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_82_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_1627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_1676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08100__S1 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09175__Y _04094_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12177_ net2139 net210 net383 vssd1 vssd1 vccd1 vccd1 _00896_ sky130_fd_sc_hd__mux2_1
XANTENNA__09616__B _04094_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10363__A2 net1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11128_ _02295_ _05839_ vssd1 vssd1 vccd1 vccd1 _05843_ sky130_fd_sc_hd__nor2_8
XFILLER_0_21_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08308__A2 _03257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11059_ _05780_ _05781_ _05761_ vssd1 vssd1 vccd1 vccd1 _05782_ sky130_fd_sc_hd__o21ai_1
XANTENNA__08947__S net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11312__A1 final_design.data_from_mem\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09351__B _04094_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1761 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14074__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10823__B1 net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08270_ final_design.cpu.reg_window\[522\] final_design.cpu.reg_window\[554\] net814
+ vssd1 vssd1 vccd1 vccd1 _03221_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07221_ final_design.cpu.reg_window\[712\] final_design.cpu.reg_window\[744\] net889
+ vssd1 vssd1 vccd1 vccd1 _02172_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07152_ final_design.cpu.reg_window\[394\] final_design.cpu.reg_window\[426\] net898
+ vssd1 vssd1 vccd1 vccd1 _02103_ sky130_fd_sc_hd__mux2_1
XANTENNA__07047__A2 net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13911__CLK clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07083_ final_design.cpu.reg_window\[332\] final_design.cpu.reg_window\[364\] net907
+ vssd1 vssd1 vccd1 vccd1 _02034_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_8_clk clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_8_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_80_1721 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_2640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_1885 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09744__A1 net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10354__A2 net1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11551__A1 net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07985_ _02935_ vssd1 vssd1 vccd1 vccd1 _02936_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout384_A net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09724_ _04641_ _04642_ net477 vssd1 vssd1 vccd1 vccd1 _04643_ sky130_fd_sc_hd__mux2_1
X_06936_ final_design.cpu.reg_window\[337\] final_design.cpu.reg_window\[369\] net928
+ vssd1 vssd1 vccd1 vccd1 _01887_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_2_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11303__A1 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12500__B1 net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1514 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09655_ _04571_ _04573_ vssd1 vssd1 vccd1 vccd1 _04574_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_65_2411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12379__S net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06867_ _01816_ _01817_ vssd1 vssd1 vccd1 vccd1 _01818_ sky130_fd_sc_hd__nand2_4
XANTENNA__11854__A2 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout551_A _01750_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_2422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_2433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout649_A net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08606_ _03555_ _03556_ _03488_ vssd1 vssd1 vccd1 vccd1 _03557_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11136__X _05851_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_3_2_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_3_2_0_clk sky130_fd_sc_hd__clkbuf_8
X_09586_ _03070_ _03101_ _04504_ _04137_ vssd1 vssd1 vccd1 vccd1 _04505_ sky130_fd_sc_hd__a31o_1
X_06798_ net752 _01748_ net883 vssd1 vssd1 vccd1 vccd1 _01749_ sky130_fd_sc_hd__o21ai_1
X_08537_ _03486_ _03487_ vssd1 vssd1 vccd1 vccd1 _03488_ sky130_fd_sc_hd__nor2_2
XANTENNA__10200__B net35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout437_X net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout816_A net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13441__CLK clknet_leaf_48_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09688__S net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07905__S1 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07997__A net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08468_ net609 _03415_ _03416_ vssd1 vssd1 vccd1 vccd1 _03419_ sky130_fd_sc_hd__a21o_2
XFILLER_0_33_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07419_ final_design.cpu.reg_window\[65\] final_design.cpu.reg_window\[97\] net916
+ vssd1 vssd1 vccd1 vccd1 _02370_ sky130_fd_sc_hd__mux2_1
X_08399_ _03346_ _03347_ _03348_ _03349_ net677 net691 vssd1 vssd1 vccd1 vccd1 _03350_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_59_2215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10430_ net1435 net1028 _05198_ net245 vssd1 vssd1 vccd1 vccd1 _00156_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_59_2226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_2237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13591__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12127__B net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10361_ net3 net1025 net1008 final_design.data_from_mem\[10\] vssd1 vssd1 vccd1 vccd1
+ _00114_ sky130_fd_sc_hd__a22o_1
X_12100_ net1923 net225 net391 vssd1 vssd1 vccd1 vccd1 _00824_ sky130_fd_sc_hd__mux2_1
XANTENNA__09717__A net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13080_ clknet_leaf_62_clk _00311_ net1120 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[68\]
+ sky130_fd_sc_hd__dfrtp_1
X_10292_ _05144_ _05145_ _01384_ vssd1 vssd1 vccd1 vccd1 _05146_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout973_X net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12031_ net2163 net240 net396 vssd1 vssd1 vccd1 vccd1 _00759_ sky130_fd_sc_hd__mux2_1
Xhold180 final_design.VGA_data_control.ready_data\[14\] vssd1 vssd1 vccd1 vccd1 net1522
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold191 final_design.reqhand.current_client\[0\] vssd1 vssd1 vccd1 vccd1 net1533
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10345__A2 net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout660 _02512_ vssd1 vssd1 vccd1 vccd1 net660 sky130_fd_sc_hd__clkbuf_4
Xfanout671 net672 vssd1 vssd1 vccd1 vccd1 net671 sky130_fd_sc_hd__buf_2
Xfanout682 net689 vssd1 vssd1 vccd1 vccd1 net682 sky130_fd_sc_hd__clkbuf_8
Xfanout693 net695 vssd1 vssd1 vccd1 vccd1 net693 sky130_fd_sc_hd__buf_4
X_13982_ clknet_leaf_13_clk _01213_ net1099 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[970\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14097__CLK clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12933_ clknet_leaf_50_clk _00171_ net1172 vssd1 vssd1 vccd1 vccd1 net157 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14238__1292 vssd1 vssd1 vccd1 vccd1 _14238__1292/HI net1292 sky130_fd_sc_hd__conb_1
XFILLER_0_70_1901 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12864_ clknet_leaf_19_clk _00102_ net1157 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.ready_data\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_11815_ net239 net2207 net264 vssd1 vssd1 vccd1 vccd1 _00567_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11746_ net217 net2347 net416 vssd1 vssd1 vccd1 vccd1 _00509_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13934__CLK clknet_leaf_45_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11677_ net226 net627 vssd1 vssd1 vccd1 vccd1 _06197_ sky130_fd_sc_hd__and2_1
XFILLER_0_37_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12558__B1 net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11222__A net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10628_ _05351_ _05370_ vssd1 vssd1 vccd1 vccd1 _05371_ sky130_fd_sc_hd__nand2_1
X_13416_ clknet_leaf_35_clk _00647_ net1241 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[404\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12022__A2 net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13347_ clknet_leaf_1_clk _00578_ net1074 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[335\]
+ sky130_fd_sc_hd__dfrtp_1
X_10559_ _05268_ _05305_ vssd1 vssd1 vccd1 vccd1 _05306_ sky130_fd_sc_hd__and2_1
XFILLER_0_52_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11781__B2 net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13278_ clknet_leaf_9_clk _00509_ net1103 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[266\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09726__A1 _01626_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12229_ net671 _06158_ _06262_ vssd1 vssd1 vccd1 vccd1 _06272_ sky130_fd_sc_hd__or3_4
XFILLER_0_75_12 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13314__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07147__A _02097_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07832__S0 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07770_ final_design.cpu.reg_window\[792\] final_design.cpu.reg_window\[824\] net864
+ vssd1 vssd1 vccd1 vccd1 _02721_ sky130_fd_sc_hd__mux2_1
X_06721_ final_design.cpu.reg_window\[408\] final_design.cpu.reg_window\[440\] net944
+ vssd1 vssd1 vccd1 vccd1 _01672_ sky130_fd_sc_hd__mux2_1
XANTENNA__11297__B1 net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13464__CLK clknet_leaf_62_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09440_ _02769_ _03597_ vssd1 vssd1 vccd1 vccd1 _04359_ sky130_fd_sc_hd__nand2_1
X_06652_ final_design.cpu.reg_window\[282\] final_design.cpu.reg_window\[314\] net943
+ vssd1 vssd1 vccd1 vccd1 _01603_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09371_ _04286_ _04288_ vssd1 vssd1 vccd1 vccd1 _04290_ sky130_fd_sc_hd__or2_1
X_06583_ net761 _01533_ vssd1 vssd1 vccd1 vccd1 _01534_ sky130_fd_sc_hd__or2_1
XANTENNA__11831__S net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08322_ _03269_ _03270_ _03271_ _03272_ net675 net697 vssd1 vssd1 vccd1 vccd1 _03273_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_75_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1805 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08253_ final_design.cpu.reg_window\[394\] final_design.cpu.reg_window\[426\] net818
+ vssd1 vssd1 vccd1 vccd1 _03204_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08560__S1 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12549__B1 net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07204_ net881 _02148_ _02154_ _02141_ _02142_ vssd1 vssd1 vccd1 vccd1 _02155_ sky130_fd_sc_hd__a32oi_2
XFILLER_0_43_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12013__A2 net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08184_ _02000_ net599 vssd1 vssd1 vccd1 vccd1 _03135_ sky130_fd_sc_hd__nand2_1
XANTENNA__09414__B1 net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1805 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07135_ final_design.cpu.reg_window\[651\] final_design.cpu.reg_window\[683\] net909
+ vssd1 vssd1 vccd1 vccd1 _02086_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_73_2702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_1849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1139_A net1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07066_ final_design.cpu.reg_window\[717\] final_design.cpu.reg_window\[749\] net934
+ vssd1 vssd1 vccd1 vccd1 _02017_ sky130_fd_sc_hd__mux2_1
XANTENNA__07440__A2 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout599_A net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10035__X _04954_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07057__A net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout766_A net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout387_X net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07968_ final_design.cpu.reg_window\[913\] final_design.cpu.reg_window\[945\] net845
+ vssd1 vssd1 vccd1 vccd1 _02919_ sky130_fd_sc_hd__mux2_1
XANTENNA__13807__CLK clknet_leaf_42_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_2506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06919_ final_design.cpu.reg_window\[786\] final_design.cpu.reg_window\[818\] net925
+ vssd1 vssd1 vccd1 vccd1 _01870_ sky130_fd_sc_hd__mux2_1
X_09707_ _04124_ _04625_ _04624_ net263 vssd1 vssd1 vccd1 vccd1 _04626_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout554_X net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07899_ net721 _02849_ vssd1 vssd1 vccd1 vccd1 _02850_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout933_A net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09638_ _02995_ net440 vssd1 vssd1 vccd1 vccd1 _04557_ sky130_fd_sc_hd__nand2_1
XANTENNA__07900__B1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13957__CLK clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09569_ net319 _04487_ vssd1 vssd1 vccd1 vccd1 _04488_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout721_X net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11741__S net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11600_ net176 net636 vssd1 vssd1 vccd1 vccd1 _06156_ sky130_fd_sc_hd__and2_2
XFILLER_0_72_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12580_ _01395_ _04037_ vssd1 vssd1 vccd1 vccd1 _06295_ sky130_fd_sc_hd__nand2b_1
X_11531_ net1546 net184 net523 vssd1 vssd1 vccd1 vccd1 _00398_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12981__CLK clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14250_ net1304 vssd1 vssd1 vccd1 vccd1 gpio_out[28] sky130_fd_sc_hd__buf_2
XFILLER_0_11_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11462_ net219 net638 vssd1 vssd1 vccd1 vccd1 _06104_ sky130_fd_sc_hd__and2_1
XANTENNA__08208__A1 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1159 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13201_ clknet_leaf_33_clk _00432_ net1238 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[189\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11212__B1 _05916_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10413_ net1430 net1027 _05189_ net246 vssd1 vssd1 vccd1 vccd1 _00148_ sky130_fd_sc_hd__a22o_1
XFILLER_0_33_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14181_ clknet_leaf_21_clk _01355_ net1161 vssd1 vssd1 vccd1 vccd1 final_design.VGA_adr\[8\]
+ sky130_fd_sc_hd__dfrtp_4
X_11393_ final_design.data_from_mem\[30\] net235 net233 vssd1 vssd1 vccd1 vccd1 _06078_
+ sky130_fd_sc_hd__a21o_2
XFILLER_0_60_160 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_683 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13132_ clknet_leaf_46_clk _00363_ net1214 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[120\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input62_A mem_adr_start[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10344_ net1534 net1012 net989 final_design.data_from_mem\[29\] vssd1 vssd1 vccd1
+ vccd1 _00101_ sky130_fd_sc_hd__a22o_1
XANTENNA__13337__CLK clknet_leaf_55_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13063_ clknet_leaf_62_clk _00294_ net1119 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[51\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10275_ _05134_ _05135_ vssd1 vssd1 vccd1 vccd1 _00025_ sky130_fd_sc_hd__nor2_1
XFILLER_0_63_1793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11515__A1 net209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12790__21_A clknet_leaf_30_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12014_ _06216_ net283 net401 net2360 vssd1 vssd1 vccd1 vccd1 _00745_ sky130_fd_sc_hd__a22o_1
XANTENNA__09184__A2 _03550_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output149_A net149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11916__S net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13487__CLK clknet_leaf_42_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10820__S net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout490 _03453_ vssd1 vssd1 vccd1 vccd1 net490 sky130_fd_sc_hd__buf_2
XANTENNA__09182__A _04097_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09567__S0 net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13965_ clknet_leaf_48_clk _01196_ net1200 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[953\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_31_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12916_ clknet_leaf_50_clk _00154_ net1168 vssd1 vssd1 vccd1 vccd1 net138 sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkload8_A clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07042__S1 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12491__A2 net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13896_ clknet_leaf_41_clk _01127_ net1225 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[884\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09892__B1 net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12847_ clknet_leaf_18_clk _00085_ net1110 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.ready_data\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_17_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12798__29 clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 net1339 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_17_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_1737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11451__A0 net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08542__S1 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11729_ net180 net628 vssd1 vssd1 vccd1 vccd1 _06223_ sky130_fd_sc_hd__and2_1
XFILLER_0_9_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_25_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14112__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09086__A1_N net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xwire880 _01473_ vssd1 vssd1 vccd1 vccd1 net880 sky130_fd_sc_hd__clkbuf_1
Xhold905 final_design.cpu.reg_window\[797\] vssd1 vssd1 vccd1 vccd1 net2247 sky130_fd_sc_hd__dlygate4sd3_1
Xhold916 final_design.cpu.reg_window\[789\] vssd1 vssd1 vccd1 vccd1 net2258 sky130_fd_sc_hd__dlygate4sd3_1
Xhold927 final_design.cpu.reg_window\[871\] vssd1 vssd1 vccd1 vccd1 net2269 sky130_fd_sc_hd__dlygate4sd3_1
Xhold938 final_design.cpu.reg_window\[386\] vssd1 vssd1 vccd1 vccd1 net2280 sky130_fd_sc_hd__dlygate4sd3_1
Xhold949 final_design.cpu.reg_window\[1015\] vssd1 vssd1 vccd1 vccd1 net2291 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06856__S1 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08940_ final_design.CPU_instr_adr\[20\] _01823_ _03753_ vssd1 vssd1 vccd1 vccd1
+ _03881_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_0_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08871_ final_design.CPU_instr_adr\[29\] _03800_ vssd1 vssd1 vccd1 vccd1 _03820_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_42_1877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07805__S0 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11826__S net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07822_ _01788_ net606 vssd1 vssd1 vccd1 vccd1 _02773_ sky130_fd_sc_hd__nand2_1
XFILLER_0_19_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07281__S1 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12854__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07753_ _02701_ _02703_ vssd1 vssd1 vccd1 vccd1 _02704_ sky130_fd_sc_hd__nor2_1
XANTENNA__08200__S net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11809__A2 net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06704_ _01651_ _01652_ _01653_ _01654_ net772 net783 vssd1 vssd1 vccd1 vccd1 _01655_
+ sky130_fd_sc_hd__mux4_1
X_07684_ _02622_ _02623_ _02634_ net878 vssd1 vssd1 vccd1 vccd1 _02635_ sky130_fd_sc_hd__a22oi_4
XANTENNA__12482__A2 net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09423_ _03627_ _04341_ vssd1 vssd1 vccd1 vccd1 _04342_ sky130_fd_sc_hd__or2_4
XFILLER_0_48_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06635_ final_design.cpu.reg_window\[987\] final_design.cpu.reg_window\[1019\] net945
+ vssd1 vssd1 vccd1 vccd1 _01586_ sky130_fd_sc_hd__mux2_1
XANTENNA__11690__B1 net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1913 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout347_A net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09354_ net492 _04231_ _04261_ _04265_ _04272_ vssd1 vssd1 vccd1 vccd1 _04273_ sky130_fd_sc_hd__o311a_1
XANTENNA_fanout1089_A net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06566_ final_design.cpu.reg_window\[29\] final_design.cpu.reg_window\[61\] net950
+ vssd1 vssd1 vccd1 vccd1 _01517_ sky130_fd_sc_hd__mux2_1
X_08305_ net707 _03255_ net874 vssd1 vssd1 vccd1 vccd1 _03256_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_79_2900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07379__A2_N net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_2911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_1793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09285_ net527 net458 _04203_ net467 vssd1 vssd1 vccd1 vccd1 _04204_ sky130_fd_sc_hd__a211o_1
X_06497_ final_design.cpu.reg_window\[606\] final_design.cpu.reg_window\[638\] net931
+ vssd1 vssd1 vccd1 vccd1 _01448_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout514_A net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08236_ final_design.cpu.reg_window\[651\] final_design.cpu.reg_window\[683\] net826
+ vssd1 vssd1 vccd1 vccd1 _03187_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09938__A1 _04222_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08167_ final_design.cpu.reg_window\[847\] final_design.cpu.reg_window\[879\] net819
+ vssd1 vssd1 vccd1 vccd1 _03118_ sky130_fd_sc_hd__mux2_1
XANTENNA__12392__S net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout302_X net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07118_ final_design.cpu.reg_window\[267\] final_design.cpu.reg_window\[299\] net916
+ vssd1 vssd1 vccd1 vccd1 _02069_ sky130_fd_sc_hd__mux2_1
X_14237__1291 vssd1 vssd1 vccd1 vccd1 _14237__1291/HI net1291 sky130_fd_sc_hd__conb_1
X_08098_ final_design.cpu.reg_window\[204\] final_design.cpu.reg_window\[236\] net815
+ vssd1 vssd1 vccd1 vccd1 _03049_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout883_A _01437_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12786__17_A clknet_leaf_27_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07049_ net743 net667 net664 _01999_ _01821_ vssd1 vssd1 vccd1 vccd1 _02000_ sky130_fd_sc_hd__o221ai_4
XFILLER_0_80_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10060_ _04967_ _04969_ _04977_ _04978_ vssd1 vssd1 vccd1 vccd1 _04979_ sky130_fd_sc_hd__and4_1
XFILLER_0_21_1917 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07177__A1 _01505_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout769_X net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11736__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_1873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10962_ _05689_ vssd1 vssd1 vccd1 vccd1 _05690_ sky130_fd_sc_hd__inv_2
X_13750_ clknet_leaf_60_clk _00981_ net1137 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[738\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12473__A2 net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07024__S1 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1868 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12701_ final_design.VGA_data_control.v_count\[5\] _06339_ _06335_ vssd1 vssd1 vccd1
+ vccd1 _06342_ sky130_fd_sc_hd__o21ai_1
XANTENNA__09730__A net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10893_ _05606_ _05622_ vssd1 vssd1 vccd1 vccd1 _05624_ sky130_fd_sc_hd__or2_1
X_13681_ clknet_leaf_35_clk _00912_ net1240 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[669\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14135__CLK clknet_leaf_17_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12632_ _06303_ net1419 net980 vssd1 vssd1 vccd1 vccd1 _01318_ sky130_fd_sc_hd__mux2_1
XANTENNA__12225__A2 _06153_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12563_ net1052 _05078_ _05066_ vssd1 vssd1 vccd1 vccd1 _06286_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_25_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11514_ net1715 net212 net521 vssd1 vssd1 vccd1 vccd1 _00383_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_43_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12494_ _06154_ net358 net332 net2308 vssd1 vssd1 vccd1 vccd1 _01200_ sky130_fd_sc_hd__a22o_1
XFILLER_0_41_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14233_ net1287 vssd1 vssd1 vccd1 vccd1 gpio_out[11] sky130_fd_sc_hd__buf_2
XFILLER_0_80_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11445_ net232 net2371 net306 vssd1 vssd1 vccd1 vccd1 _00339_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10539__A2 net1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07396__S net913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14164_ clknet_leaf_17_clk _01338_ net1109 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.data_to_VGA\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_1708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11376_ net733 _03829_ _06062_ vssd1 vssd1 vccd1 vccd1 _06063_ sky130_fd_sc_hd__o21a_1
X_10327_ net1514 net1010 net987 final_design.data_from_mem\[12\] vssd1 vssd1 vccd1
+ vccd1 _00084_ sky130_fd_sc_hd__a22o_1
X_13115_ clknet_leaf_66_clk _00346_ net1063 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[103\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14095_ clknet_leaf_9_clk _01292_ net1151 vssd1 vssd1 vccd1 vccd1 final_design.reqhand.instruction\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_13046_ clknet_leaf_61_clk _00277_ net1139 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[34\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_37_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09157__A2 net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12877__CLK clknet_leaf_17_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10258_ final_design.uart.BAUD_counter\[21\] _05123_ net797 vssd1 vssd1 vccd1 vccd1
+ _05125_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_37_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1230 net1232 vssd1 vssd1 vccd1 vccd1 net1230 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_33_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1241 net1244 vssd1 vssd1 vccd1 vccd1 net1241 sky130_fd_sc_hd__buf_2
XANTENNA__12331__A net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10189_ _05078_ vssd1 vssd1 vccd1 vccd1 _05079_ sky130_fd_sc_hd__inv_2
X_13948_ clknet_leaf_3_clk _01179_ net1079 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[936\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09865__B1 net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1214 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11672__A0 net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06679__B1 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10475__B2 final_design.CPU_instr_adr\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13879_ clknet_leaf_58_clk _01110_ net1132 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[867\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_27_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06420_ final_design.data_from_mem\[2\] vssd1 vssd1 vccd1 vccd1 _01375_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_27_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09617__B1 _04117_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1572 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_904 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12989__RESET_B net1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13502__CLK clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09070_ _03655_ _03995_ _03996_ _03993_ net1037 vssd1 vssd1 vccd1 vccd1 _03997_ sky130_fd_sc_hd__o221a_1
XFILLER_0_66_1619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08021_ net710 _02971_ vssd1 vssd1 vccd1 vccd1 _02972_ sky130_fd_sc_hd__nor2_1
XFILLER_0_4_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13652__CLK clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold702 final_design.cpu.reg_window\[441\] vssd1 vssd1 vccd1 vccd1 net2044 sky130_fd_sc_hd__dlygate4sd3_1
Xhold713 final_design.cpu.reg_window\[279\] vssd1 vssd1 vccd1 vccd1 net2055 sky130_fd_sc_hd__dlygate4sd3_1
Xhold724 final_design.cpu.reg_window\[165\] vssd1 vssd1 vccd1 vccd1 net2066 sky130_fd_sc_hd__dlygate4sd3_1
Xhold735 final_design.cpu.reg_window\[409\] vssd1 vssd1 vccd1 vccd1 net2077 sky130_fd_sc_hd__dlygate4sd3_1
Xhold746 final_design.cpu.reg_window\[994\] vssd1 vssd1 vccd1 vccd1 net2088 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkload34_A clknet_leaf_43_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold757 final_design.cpu.reg_window\[959\] vssd1 vssd1 vccd1 vccd1 net2099 sky130_fd_sc_hd__dlygate4sd3_1
Xhold768 final_design.cpu.reg_window\[898\] vssd1 vssd1 vccd1 vccd1 net2110 sky130_fd_sc_hd__dlygate4sd3_1
Xhold779 final_design.cpu.reg_window\[211\] vssd1 vssd1 vccd1 vccd1 net2121 sky130_fd_sc_hd__dlygate4sd3_1
X_09972_ _04663_ _04815_ net471 vssd1 vssd1 vccd1 vccd1 _04891_ sky130_fd_sc_hd__mux2_1
XANTENNA__14008__CLK clknet_leaf_63_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08923_ net621 _03865_ vssd1 vssd1 vccd1 vccd1 _03866_ sky130_fd_sc_hd__nor2_1
XFILLER_0_41_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout297_A _06194_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09699__A3 net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11409__X _06092_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10313__X _05166_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08854_ net256 _03804_ net1014 vssd1 vssd1 vccd1 vccd1 _03805_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout1004_A _05173_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07805_ _02752_ _02753_ _02754_ _02755_ net684 net703 vssd1 vssd1 vccd1 vccd1 _02756_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__11128__Y _05843_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08785_ _01365_ _02063_ _03685_ vssd1 vssd1 vccd1 vccd1 _03736_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout464_A _03519_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13032__CLK clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14158__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07736_ final_design.cpu.reg_window\[858\] final_design.cpu.reg_window\[890\] net863
+ vssd1 vssd1 vccd1 vccd1 _02687_ sky130_fd_sc_hd__mux2_1
XANTENNA__11258__A3 _05959_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09550__A _04072_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10466__A1 net68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10466__B2 final_design.CPU_instr_adr\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1833 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12387__S net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07667_ final_design.cpu.reg_window\[30\] final_design.cpu.reg_window\[62\] net856
+ vssd1 vssd1 vccd1 vccd1 _02618_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout252_X net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout631_A _06157_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07331__A1 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout729_A net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09406_ _01493_ _04324_ vssd1 vssd1 vccd1 vccd1 _04325_ sky130_fd_sc_hd__nor2_1
XFILLER_0_1_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06618_ net744 _01568_ vssd1 vssd1 vccd1 vccd1 _01569_ sky130_fd_sc_hd__and2_1
X_07598_ final_design.cpu.reg_window\[349\] final_design.cpu.reg_window\[381\] net871
+ vssd1 vssd1 vccd1 vccd1 _02549_ sky130_fd_sc_hd__mux2_1
XANTENNA__07882__A2 _02830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13182__CLK clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1180 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09337_ _03602_ _04254_ _02673_ vssd1 vssd1 vccd1 vccd1 _04256_ sky130_fd_sc_hd__o21ai_1
X_06549_ final_design.reqhand.instruction\[31\] net973 vssd1 vssd1 vccd1 vccd1 _01500_
+ sky130_fd_sc_hd__or2_1
XANTENNA_fanout1161_X net1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout517_X net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09268_ net75 _04186_ vssd1 vssd1 vccd1 vccd1 _04187_ sky130_fd_sc_hd__or2_1
XFILLER_0_35_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08219_ final_design.cpu.reg_window\[267\] final_design.cpu.reg_window\[299\] net836
+ vssd1 vssd1 vccd1 vccd1 _03170_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09199_ net489 net318 vssd1 vssd1 vccd1 vccd1 _04118_ sky130_fd_sc_hd__nor2_1
XANTENNA__11718__A1 net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11230_ net646 net216 vssd1 vssd1 vccd1 vccd1 _05935_ sky130_fd_sc_hd__and2_1
XANTENNA__08044__C1 _01850_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout886_X net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1416 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11161_ net653 _05871_ _05873_ vssd1 vssd1 vccd1 vccd1 _05874_ sky130_fd_sc_hd__or3_1
X_10112_ _05023_ _05024_ _05006_ vssd1 vssd1 vccd1 vccd1 final_design.vga.v_next_count\[3\]
+ sky130_fd_sc_hd__and3b_1
XANTENNA__09139__A2 net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11092_ net59 _05799_ _05810_ _05812_ vssd1 vssd1 vccd1 vccd1 _05814_ sky130_fd_sc_hd__and4_1
XFILLER_0_41_1162 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11466__S net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10043_ _04571_ _04573_ _04388_ _04425_ vssd1 vssd1 vccd1 vccd1 _04962_ sky130_fd_sc_hd__o211a_1
XFILLER_0_76_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold40 final_design.cpu.reg_window\[18\] vssd1 vssd1 vccd1 vccd1 net1382 sky130_fd_sc_hd__dlygate4sd3_1
Xhold51 net146 vssd1 vssd1 vccd1 vccd1 net1393 sky130_fd_sc_hd__dlygate4sd3_1
Xhold62 net110 vssd1 vssd1 vccd1 vccd1 net1404 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_input25_A DAT_I[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold73 final_design.cpu.reg_window\[12\] vssd1 vssd1 vccd1 vccd1 net1415 sky130_fd_sc_hd__dlygate4sd3_1
Xhold84 net150 vssd1 vssd1 vccd1 vccd1 net1426 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_37_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold95 final_design.reqhand.instruction\[30\] vssd1 vssd1 vccd1 vccd1 net1437 sky130_fd_sc_hd__dlygate4sd3_1
X_13802_ clknet_leaf_59_clk _01033_ net1142 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[790\]
+ sky130_fd_sc_hd__dfrtp_1
X_11994_ net2445 net401 _06258_ net428 vssd1 vssd1 vccd1 vccd1 _00725_ sky130_fd_sc_hd__a22o_1
XANTENNA__13525__CLK clknet_leaf_58_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10457__B2 net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13733_ clknet_leaf_50_clk _00964_ net1181 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[721\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11654__B1 net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10945_ _05508_ _05672_ _05671_ vssd1 vssd1 vccd1 vccd1 _05673_ sky130_fd_sc_hd__o21bai_4
XANTENNA__12297__S net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13664_ clknet_leaf_11_clk _00895_ net1090 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[652\]
+ sky130_fd_sc_hd__dfrtp_1
X_10876_ net1004 _05606_ _05607_ net1032 net1358 vssd1 vssd1 vccd1 vccd1 _00193_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_45_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12777__8_A clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12615_ net2013 net2048 _05080_ vssd1 vssd1 vccd1 vccd1 _01308_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_41_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13595_ clknet_leaf_66_clk _00826_ net1063 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[583\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_41_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13675__CLK clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09459__X _04378_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1917 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12546_ _06209_ net342 net322 net1871 vssd1 vssd1 vccd1 vccd1 _01250_ sky130_fd_sc_hd__a22o_1
XFILLER_0_54_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11501__Y _06120_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09619__B net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12477_ _06137_ net345 net330 net2288 vssd1 vssd1 vccd1 vccd1 _01183_ sky130_fd_sc_hd__a22o_1
XANTENNA__11230__A net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_4 _05934_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14216_ net1274 vssd1 vssd1 vccd1 vccd1 gpio_oeb[28] sky130_fd_sc_hd__buf_2
X_11428_ net1727 net201 net313 vssd1 vssd1 vccd1 vccd1 _00325_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_39_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14147_ clknet_leaf_19_clk _01321_ net1112 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.data_to_VGA\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_11359_ net737 _03844_ _06047_ vssd1 vssd1 vccd1 vccd1 _06048_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09906__Y _04825_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10393__B1 net1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14078_ clknet_leaf_19_clk _01275_ net1157 vssd1 vssd1 vccd1 vccd1 final_design.reqhand.instruction\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13055__CLK clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11229__X _05934_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13029_ clknet_leaf_49_clk _00260_ net1184 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[17\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1060 final_design.reqhand.current_client\[3\] vssd1 vssd1 vccd1 vccd1 net1060
+ sky130_fd_sc_hd__buf_4
Xfanout1071 net1072 vssd1 vssd1 vccd1 vccd1 net1071 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11893__A0 net221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_6_clk_A clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1082 net1085 vssd1 vssd1 vccd1 vccd1 net1082 sky130_fd_sc_hd__clkbuf_2
XANTENNA__13117__RESET_B net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1093 net1096 vssd1 vssd1 vccd1 vccd1 net1093 sky130_fd_sc_hd__buf_2
X_08570_ net595 _03513_ _03517_ _02389_ vssd1 vssd1 vccd1 vccd1 _03521_ sky130_fd_sc_hd__o211a_2
X_07521_ _01631_ _02471_ vssd1 vssd1 vccd1 vccd1 _02472_ sky130_fd_sc_hd__nand2_1
XFILLER_0_72_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_18_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07849__C1 net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14236__1290 vssd1 vssd1 vccd1 vccd1 _14236__1290/HI net1290 sky130_fd_sc_hd__conb_1
XFILLER_0_37_1787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07452_ final_design.cpu.reg_window\[192\] final_design.cpu.reg_window\[224\] net895
+ vssd1 vssd1 vccd1 vccd1 _02403_ sky130_fd_sc_hd__mux2_1
XANTENNA__11405__A net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06403_ final_design.CPU_instr_adr\[29\] vssd1 vssd1 vccd1 vccd1 _01358_ sky130_fd_sc_hd__inv_2
XFILLER_0_57_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07383_ final_design.cpu.reg_window\[258\] final_design.cpu.reg_window\[290\] net919
+ vssd1 vssd1 vccd1 vccd1 _02334_ sky130_fd_sc_hd__mux2_1
X_09122_ net995 _01414_ vssd1 vssd1 vccd1 vccd1 _04041_ sky130_fd_sc_hd__nand2_2
XFILLER_0_2_1763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12070__B1 net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08273__X _03224_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09053_ net254 _03981_ net1013 vssd1 vssd1 vccd1 vccd1 _03982_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_26_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout212_A net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08004_ final_design.cpu.reg_window\[720\] final_design.cpu.reg_window\[752\] net843
+ vssd1 vssd1 vccd1 vccd1 _02955_ sky130_fd_sc_hd__mux2_1
XANTENNA__11140__A net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12782__13 clknet_leaf_28_clk vssd1 vssd1 vccd1 vccd1 net1323 sky130_fd_sc_hd__inv_2
Xhold510 final_design.cpu.reg_window\[703\] vssd1 vssd1 vccd1 vccd1 net1852 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold521 final_design.cpu.reg_window\[525\] vssd1 vssd1 vccd1 vccd1 net1863 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12373__A1 net219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold532 final_design.cpu.reg_window\[910\] vssd1 vssd1 vccd1 vccd1 net1874 sky130_fd_sc_hd__dlygate4sd3_1
Xhold543 final_design.cpu.reg_window\[745\] vssd1 vssd1 vccd1 vccd1 net1885 sky130_fd_sc_hd__dlygate4sd3_1
Xhold554 final_design.cpu.reg_window\[973\] vssd1 vssd1 vccd1 vccd1 net1896 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold565 final_design.cpu.reg_window\[585\] vssd1 vssd1 vccd1 vccd1 net1907 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1121_A net1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_2070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold576 final_design.cpu.reg_window\[475\] vssd1 vssd1 vccd1 vccd1 net1918 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07764__S net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold587 final_design.cpu.reg_window\[958\] vssd1 vssd1 vccd1 vccd1 net1929 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_55_2081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11794__B net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold598 final_design.cpu.reg_window\[236\] vssd1 vssd1 vccd1 vccd1 net1940 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_55_2092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09955_ _03488_ _04087_ _04873_ vssd1 vssd1 vccd1 vccd1 _04874_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout581_A net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout679_A net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08906_ net624 _03848_ _03849_ _03850_ net256 vssd1 vssd1 vccd1 vccd1 _03851_ sky130_fd_sc_hd__a311o_1
X_09886_ net263 _04793_ _04803_ _04804_ net450 vssd1 vssd1 vccd1 vccd1 _04805_ sky130_fd_sc_hd__a32o_2
XANTENNA_fanout1007_X net1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1210 final_design.cpu.reg_window\[365\] vssd1 vssd1 vccd1 vccd1 net2552 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13548__CLK clknet_leaf_45_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08837_ final_design.CPU_instr_adr\[10\] final_design.CPU_instr_adr\[9\] _03787_
+ vssd1 vssd1 vccd1 vccd1 _03788_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout846_A net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07552__A1 net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1917 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12428__A2 net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08595__S net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08768_ _03713_ _03718_ _03712_ vssd1 vssd1 vccd1 vccd1 _03719_ sky130_fd_sc_hd__a21o_1
XANTENNA__10439__B2 net245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11636__B1 net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07719_ net605 _02668_ _02643_ _01596_ vssd1 vssd1 vccd1 vccd1 _02670_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout634_X net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08699_ _02510_ _03647_ net659 vssd1 vssd1 vccd1 vccd1 _03650_ sky130_fd_sc_hd__nand3_4
XANTENNA__13698__CLK clknet_leaf_11_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10730_ _01382_ _05446_ _05467_ vssd1 vssd1 vccd1 vccd1 _05468_ sky130_fd_sc_hd__o21bai_1
X_10661_ net67 _05382_ _05386_ vssd1 vssd1 vccd1 vccd1 _05403_ sky130_fd_sc_hd__a21o_1
XANTENNA__11034__B net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout801_X net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07939__S net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12400_ _06098_ net347 net338 net2202 vssd1 vssd1 vccd1 vccd1 _01110_ sky130_fd_sc_hd__a22o_1
XANTENNA__11602__X _06157_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13380_ clknet_leaf_52_clk _00611_ net1174 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[368\]
+ sky130_fd_sc_hd__dfrtp_1
X_10592_ _05315_ _05318_ _05335_ vssd1 vssd1 vccd1 vccd1 _05337_ sky130_fd_sc_hd__a21oi_1
X_12331_ net571 _06262_ vssd1 vssd1 vccd1 vccd1 _06277_ sky130_fd_sc_hd__nor2_2
XANTENNA__06910__S0 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12262_ net579 _06191_ net511 net374 net1513 vssd1 vssd1 vccd1 vccd1 _00978_ sky130_fd_sc_hd__a32o_1
XFILLER_0_62_1803 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12364__A1 net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13078__CLK clknet_leaf_60_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11213_ _04772_ _04786_ net651 vssd1 vssd1 vccd1 vccd1 _05920_ sky130_fd_sc_hd__a21o_1
X_14001_ clknet_leaf_34_clk _01232_ net1242 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[989\]
+ sky130_fd_sc_hd__dfrtp_1
X_12193_ net1977 net180 net382 vssd1 vssd1 vccd1 vccd1 _00912_ sky130_fd_sc_hd__mux2_1
XANTENNA__10375__B1 net1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07466__S1 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13628__RESET_B net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07674__S net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11144_ net232 net2333 net314 vssd1 vssd1 vccd1 vccd1 _00275_ sky130_fd_sc_hd__mux2_1
XANTENNA__12116__A1 net196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11075_ _01388_ _05790_ _05795_ vssd1 vssd1 vccd1 vccd1 _05797_ sky130_fd_sc_hd__o21ba_1
XANTENNA__07218__S1 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10026_ net320 _04395_ _04403_ net319 _04944_ vssd1 vssd1 vccd1 vccd1 _04945_ sky130_fd_sc_hd__a221o_1
X_14201__1259 vssd1 vssd1 vccd1 vccd1 _14201__1259/HI net1259 sky130_fd_sc_hd__conb_1
XANTENNA__10142__A3 net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12915__CLK clknet_leaf_61_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12419__A2 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09190__A net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11977_ _06179_ net281 net405 net1641 vssd1 vssd1 vccd1 vccd1 _00710_ sky130_fd_sc_hd__a22o_1
XFILLER_0_34_1927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_47_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13716_ clknet_leaf_10_clk _00947_ net1102 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[704\]
+ sky130_fd_sc_hd__dfrtp_1
X_10928_ final_design.CPU_instr_adr\[23\] net1042 net802 vssd1 vssd1 vccd1 vccd1 _05657_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_50_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13647_ clknet_leaf_44_clk _00878_ net1208 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[635\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_32_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10859_ net80 _05568_ _05590_ vssd1 vssd1 vccd1 vccd1 _05591_ sky130_fd_sc_hd__a21o_1
XFILLER_0_54_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_1059 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13578_ clknet_leaf_60_clk _00809_ net1141 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[566\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12529_ _06191_ net354 net328 net1798 vssd1 vssd1 vccd1 vccd1 _01234_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_10_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_1925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_1471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10366__B1 net1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06989__A net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout308 net309 vssd1 vssd1 vccd1 vccd1 net308 sky130_fd_sc_hd__clkbuf_8
Xfanout319 _04084_ vssd1 vssd1 vccd1 vccd1 net319 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_61_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12107__A1 net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09740_ _04183_ _04658_ vssd1 vssd1 vccd1 vccd1 _04659_ sky130_fd_sc_hd__nand2_1
X_06952_ final_design.cpu.reg_window\[657\] final_design.cpu.reg_window\[689\] net928
+ vssd1 vssd1 vccd1 vccd1 _01903_ sky130_fd_sc_hd__mux2_1
.ends

