* NGSPICE file created from team_03_Wrapper.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_4 abstract view
.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_4 abstract view
.subckt sky130_fd_sc_hd__and3b_4 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_4 abstract view
.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_8 abstract view
.subckt sky130_fd_sc_hd__inv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_8 abstract view
.subckt sky130_fd_sc_hd__clkinv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_4 abstract view
.subckt sky130_fd_sc_hd__o211a_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_4 abstract view
.subckt sky130_fd_sc_hd__o31a_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_8 abstract view
.subckt sky130_fd_sc_hd__mux2_8 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_2 abstract view
.subckt sky130_fd_sc_hd__o32ai_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinvlp_4 abstract view
.subckt sky130_fd_sc_hd__clkinvlp_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__bufinv_16 abstract view
.subckt sky130_fd_sc_hd__bufinv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_2 abstract view
.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_4 abstract view
.subckt sky130_fd_sc_hd__o221a_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_1 abstract view
.subckt sky130_fd_sc_hd__clkinv_1 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_1 abstract view
.subckt sky130_fd_sc_hd__nand4b_1 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_2 abstract view
.subckt sky130_fd_sc_hd__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_4 abstract view
.subckt sky130_fd_sc_hd__o21ba_4 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_4 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_4 abstract view
.subckt sky130_fd_sc_hd__a221oi_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_4 abstract view
.subckt sky130_fd_sc_hd__a22o_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_2 abstract view
.subckt sky130_fd_sc_hd__o41a_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_2 abstract view
.subckt sky130_fd_sc_hd__a311o_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_2 abstract view
.subckt sky130_fd_sc_hd__a2111oi_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_4 abstract view
.subckt sky130_fd_sc_hd__nand4b_4 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_4 abstract view
.subckt sky130_fd_sc_hd__and4b_4 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311ai_4 abstract view
.subckt sky130_fd_sc_hd__o311ai_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_4 abstract view
.subckt sky130_fd_sc_hd__a221o_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_1 abstract view
.subckt sky130_fd_sc_hd__o2111ai_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_2 abstract view
.subckt sky130_fd_sc_hd__o311a_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_4 abstract view
.subckt sky130_fd_sc_hd__a311oi_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_4 abstract view
.subckt sky130_fd_sc_hd__o2111ai_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_4 abstract view
.subckt sky130_fd_sc_hd__o2111a_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_2 abstract view
.subckt sky130_fd_sc_hd__or4bb_2 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_4 abstract view
.subckt sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_2 abstract view
.subckt sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_1 abstract view
.subckt sky130_fd_sc_hd__nor4b_1 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311ai_2 abstract view
.subckt sky130_fd_sc_hd__o311ai_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_4 abstract view
.subckt sky130_fd_sc_hd__nand3b_4 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

.subckt team_03_Wrapper ACK_I ADR_O[0] ADR_O[10] ADR_O[11] ADR_O[12] ADR_O[13] ADR_O[14]
+ ADR_O[15] ADR_O[16] ADR_O[17] ADR_O[18] ADR_O[19] ADR_O[1] ADR_O[20] ADR_O[21] ADR_O[22]
+ ADR_O[23] ADR_O[24] ADR_O[25] ADR_O[26] ADR_O[27] ADR_O[28] ADR_O[29] ADR_O[2] ADR_O[30]
+ ADR_O[31] ADR_O[3] ADR_O[4] ADR_O[5] ADR_O[6] ADR_O[7] ADR_O[8] ADR_O[9] CYC_O DAT_I[0]
+ DAT_I[10] DAT_I[11] DAT_I[12] DAT_I[13] DAT_I[14] DAT_I[15] DAT_I[16] DAT_I[17]
+ DAT_I[18] DAT_I[19] DAT_I[1] DAT_I[20] DAT_I[21] DAT_I[22] DAT_I[23] DAT_I[24] DAT_I[25]
+ DAT_I[26] DAT_I[27] DAT_I[28] DAT_I[29] DAT_I[2] DAT_I[30] DAT_I[31] DAT_I[3] DAT_I[4]
+ DAT_I[5] DAT_I[6] DAT_I[7] DAT_I[8] DAT_I[9] DAT_O[0] DAT_O[10] DAT_O[11] DAT_O[12]
+ DAT_O[13] DAT_O[14] DAT_O[15] DAT_O[16] DAT_O[17] DAT_O[18] DAT_O[19] DAT_O[1] DAT_O[20]
+ DAT_O[21] DAT_O[22] DAT_O[23] DAT_O[24] DAT_O[25] DAT_O[26] DAT_O[27] DAT_O[28]
+ DAT_O[29] DAT_O[2] DAT_O[30] DAT_O[31] DAT_O[3] DAT_O[4] DAT_O[5] DAT_O[6] DAT_O[7]
+ DAT_O[8] DAT_O[9] SEL_O[0] SEL_O[1] SEL_O[2] SEL_O[3] STB_O WE_O gpio_in[0] gpio_in[10]
+ gpio_in[11] gpio_in[12] gpio_in[13] gpio_in[14] gpio_in[15] gpio_in[16] gpio_in[17]
+ gpio_in[18] gpio_in[19] gpio_in[1] gpio_in[20] gpio_in[21] gpio_in[22] gpio_in[23]
+ gpio_in[24] gpio_in[25] gpio_in[26] gpio_in[27] gpio_in[28] gpio_in[29] gpio_in[2]
+ gpio_in[30] gpio_in[31] gpio_in[32] gpio_in[33] gpio_in[34] gpio_in[35] gpio_in[36]
+ gpio_in[37] gpio_in[3] gpio_in[4] gpio_in[5] gpio_in[6] gpio_in[7] gpio_in[8] gpio_in[9]
+ gpio_oeb[0] gpio_oeb[10] gpio_oeb[11] gpio_oeb[12] gpio_oeb[13] gpio_oeb[14] gpio_oeb[15]
+ gpio_oeb[16] gpio_oeb[17] gpio_oeb[18] gpio_oeb[19] gpio_oeb[1] gpio_oeb[20] gpio_oeb[21]
+ gpio_oeb[22] gpio_oeb[23] gpio_oeb[24] gpio_oeb[25] gpio_oeb[26] gpio_oeb[27] gpio_oeb[28]
+ gpio_oeb[29] gpio_oeb[2] gpio_oeb[30] gpio_oeb[31] gpio_oeb[32] gpio_oeb[33] gpio_oeb[34]
+ gpio_oeb[35] gpio_oeb[36] gpio_oeb[37] gpio_oeb[3] gpio_oeb[4] gpio_oeb[5] gpio_oeb[6]
+ gpio_oeb[7] gpio_oeb[8] gpio_oeb[9] gpio_out[0] gpio_out[10] gpio_out[11] gpio_out[12]
+ gpio_out[13] gpio_out[14] gpio_out[15] gpio_out[16] gpio_out[17] gpio_out[18] gpio_out[19]
+ gpio_out[1] gpio_out[20] gpio_out[21] gpio_out[22] gpio_out[23] gpio_out[24] gpio_out[25]
+ gpio_out[26] gpio_out[27] gpio_out[28] gpio_out[29] gpio_out[2] gpio_out[30] gpio_out[31]
+ gpio_out[32] gpio_out[33] gpio_out[34] gpio_out[35] gpio_out[36] gpio_out[37] gpio_out[3]
+ gpio_out[4] gpio_out[5] gpio_out[6] gpio_out[7] gpio_out[8] gpio_out[9] irq[0] irq[1]
+ irq[2] la_data_in[0] la_data_in[10] la_data_in[11] la_data_in[12] la_data_in[13]
+ la_data_in[14] la_data_in[15] la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19]
+ la_data_in[1] la_data_in[20] la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24]
+ la_data_in[25] la_data_in[26] la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2]
+ la_data_in[30] la_data_in[31] la_data_in[3] la_data_in[4] la_data_in[5] la_data_in[6]
+ la_data_in[7] la_data_in[8] la_data_in[9] la_data_out[0] la_data_out[10] la_data_out[11]
+ la_data_out[12] la_data_out[13] la_data_out[14] la_data_out[15] la_data_out[16]
+ la_data_out[17] la_data_out[18] la_data_out[19] la_data_out[1] la_data_out[20] la_data_out[21]
+ la_data_out[22] la_data_out[23] la_data_out[24] la_data_out[25] la_data_out[26]
+ la_data_out[27] la_data_out[28] la_data_out[29] la_data_out[2] la_data_out[30] la_data_out[31]
+ la_data_out[3] la_data_out[4] la_data_out[5] la_data_out[6] la_data_out[7] la_data_out[8]
+ la_data_out[9] la_oenb[0] la_oenb[10] la_oenb[11] la_oenb[12] la_oenb[13] la_oenb[14]
+ la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19] la_oenb[1] la_oenb[20]
+ la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25] la_oenb[26] la_oenb[27]
+ la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31] la_oenb[3] la_oenb[4]
+ la_oenb[5] la_oenb[6] la_oenb[7] la_oenb[8] la_oenb[9] vccd1 vssd1 wb_clk_i wb_rst_i
+ wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14]
+ wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1]
+ wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25]
+ wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30]
+ wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8]
+ wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13]
+ wbs_dat_i[14] wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19]
+ wbs_dat_i[1] wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24]
+ wbs_dat_i[25] wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2]
+ wbs_dat_i[30] wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6]
+ wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11]
+ wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17]
+ wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22]
+ wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28]
+ wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4]
+ wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0] wbs_sel_i[1]
+ wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
XANTENNA__08326__A3 _04267_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09671_ _05089_ _05091_ _05095_ _05098_ net554 net567 vssd1 vssd1 vccd1 vccd1 _05613_
+ sky130_fd_sc_hd__mux4_1
X_06883_ team_03_WB.instance_to_wrap.core.decoder.inst\[28\] team_03_WB.instance_to_wrap.core.decoder.inst\[27\]
+ _02824_ vssd1 vssd1 vccd1 vccd1 _02825_ sky130_fd_sc_hd__or3_1
XANTENNA__11866__B1 net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08731__B1 net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13615__A net1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08622_ _04558_ _04563_ net874 vssd1 vssd1 vccd1 vccd1 _04564_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10958__B _05784_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11881__A3 net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11618__B1 net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08553_ net854 _04493_ _04494_ vssd1 vssd1 vccd1 vccd1 _04495_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_46_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07298__B1 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07504_ _03443_ _03445_ net810 vssd1 vssd1 vccd1 vccd1 _03446_ sky130_fd_sc_hd__o21a_1
X_08484_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[827\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[795\]
+ net988 vssd1 vssd1 vccd1 vccd1 _04426_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07435_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[148\] net764
+ net726 _03376_ vssd1 vssd1 vccd1 vccd1 _03377_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_21_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1071_A net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_174_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout427_A _04079_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13350__A net1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09099__X _05041_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_851 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08247__C1 net1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07366_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[828\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[796\]
+ net759 vssd1 vssd1 vccd1 vccd1 _03308_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_135_3141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_135_3152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09105_ net1051 team_03_WB.instance_to_wrap.core.register_file.registers_state\[78\]
+ net1001 team_03_WB.instance_to_wrap.core.register_file.registers_state\[110\] net940
+ vssd1 vssd1 vccd1 vccd1 _05047_ sky130_fd_sc_hd__a221o_1
XFILLER_0_73_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_150_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_165_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_hold1277_A team_03_WB.instance_to_wrap.CPU_DAT_O\[2\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_07297_ net1167 _03237_ _03238_ _03234_ vssd1 vssd1 vccd1 vccd1 _03239_ sky130_fd_sc_hd__o22a_1
XFILLER_0_32_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_761 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_463 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1336_A net1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09974__S net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09036_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[880\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[848\]
+ net984 vssd1 vssd1 vccd1 vccd1 _04978_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout796_A net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11149__A2 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold340 net181 vssd1 vssd1 vccd1 vccd1 net1833 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06899__A _02837_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1124_X net1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold351 team_03_WB.instance_to_wrap.core.register_file.registers_state\[388\] vssd1
+ vssd1 vccd1 vccd1 net1844 sky130_fd_sc_hd__dlygate4sd3_1
Xhold362 team_03_WB.instance_to_wrap.CPU_DAT_I\[29\] vssd1 vssd1 vccd1 vccd1 net1855
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07494__S net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold373 net192 vssd1 vssd1 vccd1 vccd1 net1866 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_159_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold384 _02599_ vssd1 vssd1 vccd1 vccd1 net1877 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09275__A _04954_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07222__B1 net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09762__A2 _05073_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold395 team_03_WB.instance_to_wrap.core.register_file.registers_state\[391\] vssd1
+ vssd1 vccd1 vccd1 net1888 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout963_A net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout584_X net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07773__A1 net1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout820 _02847_ vssd1 vssd1 vccd1 vccd1 net820 sky130_fd_sc_hd__buf_6
XANTENNA__08970__B1 net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout831 _06558_ vssd1 vssd1 vccd1 vccd1 net831 sky130_fd_sc_hd__clkbuf_8
X_09938_ _05873_ net1750 net292 vssd1 vssd1 vccd1 vccd1 _02758_ sky130_fd_sc_hd__mux2_1
Xfanout842 net843 vssd1 vssd1 vccd1 vccd1 net842 sky130_fd_sc_hd__buf_4
Xfanout853 _04096_ vssd1 vssd1 vccd1 vccd1 net853 sky130_fd_sc_hd__buf_4
Xfanout864 net866 vssd1 vssd1 vccd1 vccd1 net864 sky130_fd_sc_hd__clkbuf_8
Xfanout875 _04081_ vssd1 vssd1 vccd1 vccd1 net875 sky130_fd_sc_hd__buf_4
Xfanout886 net887 vssd1 vssd1 vccd1 vccd1 net886 sky130_fd_sc_hd__buf_4
XANTENNA__11029__B net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11857__B1 net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09869_ net581 _05597_ _05804_ _05810_ vssd1 vssd1 vccd1 vccd1 _05811_ sky130_fd_sc_hd__a31oi_4
Xfanout897 net900 vssd1 vssd1 vccd1 vccd1 net897 sky130_fd_sc_hd__buf_2
XANTENNA_fanout751_X net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07525__A1 net1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1040 team_03_WB.instance_to_wrap.core.register_file.registers_state\[734\] vssd1
+ vssd1 vccd1 vccd1 net2533 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout849_X net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1051 team_03_WB.instance_to_wrap.core.register_file.registers_state\[493\] vssd1
+ vssd1 vccd1 vccd1 net2544 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1062 team_03_WB.instance_to_wrap.core.register_file.registers_state\[688\] vssd1
+ vssd1 vccd1 vccd1 net2555 sky130_fd_sc_hd__dlygate4sd3_1
X_11900_ net645 _06709_ net477 net374 net2120 vssd1 vssd1 vccd1 vccd1 _01641_ sky130_fd_sc_hd__a32o_1
XFILLER_0_169_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1073 team_03_WB.instance_to_wrap.core.register_file.registers_state\[715\] vssd1
+ vssd1 vccd1 vccd1 net2566 sky130_fd_sc_hd__dlygate4sd3_1
X_12880_ net1409 vssd1 vssd1 vccd1 vccd1 _00644_ sky130_fd_sc_hd__inv_2
Xhold1084 net205 vssd1 vssd1 vccd1 vccd1 net2577 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_107_2564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_2575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1095 team_03_WB.instance_to_wrap.core.register_file.registers_state\[155\] vssd1
+ vssd1 vccd1 vccd1 net2588 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_29_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11831_ net647 _06666_ net453 net323 net1872 vssd1 vssd1 vccd1 vccd1 _01708_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_159_3631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_159_3642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14550_ clknet_leaf_151_wb_clk_i _02314_ _00915_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[904\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_96_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07289__B1 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11762_ _06590_ net469 net333 net2661 vssd1 vssd1 vccd1 vccd1 _01775_ sky130_fd_sc_hd__a22o_1
XFILLER_0_68_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13501_ net1327 vssd1 vssd1 vccd1 vccd1 _01265_ sky130_fd_sc_hd__inv_2
X_10713_ team_03_WB.instance_to_wrap.core.pc.current_pc\[23\] _05518_ net603 vssd1
+ vssd1 vccd1 vccd1 _06347_ sky130_fd_sc_hd__mux2_1
X_14481_ clknet_leaf_139_wb_clk_i _02245_ _00846_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[835\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_165_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_339 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11693_ _06735_ net382 net339 net2035 vssd1 vssd1 vccd1 vccd1 _01841_ sky130_fd_sc_hd__a22o_1
XFILLER_0_153_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11332__X _06718_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13260__A net1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13432_ net1432 vssd1 vssd1 vccd1 vccd1 _01196_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12034__B1 net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input92_A wbs_adr_i[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10644_ net1212 team_03_WB.instance_to_wrap.CPU_DAT_O\[17\] net844 vssd1 vssd1 vccd1
+ vccd1 _02484_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_884 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11388__A2 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_172_3897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13363_ net1329 vssd1 vssd1 vccd1 vccd1 _01127_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10575_ net1718 net534 net601 _05885_ vssd1 vssd1 vccd1 vccd1 _02548_ sky130_fd_sc_hd__a22o_1
XFILLER_0_23_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15102_ net912 vssd1 vssd1 vccd1 vccd1 net261 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12314_ net1377 vssd1 vssd1 vccd1 vccd1 _00078_ sky130_fd_sc_hd__inv_2
XFILLER_0_51_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07461__B1 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13294_ net1328 vssd1 vssd1 vccd1 vccd1 _01058_ sky130_fd_sc_hd__inv_2
XFILLER_0_121_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15033_ clknet_leaf_91_wb_clk_i _02753_ _01398_ vssd1 vssd1 vccd1 vccd1 net189 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_146_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11919__S net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_792 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12245_ net1703 vssd1 vssd1 vccd1 vccd1 _01412_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09753__A2 _03724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12176_ net1592 vssd1 vssd1 vccd1 vccd1 _02377_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__08961__B1 net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11560__A2 net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11127_ net627 _06638_ vssd1 vssd1 vccd1 vccd1 _06639_ sky130_fd_sc_hd__nor2_1
XANTENNA__06972__C1 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11848__A0 net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11058_ net506 net653 _06606_ net422 net2100 vssd1 vssd1 vccd1 vccd1 _02276_ sky130_fd_sc_hd__a32o_1
XFILLER_0_3_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07516__A1 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_60_wb_clk_i clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_60_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08713__B1 net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11654__S net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10009_ _02888_ net1890 net290 vssd1 vssd1 vccd1 vccd1 _02705_ sky130_fd_sc_hd__mux2_1
XANTENNA__10520__B1 net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14817_ clknet_leaf_89_wb_clk_i net1783 _01182_ vssd1 vssd1 vccd1 vccd1 net137 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_118_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_171_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14748_ clknet_leaf_62_wb_clk_i net1669 _01113_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08477__C1 net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07819__A2 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_48_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_15_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14679_ clknet_leaf_83_wb_clk_i _02443_ _01044_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.ADR_I\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_156_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06991__B net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_926 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07220_ _03160_ _03161_ net1160 vssd1 vssd1 vccd1 vccd1 _03162_ sky130_fd_sc_hd__o21a_1
XFILLER_0_129_599 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_15_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12025__B1 net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08229__C1 net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07151_ net1204 team_03_WB.instance_to_wrap.core.register_file.registers_state\[352\]
+ net885 _03092_ vssd1 vssd1 vccd1 vccd1 _03093_ sky130_fd_sc_hd__a31o_1
XFILLER_0_89_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_171_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10587__B1 net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07082_ net614 _03023_ _02995_ vssd1 vssd1 vccd1 vccd1 _03024_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_120_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_152_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_1144 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12514__A net1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1132 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_628 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11000__A1 net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_39_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11551__A2 net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07984_ net1107 team_03_WB.instance_to_wrap.core.register_file.registers_state\[880\]
+ net901 vssd1 vssd1 vccd1 vccd1 _03926_ sky130_fd_sc_hd__or3_1
X_09723_ _03759_ _04893_ vssd1 vssd1 vccd1 vccd1 _05665_ sky130_fd_sc_hd__nor2_1
XANTENNA__11839__B1 net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06935_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[548\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[516\]
+ net775 vssd1 vssd1 vccd1 vccd1 _02877_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_87_wb_clk_i_A clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout377_A _06812_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_87_2158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09654_ net594 _05584_ _05585_ _05595_ vssd1 vssd1 vccd1 vccd1 _05596_ sky130_fd_sc_hd__o31a_2
XTAP_TAPCELL_ROW_87_2169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10511__B1 net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06866_ team_03_WB.instance_to_wrap.core.control_logic.instruction\[5\] _02794_ _02806_
+ vssd1 vssd1 vccd1 vccd1 _02808_ sky130_fd_sc_hd__and3_4
XFILLER_0_97_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08605_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[933\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[901\]
+ net992 vssd1 vssd1 vccd1 vccd1 _04547_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_26_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09585_ _05420_ _05525_ net568 vssd1 vssd1 vccd1 vccd1 _05527_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_26_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_65_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1286_A net1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08536_ net542 _04476_ vssd1 vssd1 vccd1 vccd1 _04478_ sky130_fd_sc_hd__nor2_1
XANTENNA__08468__C1 net1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_102_2461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_2472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout711_A net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout332_X net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08467_ net1226 team_03_WB.instance_to_wrap.core.register_file.registers_state\[348\]
+ net951 team_03_WB.instance_to_wrap.core.register_file.registers_state\[380\] net1070
+ vssd1 vssd1 vccd1 vccd1 _04409_ sky130_fd_sc_hd__o221a_1
XFILLER_0_18_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout809_A net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1074_X net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_163_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07418_ net1084 team_03_WB.instance_to_wrap.core.register_file.registers_state\[660\]
+ net889 net1125 vssd1 vssd1 vccd1 vccd1 _03360_ sky130_fd_sc_hd__a211o_1
XANTENNA__12016__B1 net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08398_ _04334_ _04339_ net874 vssd1 vssd1 vccd1 vccd1 _04340_ sky130_fd_sc_hd__mux2_1
XANTENNA__07691__B1 net1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_350 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07349_ net1170 team_03_WB.instance_to_wrap.core.register_file.registers_state\[348\]
+ net757 team_03_WB.instance_to_wrap.core.register_file.registers_state\[380\] net1123
+ vssd1 vssd1 vccd1 vccd1 _03291_ sky130_fd_sc_hd__o221a_1
XFILLER_0_163_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10578__B1 net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1241_X net1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_150_3447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_150_3458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1339_X net1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10360_ _06092_ _06187_ _06101_ vssd1 vssd1 vccd1 vccd1 _06193_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_143_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11739__S net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout799_X net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07994__A1 net1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09019_ _04959_ _04960_ net864 vssd1 vssd1 vccd1 vccd1 _04961_ sky130_fd_sc_hd__a21o_1
X_10291_ _06131_ _06132_ vssd1 vssd1 vccd1 vccd1 _06133_ sky130_fd_sc_hd__or2_1
XANTENNA__10643__S net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12424__A net1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12030_ _06771_ net475 net362 net2587 vssd1 vssd1 vccd1 vccd1 _01515_ sky130_fd_sc_hd__a22o_1
XANTENNA__07518__A team_03_WB.instance_to_wrap.core.decoder.inst\[26\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold170 net174 vssd1 vssd1 vccd1 vccd1 net1663 sky130_fd_sc_hd__dlygate4sd3_1
Xhold181 _02614_ vssd1 vssd1 vccd1 vccd1 net1674 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout966_X net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold192 _02587_ vssd1 vssd1 vccd1 vccd1 net1685 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11542__A2 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08943__B1 net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout650 net651 vssd1 vssd1 vccd1 vccd1 net650 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_109_2615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout661 net663 vssd1 vssd1 vccd1 vccd1 net661 sky130_fd_sc_hd__buf_4
Xfanout672 net673 vssd1 vssd1 vccd1 vccd1 net672 sky130_fd_sc_hd__clkbuf_4
Xfanout683 _05915_ vssd1 vssd1 vccd1 vccd1 net683 sky130_fd_sc_hd__buf_2
X_13981_ clknet_leaf_25_wb_clk_i _01745_ _00346_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[335\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout694 _06562_ vssd1 vssd1 vccd1 vccd1 net694 sky130_fd_sc_hd__buf_6
XFILLER_0_137_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12932_ net1366 vssd1 vssd1 vccd1 vccd1 _00696_ sky130_fd_sc_hd__inv_2
XFILLER_0_77_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_126_2962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10502__B1 net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08349__A net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08171__A1 net1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_228 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12863_ net1347 vssd1 vssd1 vccd1 vccd1 _00627_ sky130_fd_sc_hd__inv_2
XFILLER_0_38_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11058__A1 net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14602_ clknet_leaf_6_wb_clk_i _02366_ _00967_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[956\]
+ sky130_fd_sc_hd__dfstp_1
X_11814_ _06642_ net475 net326 net1836 vssd1 vssd1 vccd1 vccd1 _01725_ sky130_fd_sc_hd__a22o_1
X_12794_ net1372 vssd1 vssd1 vccd1 vccd1 _00558_ sky130_fd_sc_hd__inv_2
XFILLER_0_69_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_164_Left_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_174_3937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14533_ clknet_leaf_39_wb_clk_i _02297_ _00898_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[887\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_174_3948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11745_ _06566_ net462 net331 net2426 vssd1 vssd1 vccd1 vccd1 _01792_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_174_3959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14464_ clknet_leaf_2_wb_clk_i _02228_ _00829_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[818\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_12_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11676_ net1042 net694 _06803_ vssd1 vssd1 vccd1 vccd1 _06806_ sky130_fd_sc_hd__or3_4
XFILLER_0_36_350 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13415_ net1428 vssd1 vssd1 vccd1 vccd1 _01179_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10627_ net1574 team_03_WB.instance_to_wrap.CPU_DAT_O\[2\] net842 vssd1 vssd1 vccd1
+ vccd1 _02501_ sky130_fd_sc_hd__mux2_1
X_14395_ clknet_leaf_123_wb_clk_i _02159_ _00760_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[749\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10569__B1 net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_528 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_1132 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10324__B1_N net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13346_ net1325 vssd1 vssd1 vccd1 vccd1 _01110_ sky130_fd_sc_hd__inv_2
X_10558_ net1729 net533 net600 _05868_ vssd1 vssd1 vccd1 vccd1 _02565_ sky130_fd_sc_hd__a22o_1
XFILLER_0_24_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11649__S net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13277_ net1406 vssd1 vssd1 vccd1 vccd1 _01041_ sky130_fd_sc_hd__inv_2
X_10489_ net1812 net1029 net906 team_03_WB.instance_to_wrap.ADR_I\[17\] vssd1 vssd1
+ vccd1 vccd1 _02620_ sky130_fd_sc_hd__a22o_1
XANTENNA__09187__B1 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_173_Left_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15016_ clknet_leaf_95_wb_clk_i _02736_ _01381_ vssd1 vssd1 vccd1 vccd1 net203 sky130_fd_sc_hd__dfrtp_1
XANTENNA__09119__S net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07428__A net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12228_ net1567 vssd1 vssd1 vccd1 vccd1 _01429_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_clkbuf_leaf_121_wb_clk_i_A clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__07737__A1 team_03_WB.instance_to_wrap.core.decoder.inst\[13\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11533__A2 net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12159_ net1542 vssd1 vssd1 vccd1 vccd1 _02394_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__10741__B1 net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07832__S1 net1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_34_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08698__C1 net1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11836__A3 net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_4_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_87_740 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09370_ _04071_ _05159_ vssd1 vssd1 vccd1 vccd1 _05312_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_82_2055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_89 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14992__Q team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[11\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08321_ net944 _04262_ vssd1 vssd1 vccd1 vccd1 _04263_ sky130_fd_sc_hd__or2_1
XANTENNA__10728__S net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_363 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08252_ net1226 team_03_WB.instance_to_wrap.core.register_file.registers_state\[594\]
+ net950 team_03_WB.instance_to_wrap.core.register_file.registers_state\[626\] net916
+ vssd1 vssd1 vccd1 vccd1 _04194_ sky130_fd_sc_hd__o221a_1
XFILLER_0_7_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11413__A _06478_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07673__B1 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07203_ net806 _03143_ _03144_ vssd1 vssd1 vccd1 vccd1 _03145_ sky130_fd_sc_hd__or3_1
X_08183_ net1231 team_03_WB.instance_to_wrap.core.register_file.registers_state\[83\]
+ net957 team_03_WB.instance_to_wrap.core.register_file.registers_state\[115\] net918
+ vssd1 vssd1 vccd1 vccd1 _04125_ sky130_fd_sc_hd__o221a_1
XFILLER_0_144_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_160_wb_clk_i_A clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12013__A3 net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08848__S0 net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_854 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_848 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07134_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[928\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[896\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[800\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[768\]
+ net785 net1135 vssd1 vssd1 vccd1 vccd1 _03076_ sky130_fd_sc_hd__mux4_1
XANTENNA__07425__B1 net1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11221__B2 net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07976__A1 net1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11772__A2 net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07065_ net1193 team_03_WB.instance_to_wrap.core.register_file.registers_state\[130\]
+ vssd1 vssd1 vccd1 vccd1 _03007_ sky130_fd_sc_hd__or2_1
Xoutput220 net220 vssd1 vssd1 vccd1 vccd1 gpio_out[23] sky130_fd_sc_hd__buf_2
Xoutput231 net231 vssd1 vssd1 vccd1 vccd1 gpio_out[34] sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout1034_A net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput242 net242 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[12] sky130_fd_sc_hd__buf_2
XFILLER_0_11_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_58_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput253 net253 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[27] sky130_fd_sc_hd__buf_2
XANTENNA_clkbuf_4_15__f_wb_clk_i_A clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout494_A net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07728__A1 net1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08925__B1 net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_2209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1201_A net1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout661_A net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07967_ net750 _03905_ _03906_ _03907_ _03908_ vssd1 vssd1 vccd1 vccd1 _03909_ sky130_fd_sc_hd__o32a_1
XANTENNA__09025__S0 net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_156_70 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout759_A net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09706_ _05211_ _05276_ _05209_ vssd1 vssd1 vccd1 vccd1 _05648_ sky130_fd_sc_hd__a21oi_2
XANTENNA__13075__A net1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11288__A1 net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06918_ net1106 team_03_WB.instance_to_wrap.core.register_file.registers_state\[196\]
+ net804 team_03_WB.instance_to_wrap.core.register_file.registers_state\[228\] net734
+ vssd1 vssd1 vccd1 vccd1 _02860_ sky130_fd_sc_hd__a221o_1
XANTENNA__08153__A1 net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07898_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[399\] net781
+ _03839_ vssd1 vssd1 vccd1 vccd1 _03840_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_104_2512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09637_ _05406_ _05408_ net553 vssd1 vssd1 vccd1 vccd1 _05579_ sky130_fd_sc_hd__mux2_1
X_06849_ team_03_WB.instance_to_wrap.core.decoder.inst\[13\] vssd1 vssd1 vccd1 vccd1
+ _02792_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout1191_X net1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout926_A net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09568_ _03904_ _04235_ _05509_ _02945_ vssd1 vssd1 vccd1 vccd1 _05510_ sky130_fd_sc_hd__o22a_1
XANTENNA__09102__B1 net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_2870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08519_ net867 _04460_ _04455_ vssd1 vssd1 vccd1 vccd1 _04461_ sky130_fd_sc_hd__o21ai_1
XANTENNA__10638__S net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09499_ net568 _05440_ _05439_ vssd1 vssd1 vccd1 vccd1 _05441_ sky130_fd_sc_hd__a21oi_2
XANTENNA__09653__A1 net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout714_X net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10865__C _06463_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11530_ net2226 net485 _06783_ net512 vssd1 vssd1 vccd1 vccd1 _01981_ sky130_fd_sc_hd__a22o_1
XANTENNA__11460__A1 net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08861__C1 net1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_137_Right_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11461_ net630 _06586_ vssd1 vssd1 vccd1 vccd1 _06767_ sky130_fd_sc_hd__and2_1
XFILLER_0_52_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13200_ net1412 vssd1 vssd1 vccd1 vccd1 _00964_ sky130_fd_sc_hd__inv_2
XANTENNA__11610__X _06804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10412_ net304 net303 _06234_ _06235_ vssd1 vssd1 vccd1 vccd1 _06236_ sky130_fd_sc_hd__a22o_1
XFILLER_0_151_859 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11392_ net506 net634 _06748_ net402 net2007 vssd1 vssd1 vccd1 vccd1 _02084_ sky130_fd_sc_hd__a32o_1
X_14180_ clknet_leaf_15_wb_clk_i _01944_ _00545_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[534\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_34_898 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07967__A1 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_150_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13131_ net1288 vssd1 vssd1 vccd1 vccd1 _00895_ sky130_fd_sc_hd__inv_2
XANTENNA__11763__A2 net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_1979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10343_ _06148_ _06149_ _06178_ vssd1 vssd1 vccd1 vccd1 _06179_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_131_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10971__A0 net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_1052 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10274_ _06115_ vssd1 vssd1 vccd1 vccd1 _06116_ sky130_fd_sc_hd__inv_2
XFILLER_0_143_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input55_A gpio_in[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13062_ net1300 vssd1 vssd1 vccd1 vccd1 _00826_ sky130_fd_sc_hd__inv_2
XFILLER_0_143_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07719__A1 net1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12013_ net619 _06572_ net452 net359 net2117 vssd1 vssd1 vccd1 vccd1 _01532_ sky130_fd_sc_hd__a32o_1
XFILLER_0_40_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1401 net1408 vssd1 vssd1 vccd1 vccd1 net1401 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_167_3796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1412 net1413 vssd1 vssd1 vccd1 vccd1 net1412 sky130_fd_sc_hd__buf_4
Xfanout1423 net1426 vssd1 vssd1 vccd1 vccd1 net1423 sky130_fd_sc_hd__buf_4
XFILLER_0_100_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1434 net1435 vssd1 vssd1 vccd1 vccd1 net1434 sky130_fd_sc_hd__buf_2
XANTENNA__08392__A1 net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout480 net481 vssd1 vssd1 vccd1 vccd1 net480 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_75_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_6_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout491 net492 vssd1 vssd1 vccd1 vccd1 net491 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09182__B _03062_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13964_ clknet_leaf_16_wb_clk_i _01728_ _00329_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[318\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input10_X net10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12915_ net1271 vssd1 vssd1 vccd1 vccd1 _00679_ sky130_fd_sc_hd__inv_2
X_13895_ clknet_leaf_113_wb_clk_i _01659_ _00260_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[249\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_115_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11932__S net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12846_ net1303 vssd1 vssd1 vccd1 vccd1 _00610_ sky130_fd_sc_hd__inv_2
XFILLER_0_61_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12777_ net1257 vssd1 vssd1 vccd1 vccd1 _00541_ sky130_fd_sc_hd__inv_2
XANTENNA__07104__C1 net1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12329__A net1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_659 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_1126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14516_ clknet_leaf_132_wb_clk_i _02280_ _00881_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[870\]
+ sky130_fd_sc_hd__dfrtp_1
X_11728_ net1894 _06491_ net336 vssd1 vssd1 vccd1 vccd1 _01808_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08852__C1 net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11451__B2 net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14447_ clknet_leaf_143_wb_clk_i _02211_ _00812_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[801\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_104_Right_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11659_ net2460 _06622_ net345 vssd1 vssd1 vccd1 vccd1 _01874_ sky130_fd_sc_hd__mux2_1
XFILLER_0_141_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_331 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07407__B1 net1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_876 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14378_ clknet_leaf_0_wb_clk_i _02142_ _00743_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[732\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold906 team_03_WB.instance_to_wrap.core.register_file.registers_state\[78\] vssd1
+ vssd1 vccd1 vccd1 net2399 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold917 team_03_WB.instance_to_wrap.core.register_file.registers_state\[383\] vssd1
+ vssd1 vccd1 vccd1 net2410 sky130_fd_sc_hd__dlygate4sd3_1
X_13329_ net1325 vssd1 vssd1 vccd1 vccd1 _01093_ sky130_fd_sc_hd__inv_2
XANTENNA__09698__A2_N _03864_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold928 team_03_WB.instance_to_wrap.core.register_file.registers_state\[859\] vssd1
+ vssd1 vccd1 vccd1 net2421 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08080__B1 net1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold939 team_03_WB.instance_to_wrap.core.register_file.registers_state\[188\] vssd1
+ vssd1 vccd1 vccd1 net2432 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_150_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07422__A3 net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09925__X _05867_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_36_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12999__A net1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08907__B1 net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08870_ _04809_ _04810_ _04770_ vssd1 vssd1 vccd1 vccd1 _04812_ sky130_fd_sc_hd__o21ai_1
XANTENNA__10714__B1 net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06918__C1 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14987__Q team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[6\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07821_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[170\] net764
+ net741 _03762_ vssd1 vssd1 vccd1 vccd1 _03763_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_32_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07164__Y _03106_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12003__S net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07752_ net1195 team_03_WB.instance_to_wrap.core.register_file.registers_state\[332\]
+ vssd1 vssd1 vccd1 vccd1 _03694_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_84_2106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07683_ net1174 team_03_WB.instance_to_wrap.core.register_file.registers_state\[574\]
+ net880 vssd1 vssd1 vccd1 vccd1 _03625_ sky130_fd_sc_hd__and3_1
XFILLER_0_79_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09422_ _04816_ _05343_ _05361_ _05362_ vssd1 vssd1 vccd1 vccd1 _05364_ sky130_fd_sc_hd__o211a_1
XANTENNA__10493__A2 net1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_436 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06936__S net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09353_ _05294_ vssd1 vssd1 vccd1 vccd1 _05295_ sky130_fd_sc_hd__inv_2
XANTENNA__10458__S net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09635__A1 net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11143__A net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08304_ net1237 team_03_WB.instance_to_wrap.core.register_file.registers_state\[344\]
+ net972 team_03_WB.instance_to_wrap.core.register_file.registers_state\[376\] net1073
+ vssd1 vssd1 vccd1 vccd1 _04246_ sky130_fd_sc_hd__o221a_1
XANTENNA__07646__B1 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11442__A1 net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09284_ _04922_ _05225_ vssd1 vssd1 vccd1 vccd1 _05226_ sky130_fd_sc_hd__and2_1
XFILLER_0_7_520 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08843__C1 net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08235_ net850 _04170_ _04176_ vssd1 vssd1 vccd1 vccd1 _04177_ sky130_fd_sc_hd__and3_1
XANTENNA__10982__A net1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_686 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1151_A net1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout507_A net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_848 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1249_A net1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_166_1074 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08166_ net1230 team_03_WB.instance_to_wrap.core.register_file.registers_state\[724\]
+ net959 team_03_WB.instance_to_wrap.core.register_file.registers_state\[756\] net935
+ vssd1 vssd1 vccd1 vccd1 _04108_ sky130_fd_sc_hd__o221a_1
XFILLER_0_67_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07949__A1 net1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11745__A2 net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07117_ net723 _03058_ _03043_ vssd1 vssd1 vccd1 vccd1 _03059_ sky130_fd_sc_hd__o21a_4
XFILLER_0_31_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08097_ net1173 team_03_WB.instance_to_wrap.core.register_file.registers_state\[218\]
+ net760 team_03_WB.instance_to_wrap.core.register_file.registers_state\[250\] net739
+ vssd1 vssd1 vccd1 vccd1 _04039_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_56_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09982__S net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07048_ team_03_WB.instance_to_wrap.core.decoder.inst\[10\] _02808_ _02818_ net1148
+ vssd1 vssd1 vccd1 vccd1 _02990_ sky130_fd_sc_hd__a22oi_4
Xclkload90 clknet_leaf_72_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload90/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_24_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout876_A net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout497_X net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09166__A3 _04893_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10921__S net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09020__C1 net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1204_X net1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08374__A1 net1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_3346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input2_X net2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_3357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout664_X net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08999_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[810\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[778\]
+ net955 vssd1 vssd1 vccd1 vccd1 _04941_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_188_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_188_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_3_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_162_3693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08126__A1 net1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_2910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_117_wb_clk_i clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_117_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_168_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10961_ team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[2\] net306 vssd1 vssd1
+ vccd1 vccd1 _06542_ sky130_fd_sc_hd__and2_1
XANTENNA__07234__C net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout831_X net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11130__B1 net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout929_X net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12700_ net1418 vssd1 vssd1 vccd1 vccd1 _00464_ sky130_fd_sc_hd__inv_2
XANTENNA__10484__A2 net1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13680_ clknet_leaf_160_wb_clk_i _01444_ _00045_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[34\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07885__B1 net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10892_ team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[15\] _05865_ net317 _06403_
+ net686 vssd1 vssd1 vccd1 vccd1 _06486_ sky130_fd_sc_hd__a41o_1
XFILLER_0_35_1148 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12631_ net1386 vssd1 vssd1 vccd1 vccd1 _00395_ sky130_fd_sc_hd__inv_2
XFILLER_0_109_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09087__C1 net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09626__A1 _03024_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11053__A net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07637__B1 net1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12562_ net1397 vssd1 vssd1 vccd1 vccd1 _00326_ sky130_fd_sc_hd__inv_2
XFILLER_0_93_584 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14301_ clknet_leaf_26_wb_clk_i _02065_ _00666_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[655\]
+ sky130_fd_sc_hd__dfrtp_1
X_11513_ _06629_ net2596 net391 vssd1 vssd1 vccd1 vccd1 _01993_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12493_ net1332 vssd1 vssd1 vccd1 vccd1 _00257_ sky130_fd_sc_hd__inv_2
XFILLER_0_124_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_150_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14232_ clknet_leaf_3_wb_clk_i _01996_ _00597_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[586\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_117_2769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11444_ net2373 net394 _06761_ net512 vssd1 vssd1 vccd1 vccd1 _02045_ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_684 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11199__S net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11736__A2 net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14163_ clknet_leaf_98_wb_clk_i _01927_ _00528_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[517\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_169_3836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11375_ net1247 net837 net270 net668 vssd1 vssd1 vccd1 vccd1 _06740_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_169_3847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10944__B1 net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13114_ net1377 vssd1 vssd1 vccd1 vccd1 _00878_ sky130_fd_sc_hd__inv_2
XFILLER_0_81_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10326_ _06164_ _06165_ team_03_WB.instance_to_wrap.core.pc.current_pc\[29\] net677
+ vssd1 vssd1 vccd1 vccd1 _02663_ sky130_fd_sc_hd__o2bb2a_1
X_14094_ clknet_leaf_131_wb_clk_i _01858_ _00459_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[448\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11927__S net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13045_ net1277 vssd1 vssd1 vccd1 vccd1 _00809_ sky130_fd_sc_hd__inv_2
X_10257_ _04324_ team_03_WB.instance_to_wrap.core.pc.current_pc\[22\] net672 vssd1
+ vssd1 vccd1 vccd1 _06099_ sky130_fd_sc_hd__mux2_1
XANTENNA__09905__B _05623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1220 net1225 vssd1 vssd1 vccd1 vccd1 net1220 sky130_fd_sc_hd__buf_4
XFILLER_0_79_1020 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1231 net1233 vssd1 vssd1 vccd1 vccd1 net1231 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07706__A net1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10188_ _03460_ _06029_ vssd1 vssd1 vccd1 vccd1 _06030_ sky130_fd_sc_hd__nand2_1
Xfanout1242 net1243 vssd1 vssd1 vccd1 vccd1 net1242 sky130_fd_sc_hd__buf_4
Xfanout1253 net1264 vssd1 vssd1 vccd1 vccd1 net1253 sky130_fd_sc_hd__buf_4
Xfanout1264 net1278 vssd1 vssd1 vccd1 vccd1 net1264 sky130_fd_sc_hd__clkbuf_2
XANTENNA__06915__A2 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_14__f_wb_clk_i_X clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout1275 net1277 vssd1 vssd1 vccd1 vccd1 net1275 sky130_fd_sc_hd__buf_4
Xfanout1286 net1302 vssd1 vssd1 vccd1 vccd1 net1286 sky130_fd_sc_hd__clkbuf_4
X_14996_ clknet_leaf_64_wb_clk_i net44 _01361_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[15\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1297 net1301 vssd1 vssd1 vccd1 vccd1 net1297 sky130_fd_sc_hd__buf_4
XANTENNA__08117__A1 net1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_1107 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13947_ clknet_leaf_122_wb_clk_i _01711_ _00312_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[301\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09865__B2 _02804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07325__C1 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11662__S net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09882__D_N net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07876__B1 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_58 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13878_ clknet_leaf_178_wb_clk_i _01642_ _00243_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[232\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10786__B net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_767 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_147_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12829_ net1388 vssd1 vssd1 vccd1 vccd1 _00593_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_173_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_916 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08971__S net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_62 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08020_ net1141 _03956_ _03960_ _03961_ vssd1 vssd1 vccd1 vccd1 _03962_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_25_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_170_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold703 team_03_WB.instance_to_wrap.core.register_file.registers_state\[361\] vssd1
+ vssd1 vccd1 vccd1 net2196 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_170_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold714 team_03_WB.instance_to_wrap.core.register_file.registers_state\[294\] vssd1
+ vssd1 vccd1 vccd1 net2207 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08053__B1 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold725 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[17\] vssd1 vssd1 vccd1
+ vccd1 net2218 sky130_fd_sc_hd__dlygate4sd3_1
Xhold736 team_03_WB.instance_to_wrap.core.register_file.registers_state\[246\] vssd1
+ vssd1 vccd1 vccd1 net2229 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold747 team_03_WB.instance_to_wrap.core.register_file.registers_state\[906\] vssd1
+ vssd1 vccd1 vccd1 net2240 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold758 team_03_WB.instance_to_wrap.core.register_file.registers_state\[506\] vssd1
+ vssd1 vccd1 vccd1 net2251 sky130_fd_sc_hd__dlygate4sd3_1
X_09971_ _03205_ net661 vssd1 vssd1 vccd1 vccd1 _05890_ sky130_fd_sc_hd__nor2_1
XFILLER_0_110_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold769 team_03_WB.instance_to_wrap.core.register_file.registers_state\[575\] vssd1
+ vssd1 vccd1 vccd1 net2262 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07319__C net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10026__B net99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13618__A net1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08922_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[43\] net977
+ vssd1 vssd1 vccd1 vccd1 _04864_ sky130_fd_sc_hd__or2_1
XANTENNA__09148__A3 _04119_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08356__A1 net1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_51_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08356__B2 net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08853_ net1056 team_03_WB.instance_to_wrap.core.register_file.registers_state\[576\]
+ net1009 team_03_WB.instance_to_wrap.core.register_file.registers_state\[608\] net946
+ vssd1 vssd1 vccd1 vccd1 _04795_ sky130_fd_sc_hd__a221o_1
XANTENNA__11360__B1 net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11138__A net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07804_ net1097 team_03_WB.instance_to_wrap.core.register_file.registers_state\[203\]
+ net797 team_03_WB.instance_to_wrap.core.register_file.registers_state\[235\] net730
+ vssd1 vssd1 vccd1 vccd1 _03746_ sky130_fd_sc_hd__a221o_1
X_08784_ _04724_ _04725_ net868 vssd1 vssd1 vccd1 vccd1 _04726_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08108__A1 net1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_140_3243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07735_ team_03_WB.instance_to_wrap.core.decoder.inst\[23\] _03672_ _03674_ _03676_
+ net718 vssd1 vssd1 vccd1 vccd1 _03677_ sky130_fd_sc_hd__a41o_1
XANTENNA__11112__A0 net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_140_3254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08203__S1 net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout457_A net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1199_A net1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07867__B1 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07666_ net1174 team_03_WB.instance_to_wrap.core.register_file.registers_state\[190\]
+ net888 net1127 vssd1 vssd1 vccd1 vccd1 _03608_ sky130_fd_sc_hd__a211o_1
XFILLER_0_94_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_49_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09405_ _05164_ _05340_ _05345_ net582 vssd1 vssd1 vccd1 vccd1 _05347_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_49_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07597_ net1112 team_03_WB.instance_to_wrap.core.register_file.registers_state\[377\]
+ net902 vssd1 vssd1 vccd1 vccd1 _03539_ sky130_fd_sc_hd__or3_1
XANTENNA_fanout624_A net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1366_A net1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09977__S net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_759 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09336_ _05235_ _05275_ _05277_ vssd1 vssd1 vccd1 vccd1 _05278_ sky130_fd_sc_hd__a21o_2
XANTENNA__10983__Y _06561_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09267_ _05207_ _05208_ vssd1 vssd1 vccd1 vccd1 _05209_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_106_815 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout412_X net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_768 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1154_X net1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09278__A _04893_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08218_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[433\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[401\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[305\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[273\]
+ net961 net1071 vssd1 vssd1 vccd1 vccd1 _04160_ sky130_fd_sc_hd__mux4_1
XFILLER_0_65_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09198_ net565 _05134_ _05139_ vssd1 vssd1 vccd1 vccd1 _05140_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout993_A net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08149_ net936 _04089_ _04090_ vssd1 vssd1 vccd1 vccd1 _04091_ sky130_fd_sc_hd__o21a_1
XFILLER_0_43_492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_1916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10926__A0 _06513_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_1927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11160_ net651 _06657_ vssd1 vssd1 vccd1 vccd1 _06658_ sky130_fd_sc_hd__and2_1
XANTENNA__07229__C net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout781_X net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_2666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout879_X net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_2677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10111_ _04807_ net660 vssd1 vssd1 vccd1 vccd1 _05955_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_8_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10651__S net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11091_ net834 net272 vssd1 vssd1 vccd1 vccd1 _06622_ sky130_fd_sc_hd__and2_2
XTAP_TAPCELL_ROW_164_3733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_164_3744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08347__A1 net1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10042_ net15 net1040 _05906_ net2736 vssd1 vssd1 vccd1 vccd1 _02689_ sky130_fd_sc_hd__a22o_1
Xhold30 team_03_WB.instance_to_wrap.core.register_file.registers_state\[983\] vssd1
+ vssd1 vccd1 vccd1 net1523 sky130_fd_sc_hd__dlygate4sd3_1
Xhold41 team_03_WB.instance_to_wrap.core.register_file.registers_state\[939\] vssd1
+ vssd1 vccd1 vccd1 net1534 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07555__C1 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14850_ clknet_leaf_81_wb_clk_i net1674 _01215_ vssd1 vssd1 vccd1 vccd1 net105 sky130_fd_sc_hd__dfrtp_1
Xhold52 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[3\] vssd1 vssd1 vccd1
+ vccd1 net1545 sky130_fd_sc_hd__dlygate4sd3_1
Xhold63 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[19\] vssd1 vssd1 vccd1
+ vccd1 net1556 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold74 team_03_WB.instance_to_wrap.core.register_file.registers_state\[19\] vssd1
+ vssd1 vccd1 vccd1 net1567 sky130_fd_sc_hd__dlygate4sd3_1
Xhold85 team_03_WB.instance_to_wrap.core.ru.state\[1\] vssd1 vssd1 vccd1 vccd1 net1578
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13801_ clknet_leaf_72_wb_clk_i _01565_ _00166_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[155\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold96 team_03_WB.instance_to_wrap.core.register_file.registers_state\[20\] vssd1
+ vssd1 vccd1 vccd1 net1589 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14781_ clknet_leaf_89_wb_clk_i _02545_ _01146_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_I\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input18_A DAT_I[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11993_ net298 net2603 net445 vssd1 vssd1 vccd1 vccd1 _01551_ sky130_fd_sc_hd__mux2_1
XANTENNA__13263__A net1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13732_ clknet_leaf_28_wb_clk_i _01496_ _00097_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[86\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_168_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07858__B1 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10944_ net508 net597 net265 net520 net1820 vssd1 vssd1 vccd1 vccd1 _02312_ sky130_fd_sc_hd__a32o_1
XFILLER_0_97_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07322__A2 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13663_ clknet_leaf_21_wb_clk_i _01427_ _00028_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_10875_ net691 net315 net585 vssd1 vssd1 vccd1 vccd1 _06472_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_112_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_231 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12614_ net1299 vssd1 vssd1 vccd1 vccd1 _00378_ sky130_fd_sc_hd__inv_2
XFILLER_0_155_247 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08807__C1 net1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13594_ net1268 vssd1 vssd1 vccd1 vccd1 _01358_ sky130_fd_sc_hd__inv_2
XFILLER_0_94_882 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_85_wb_clk_i clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_85_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_109_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07086__A1 net1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12545_ net1272 vssd1 vssd1 vccd1 vccd1 _00309_ sky130_fd_sc_hd__inv_2
XFILLER_0_170_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_152_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_14_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_14_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_124_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_431 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12476_ net1414 vssd1 vssd1 vccd1 vccd1 _00240_ sky130_fd_sc_hd__inv_2
XANTENNA__07200__S net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14215_ clknet_leaf_99_wb_clk_i _01979_ _00580_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[569\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08035__B1 net1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_5 team_03_WB.instance_to_wrap.core.decoder.inst\[23\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_11427_ net639 net708 _06463_ vssd1 vssd1 vccd1 vccd1 _06756_ sky130_fd_sc_hd__and3_4
XFILLER_0_22_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10917__B1 net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07389__A2 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09916__A _02837_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09783__B1 _04816_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14146_ clknet_leaf_175_wb_clk_i _01910_ _00511_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[500\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_104_380 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11358_ net493 net622 _06731_ net400 net2088 vssd1 vssd1 vccd1 vccd1 _02101_ sky130_fd_sc_hd__a32o_1
XFILLER_0_1_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11590__A0 _06477_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07794__C1 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11657__S net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10309_ team_03_WB.instance_to_wrap.core.pc.current_pc\[27\] _06150_ vssd1 vssd1
+ vccd1 vccd1 _06151_ sky130_fd_sc_hd__and2_1
X_14077_ clknet_leaf_26_wb_clk_i _01841_ _00442_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[431\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11289_ net1249 net838 _06536_ net671 vssd1 vssd1 vccd1 vccd1 _06712_ sky130_fd_sc_hd__and4_1
XPHY_EDGE_ROW_5_Left_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13028_ net1366 vssd1 vssd1 vccd1 vccd1 _00792_ sky130_fd_sc_hd__inv_2
XANTENNA__11342__B1 net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1050 net1055 vssd1 vssd1 vccd1 vccd1 net1050 sky130_fd_sc_hd__clkbuf_4
Xfanout1061 net1062 vssd1 vssd1 vccd1 vccd1 net1061 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_83_13 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11893__A1 net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1072 net1073 vssd1 vssd1 vccd1 vccd1 net1072 sky130_fd_sc_hd__buf_4
XANTENNA__08966__S net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1083 net1093 vssd1 vssd1 vccd1 vccd1 net1083 sky130_fd_sc_hd__buf_2
Xfanout1094 net1095 vssd1 vssd1 vccd1 vccd1 net1094 sky130_fd_sc_hd__buf_2
XFILLER_0_83_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10797__A net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14979_ clknet_leaf_87_wb_clk_i _02731_ _01344_ vssd1 vssd1 vccd1 vccd1 net231 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_117_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07520_ net1102 team_03_WB.instance_to_wrap.core.register_file.registers_state\[966\]
+ net800 team_03_WB.instance_to_wrap.core.register_file.registers_state\[998\] net1134
+ vssd1 vssd1 vccd1 vccd1 _03462_ sky130_fd_sc_hd__a221o_1
XFILLER_0_18_1132 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08510__A1 net1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_704 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_575 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07451_ net1184 team_03_WB.instance_to_wrap.core.register_file.registers_state\[53\]
+ net876 vssd1 vssd1 vccd1 vccd1 _03393_ sky130_fd_sc_hd__and3_1
XFILLER_0_88_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_114 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07382_ net811 _03319_ _03320_ _03323_ vssd1 vssd1 vccd1 vccd1 _03324_ sky130_fd_sc_hd__o22a_1
XFILLER_0_57_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11124__C net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_61 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_2005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09121_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[558\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[526\]
+ net978 vssd1 vssd1 vccd1 vccd1 _05063_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_44_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10736__S net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08274__B1 net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09052_ net1047 team_03_WB.instance_to_wrap.core.register_file.registers_state\[463\]
+ net998 team_03_WB.instance_to_wrap.core.register_file.registers_state\[495\] net1073
+ vssd1 vssd1 vccd1 vccd1 _04994_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_96_2341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_96_2352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_656 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08206__S net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08003_ net613 _03943_ vssd1 vssd1 vccd1 vccd1 _03945_ sky130_fd_sc_hd__nor2_1
XANTENNA__08026__B1 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11140__B net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold500 team_03_WB.instance_to_wrap.core.register_file.registers_state\[890\] vssd1
+ vssd1 vccd1 vccd1 net1993 sky130_fd_sc_hd__dlygate4sd3_1
Xhold511 team_03_WB.instance_to_wrap.core.i_hit vssd1 vssd1 vccd1 vccd1 net2004 sky130_fd_sc_hd__dlygate4sd3_1
Xhold522 team_03_WB.instance_to_wrap.core.register_file.registers_state\[225\] vssd1
+ vssd1 vccd1 vccd1 net2015 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08577__A1 net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_974 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold533 team_03_WB.instance_to_wrap.core.register_file.registers_state\[389\] vssd1
+ vssd1 vccd1 vccd1 net2026 sky130_fd_sc_hd__dlygate4sd3_1
Xhold544 team_03_WB.instance_to_wrap.core.register_file.registers_state\[899\] vssd1
+ vssd1 vccd1 vccd1 net2037 sky130_fd_sc_hd__dlygate4sd3_1
Xhold555 team_03_WB.instance_to_wrap.core.register_file.registers_state\[569\] vssd1
+ vssd1 vccd1 vccd1 net2048 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11581__A0 net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold566 team_03_WB.instance_to_wrap.core.register_file.registers_state\[626\] vssd1
+ vssd1 vccd1 vccd1 net2059 sky130_fd_sc_hd__dlygate4sd3_1
Xhold577 team_03_WB.instance_to_wrap.core.register_file.registers_state\[277\] vssd1
+ vssd1 vccd1 vccd1 net2070 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10923__A3 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13348__A net1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold588 team_03_WB.instance_to_wrap.core.register_file.registers_state\[822\] vssd1
+ vssd1 vccd1 vccd1 net2081 sky130_fd_sc_hd__dlygate4sd3_1
X_09954_ _05881_ net1981 net291 vssd1 vssd1 vccd1 vccd1 _02750_ sky130_fd_sc_hd__mux2_1
Xhold599 team_03_WB.instance_to_wrap.core.register_file.registers_state\[170\] vssd1
+ vssd1 vccd1 vccd1 net2092 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_70_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1114_A net1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09037__S net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08905_ _04841_ _04846_ net873 vssd1 vssd1 vccd1 vccd1 _04847_ sky130_fd_sc_hd__mux2_1
XANTENNA__07346__A net1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09885_ _03137_ _04148_ vssd1 vssd1 vccd1 vccd1 _05827_ sky130_fd_sc_hd__nor2_1
Xhold1200 team_03_WB.instance_to_wrap.core.register_file.registers_state\[69\] vssd1
+ vssd1 vccd1 vccd1 net2693 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1211 team_03_WB.instance_to_wrap.core.register_file.registers_state\[648\] vssd1
+ vssd1 vccd1 vccd1 net2704 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_57_91 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08836_ net578 net353 vssd1 vssd1 vccd1 vccd1 _04778_ sky130_fd_sc_hd__nand2_2
Xhold1222 team_03_WB.instance_to_wrap.core.register_file.registers_state\[909\] vssd1
+ vssd1 vccd1 vccd1 net2715 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1233 team_03_WB.instance_to_wrap.core.register_file.registers_state\[709\] vssd1
+ vssd1 vccd1 vccd1 net2726 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11884__A1 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1244 team_03_WB.instance_to_wrap.core.register_file.registers_state\[76\] vssd1
+ vssd1 vccd1 vccd1 net2737 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1255 team_03_WB.instance_to_wrap.core.register_file.registers_state\[349\] vssd1
+ vssd1 vccd1 vccd1 net2748 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1266 team_03_WB.instance_to_wrap.core.register_file.registers_state\[731\] vssd1
+ vssd1 vccd1 vccd1 net2759 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1277 team_03_WB.instance_to_wrap.CPU_DAT_O\[2\] vssd1 vssd1 vccd1 vccd1 net2770
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08767_ net1214 _04703_ _04705_ _04708_ vssd1 vssd1 vccd1 vccd1 _04709_ sky130_fd_sc_hd__a31o_1
Xhold1288 team_03_WB.instance_to_wrap.CPU_DAT_O\[14\] vssd1 vssd1 vccd1 vccd1 net2781
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout741_A net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout362_X net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout839_A _06386_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13083__A net1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07718_ net824 _03651_ _03654_ _03659_ net718 vssd1 vssd1 vccd1 vccd1 _03660_ sky130_fd_sc_hd__o221ai_4
XTAP_TAPCELL_ROW_68_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08698_ net1241 team_03_WB.instance_to_wrap.core.register_file.registers_state\[328\]
+ net976 team_03_WB.instance_to_wrap.core.register_file.registers_state\[360\] net1071
+ vssd1 vssd1 vccd1 vccd1 _04640_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_68_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07649_ net1192 team_03_WB.instance_to_wrap.core.register_file.registers_state\[686\]
+ vssd1 vssd1 vccd1 vccd1 _03591_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout627_X net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1369_X net1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10660_ team_03_WB.instance_to_wrap.core.control_logic.instruction\[1\] team_03_WB.instance_to_wrap.CPU_DAT_O\[1\]
+ net846 vssd1 vssd1 vccd1 vccd1 _02468_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_882 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_24_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_157_3592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09319_ net592 _05258_ vssd1 vssd1 vccd1 vccd1 _05261_ sky130_fd_sc_hd__nand2_1
XFILLER_0_134_910 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10646__S net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10591_ _06293_ _06300_ net1144 net1145 vssd1 vssd1 vccd1 vccd1 _06301_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_36_768 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12330_ net1285 vssd1 vssd1 vccd1 vccd1 _00094_ sky130_fd_sc_hd__inv_2
XFILLER_0_69_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout996_X net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_114_2717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08017__B1 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_998 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12261_ net1353 vssd1 vssd1 vccd1 vccd1 _00025_ sky130_fd_sc_hd__inv_2
XFILLER_0_32_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14000_ clknet_leaf_157_wb_clk_i _01764_ _00365_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[354\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08568__A1 net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11212_ net273 net2296 net486 vssd1 vssd1 vccd1 vccd1 _02196_ sky130_fd_sc_hd__mux2_1
X_12192_ net1646 vssd1 vssd1 vccd1 vccd1 _02361_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__08032__A3 net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07776__C1 net1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07240__A1 net1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11143_ net711 net694 net300 vssd1 vssd1 vccd1 vccd1 _06648_ sky130_fd_sc_hd__or3b_1
XFILLER_0_102_895 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07256__A net1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_132_wb_clk_i clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_132_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_11074_ net832 net278 vssd1 vssd1 vccd1 vccd1 _06615_ sky130_fd_sc_hd__and2_1
X_14902_ clknet_leaf_58_wb_clk_i _02665_ _01267_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.pc.current_pc\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_10025_ net914 vssd1 vssd1 vccd1 vccd1 _05902_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14833_ clknet_leaf_87_wb_clk_i net1838 _01198_ vssd1 vssd1 vccd1 vccd1 net154 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_99_963 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14764_ clknet_leaf_61_wb_clk_i _02528_ _01129_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_11976_ net280 net2536 net443 vssd1 vssd1 vccd1 vccd1 _01568_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13715_ clknet_leaf_102_wb_clk_i _01479_ _00080_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[69\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_38_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_168_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10927_ net693 _05718_ net586 vssd1 vssd1 vccd1 vccd1 _06514_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_58_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_169_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14695_ clknet_leaf_63_wb_clk_i _02459_ _01060_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.ADR_I\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11940__S net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13646_ clknet_leaf_124_wb_clk_i _01410_ _00011_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_156_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10858_ team_03_WB.instance_to_wrap.core.decoder.inst\[10\] _06389_ _06390_ vssd1
+ vssd1 vccd1 vccd1 _06457_ sky130_fd_sc_hd__a21o_1
XFILLER_0_73_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08256__B1 net995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13577_ net1435 vssd1 vssd1 vccd1 vccd1 _01341_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10789_ _02932_ _06391_ vssd1 vssd1 vccd1 vccd1 _06399_ sky130_fd_sc_hd__and2_4
XANTENNA__08534__B net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10063__B1 net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11241__A net1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12528_ net1402 vssd1 vssd1 vccd1 vccd1 _00292_ sky130_fd_sc_hd__inv_2
XFILLER_0_125_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12459_ net1282 vssd1 vssd1 vccd1 vccd1 _00223_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_10_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08559__A1 net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09646__A _03428_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09220__A2 _03314_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14129_ clknet_leaf_138_wb_clk_i _01893_ _00494_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[483\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07231__A1 net1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout309 _05846_ vssd1 vssd1 vccd1 vccd1 net309 sky130_fd_sc_hd__buf_2
X_06951_ team_03_WB.instance_to_wrap.core.decoder.inst\[25\] net826 vssd1 vssd1 vccd1
+ vccd1 _02893_ sky130_fd_sc_hd__nand2_2
XFILLER_0_158_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07519__C1 net1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09670_ _05187_ _05302_ _05305_ vssd1 vssd1 vccd1 vccd1 _05612_ sky130_fd_sc_hd__nand3_1
XANTENNA_clkbuf_leaf_77_wb_clk_i_A clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_06882_ team_03_WB.instance_to_wrap.core.decoder.inst\[29\] team_03_WB.instance_to_wrap.core.decoder.inst\[26\]
+ team_03_WB.instance_to_wrap.core.decoder.inst\[25\] vssd1 vssd1 vccd1 vccd1 _02824_
+ sky130_fd_sc_hd__or3_1
XANTENNA__12800__A net1402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08731__A1 net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14995__Q team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[14\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09381__A _04354_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08621_ net1068 _04561_ _04562_ vssd1 vssd1 vccd1 vccd1 _04563_ sky130_fd_sc_hd__a21o_1
XANTENNA__08709__B net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08552_ net1229 team_03_WB.instance_to_wrap.core.register_file.registers_state\[94\]
+ net955 team_03_WB.instance_to_wrap.core.register_file.registers_state\[126\] net917
+ vssd1 vssd1 vccd1 vccd1 _04494_ sky130_fd_sc_hd__o221a_1
XFILLER_0_166_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_51 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_59_Left_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07503_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[167\] net785
+ net752 _03444_ vssd1 vssd1 vccd1 vccd1 _03445_ sky130_fd_sc_hd__o211a_1
XANTENNA__07298__A1 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08483_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[955\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[923\]
+ net988 vssd1 vssd1 vccd1 vccd1 _04425_ sky130_fd_sc_hd__mux2_1
XANTENNA__11850__S net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07434_ net1177 team_03_WB.instance_to_wrap.core.register_file.registers_state\[180\]
+ vssd1 vssd1 vccd1 vccd1 _03376_ sky130_fd_sc_hd__and2_1
XFILLER_0_119_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_21_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_543 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07365_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[924\] net792
+ _03306_ vssd1 vssd1 vccd1 vccd1 _03307_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_135_3142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_863 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_3153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1064_A net1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10054__B1 net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09104_ _05044_ _05045_ net857 vssd1 vssd1 vccd1 vccd1 _05046_ sky130_fd_sc_hd__o21a_1
XFILLER_0_33_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07296_ net1158 _03235_ _03236_ net1120 vssd1 vssd1 vccd1 vccd1 _03238_ sky130_fd_sc_hd__a31o_1
XFILLER_0_33_749 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09035_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[816\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[784\]
+ net984 vssd1 vssd1 vccd1 vccd1 _04977_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_475 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1231_A net1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1329_A net1330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_760 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_68_Left_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold330 net126 vssd1 vssd1 vccd1 vccd1 net1823 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold341 team_03_WB.instance_to_wrap.core.register_file.registers_state\[562\] vssd1
+ vssd1 vccd1 vccd1 net1834 sky130_fd_sc_hd__dlygate4sd3_1
Xhold352 team_03_WB.instance_to_wrap.core.ru.state\[6\] vssd1 vssd1 vccd1 vccd1 net1845
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout691_A net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold363 _02600_ vssd1 vssd1 vccd1 vccd1 net1856 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout789_A net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold374 net220 vssd1 vssd1 vccd1 vccd1 net1867 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold385 team_03_WB.instance_to_wrap.core.register_file.registers_state\[180\] vssd1
+ vssd1 vccd1 vccd1 net1878 sky130_fd_sc_hd__dlygate4sd3_1
Xhold396 team_03_WB.instance_to_wrap.core.register_file.registers_state\[404\] vssd1
+ vssd1 vccd1 vccd1 net1889 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09990__S net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1117_X net1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout810 _02849_ vssd1 vssd1 vccd1 vccd1 net810 sky130_fd_sc_hd__clkbuf_8
XANTENNA__08970__A1 net1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout821 net825 vssd1 vssd1 vccd1 vccd1 net821 sky130_fd_sc_hd__buf_6
X_09937_ _03563_ net661 vssd1 vssd1 vccd1 vccd1 _05873_ sky130_fd_sc_hd__nor2_1
Xfanout832 _06387_ vssd1 vssd1 vccd1 vccd1 net832 sky130_fd_sc_hd__clkbuf_8
XANTENNA__10109__A1 _04770_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout843 _06304_ vssd1 vssd1 vccd1 vccd1 net843 sky130_fd_sc_hd__buf_2
XANTENNA__11306__A0 _06616_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout854 net855 vssd1 vssd1 vccd1 vccd1 net854 sky130_fd_sc_hd__buf_4
XANTENNA_fanout956_A net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout865 net866 vssd1 vssd1 vccd1 vccd1 net865 sky130_fd_sc_hd__buf_4
XFILLER_0_99_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout876 net879 vssd1 vssd1 vccd1 vccd1 net876 sky130_fd_sc_hd__clkbuf_4
X_09868_ net352 _05107_ _05809_ vssd1 vssd1 vccd1 vccd1 _05810_ sky130_fd_sc_hd__a21o_1
Xfanout887 _02845_ vssd1 vssd1 vccd1 vccd1 net887 sky130_fd_sc_hd__clkbuf_8
Xfanout898 net900 vssd1 vssd1 vccd1 vccd1 net898 sky130_fd_sc_hd__clkbuf_2
Xhold1030 team_03_WB.instance_to_wrap.core.register_file.registers_state\[484\] vssd1
+ vssd1 vccd1 vccd1 net2523 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1041 team_03_WB.instance_to_wrap.core.register_file.registers_state\[857\] vssd1
+ vssd1 vccd1 vccd1 net2534 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08183__C1 net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08819_ net1215 _04757_ _04758_ _04760_ vssd1 vssd1 vccd1 vccd1 _04761_ sky130_fd_sc_hd__a31o_1
Xhold1052 team_03_WB.instance_to_wrap.core.register_file.registers_state\[453\] vssd1
+ vssd1 vccd1 vccd1 net2545 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1063 team_03_WB.instance_to_wrap.core.register_file.registers_state\[123\] vssd1
+ vssd1 vccd1 vccd1 net2556 sky130_fd_sc_hd__dlygate4sd3_1
X_09799_ _03489_ _04591_ vssd1 vssd1 vccd1 vccd1 _05741_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout744_X net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1074 team_03_WB.instance_to_wrap.core.register_file.registers_state\[647\] vssd1
+ vssd1 vccd1 vccd1 net2567 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1085 team_03_WB.instance_to_wrap.core.register_file.registers_state\[637\] vssd1
+ vssd1 vccd1 vccd1 net2578 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_107_2565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07930__C1 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07082__Y _03024_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_2576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11830_ _06665_ net456 net323 net2057 vssd1 vssd1 vccd1 vccd1 _01709_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_77_Left_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1096 team_03_WB.instance_to_wrap.core.register_file.registers_state\[728\] vssd1
+ vssd1 vccd1 vccd1 net2589 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10230__A net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_159_3632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_159_3643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07289__A1 net1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11761_ net653 _06588_ net464 net333 net2042 vssd1 vssd1 vccd1 vccd1 _01776_ sky130_fd_sc_hd__a32o_1
XFILLER_0_166_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13500_ net1328 vssd1 vssd1 vccd1 vccd1 _01264_ sky130_fd_sc_hd__inv_2
X_10712_ net1765 net528 net523 _06346_ vssd1 vssd1 vccd1 vccd1 _02458_ sky130_fd_sc_hd__a22o_1
XANTENNA__13541__A net1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08769__A1_N net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14480_ clknet_leaf_156_wb_clk_i _02244_ _00845_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[834\]
+ sky130_fd_sc_hd__dfrtp_1
X_11692_ _06734_ net385 net341 net2550 vssd1 vssd1 vccd1 vccd1 _01842_ sky130_fd_sc_hd__a22o_1
XANTENNA__08635__A net1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13431_ net1406 vssd1 vssd1 vccd1 vccd1 _01195_ sky130_fd_sc_hd__inv_2
X_10643_ net1209 net2745 net845 vssd1 vssd1 vccd1 vccd1 _02485_ sky130_fd_sc_hd__mux2_1
XANTENNA__12034__A1 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08354__B net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11061__A net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13362_ net1319 vssd1 vssd1 vccd1 vccd1 _01126_ sky130_fd_sc_hd__inv_2
XANTENNA_input85_A wbs_adr_i[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_172_3898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10574_ net1773 net532 net599 _05884_ vssd1 vssd1 vccd1 vccd1 _02549_ sky130_fd_sc_hd__a22o_1
XFILLER_0_134_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15101_ net912 vssd1 vssd1 vccd1 vccd1 net260 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12313_ net1355 vssd1 vssd1 vccd1 vccd1 _00077_ sky130_fd_sc_hd__inv_2
XFILLER_0_121_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_86_Left_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07461__A1 net1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13293_ net1328 vssd1 vssd1 vccd1 vccd1 _01057_ sky130_fd_sc_hd__inv_2
XFILLER_0_146_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15032_ clknet_leaf_104_wb_clk_i _02752_ _01397_ vssd1 vssd1 vccd1 vccd1 net188 sky130_fd_sc_hd__dfrtp_1
X_12244_ net1815 vssd1 vssd1 vccd1 vccd1 _01413_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_111_wb_clk_i_A clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_48_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12175_ net1590 vssd1 vssd1 vccd1 vccd1 _02378_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__10405__A net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08961__A1 net1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11126_ net1247 net832 _06414_ net670 vssd1 vssd1 vccd1 vccd1 _06638_ sky130_fd_sc_hd__or4_1
XANTENNA__07417__C net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06972__B1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11935__S net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09913__B _05718_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11057_ net1043 net838 _06545_ net671 vssd1 vssd1 vccd1 vccd1 _06606_ sky130_fd_sc_hd__and4_1
XANTENNA__08174__C1 net1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08713__A1 net1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10008_ _02921_ net2194 net289 vssd1 vssd1 vccd1 vccd1 _02706_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_95_Left_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_900 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14816_ clknet_leaf_92_wb_clk_i net1722 _01181_ vssd1 vssd1 vccd1 vccd1 net167 sky130_fd_sc_hd__dfrtp_1
XANTENNA__10140__A _03390_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_153_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14747_ clknet_leaf_48_wb_clk_i _02511_ _01112_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08477__B1 net999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11959_ net632 _06736_ net465 net365 net2110 vssd1 vssd1 vccd1 vccd1 _01584_ sky130_fd_sc_hd__a32o_1
XFILLER_0_114_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11670__S net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14678_ clknet_leaf_82_wb_clk_i _02442_ _01043_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.ADR_I\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10794__B _05867_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13629_ net1422 vssd1 vssd1 vccd1 vccd1 _01393_ sky130_fd_sc_hd__inv_2
XFILLER_0_117_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12025__A1 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_938 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08229__B1 net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_15_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10036__B1 net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09977__A0 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_150_wb_clk_i_A clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_07150_ net1109 team_03_WB.instance_to_wrap.core.register_file.registers_state\[320\]
+ net1155 vssd1 vssd1 vccd1 vccd1 _03092_ sky130_fd_sc_hd__a21o_1
XFILLER_0_42_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10587__B2 _03059_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07988__C1 net1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07452__A1 net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07081_ net718 _03006_ _03015_ _03022_ vssd1 vssd1 vccd1 vccd1 _03023_ sky130_fd_sc_hd__o22a_4
XFILLER_0_30_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_140_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_130_3050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12073__Y _06819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07167__Y _03109_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07204__A1 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_1144 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11000__A2 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08401__B1 net1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12006__S net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07983_ net823 _03914_ _03924_ vssd1 vssd1 vccd1 vccd1 _03925_ sky130_fd_sc_hd__o21ai_1
XANTENNA__11845__S net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09722_ _05216_ _05662_ _05221_ vssd1 vssd1 vccd1 vccd1 _05664_ sky130_fd_sc_hd__o21ai_1
X_06934_ net823 _02875_ net724 vssd1 vssd1 vccd1 vccd1 _02876_ sky130_fd_sc_hd__a21o_1
XANTENNA__08165__C1 net1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09901__B1 _05833_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09653_ net352 _05587_ _05594_ vssd1 vssd1 vccd1 vccd1 _05595_ sky130_fd_sc_hd__a21oi_2
XTAP_TAPCELL_ROW_87_2159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06865_ team_03_WB.instance_to_wrap.core.control_logic.instruction\[3\] team_03_WB.instance_to_wrap.core.control_logic.instruction\[2\]
+ team_03_WB.instance_to_wrap.core.control_logic.instruction\[1\] team_03_WB.instance_to_wrap.core.control_logic.instruction\[0\]
+ vssd1 vssd1 vccd1 vccd1 _02807_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_59_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout272_A _06483_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08604_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[869\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[837\]
+ net992 vssd1 vssd1 vccd1 vccd1 _04546_ sky130_fd_sc_hd__mux2_1
XANTENNA__11146__A net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09584_ _05525_ vssd1 vssd1 vccd1 vccd1 _05526_ sky130_fd_sc_hd__inv_2
XFILLER_0_167_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_26_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_26_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_118_Right_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_167_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08535_ _04476_ vssd1 vssd1 vccd1 vccd1 _04477_ sky130_fd_sc_hd__inv_2
XFILLER_0_166_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10275__A0 _04444_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11580__S net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1181_A net1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1279_A net1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_2462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15124__1489 vssd1 vssd1 vccd1 vccd1 _15124__1489/HI net1489 sky130_fd_sc_hd__conb_1
XFILLER_0_159_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08466_ net859 _04404_ _04407_ vssd1 vssd1 vccd1 vccd1 _04408_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_102_2473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_147_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07417_ net1175 team_03_WB.instance_to_wrap.core.register_file.registers_state\[692\]
+ net880 vssd1 vssd1 vccd1 vccd1 _03359_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_154_3540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08397_ net1223 _04337_ _04338_ vssd1 vssd1 vccd1 vccd1 _04339_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout704_A net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout325_X net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09968__A0 _05888_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_800 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1067_X net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09985__S net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07348_ net811 _03285_ _03286_ _03289_ vssd1 vssd1 vccd1 vccd1 _03290_ sky130_fd_sc_hd__o22a_1
XANTENNA__10578__B2 _05888_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11775__B1 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_150_3448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_150_3459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07279_ net1108 team_03_WB.instance_to_wrap.core.register_file.registers_state\[649\]
+ net804 team_03_WB.instance_to_wrap.core.register_file.registers_state\[681\] net734
+ vssd1 vssd1 vccd1 vccd1 _03221_ sky130_fd_sc_hd__a221o_1
XFILLER_0_27_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1234_X net1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09286__A _04922_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09018_ net1242 team_03_WB.instance_to_wrap.core.register_file.registers_state\[176\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[144\] net984 net928
+ vssd1 vssd1 vccd1 vccd1 _04960_ sky130_fd_sc_hd__a221o_1
X_10290_ _05963_ _06128_ _06130_ net303 net304 vssd1 vssd1 vccd1 vccd1 _06132_ sky130_fd_sc_hd__a32o_1
XANTENNA__08190__A net1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout694_X net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold160 net235 vssd1 vssd1 vccd1 vccd1 net1653 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07518__B net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold171 team_03_WB.instance_to_wrap.core.register_file.registers_state\[814\] vssd1
+ vssd1 vccd1 vccd1 net1664 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1401_X net1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold182 team_03_WB.instance_to_wrap.core.register_file.registers_state\[989\] vssd1
+ vssd1 vccd1 vccd1 net1675 sky130_fd_sc_hd__dlygate4sd3_1
Xhold193 net131 vssd1 vssd1 vccd1 vccd1 net1686 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08943__A1 net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout861_X net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout640 net641 vssd1 vssd1 vccd1 vccd1 net640 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_109_2605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout959_X net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout651 net652 vssd1 vssd1 vccd1 vccd1 net651 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_109_2616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout662 net663 vssd1 vssd1 vccd1 vccd1 net662 sky130_fd_sc_hd__buf_2
X_13980_ clknet_leaf_146_wb_clk_i _01744_ _00345_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[334\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout673 net674 vssd1 vssd1 vccd1 vccd1 net673 sky130_fd_sc_hd__clkbuf_4
Xfanout684 _03278_ vssd1 vssd1 vccd1 vccd1 net684 sky130_fd_sc_hd__buf_4
XANTENNA__08156__C1 net1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout695 net696 vssd1 vssd1 vccd1 vccd1 net695 sky130_fd_sc_hd__clkbuf_4
X_12931_ net1356 vssd1 vssd1 vccd1 vccd1 _00695_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_126_2963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07903__C1 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12862_ net1414 vssd1 vssd1 vccd1 vccd1 _00626_ sky130_fd_sc_hd__inv_2
XFILLER_0_34_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14601_ clknet_leaf_78_wb_clk_i _02365_ _00966_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[955\]
+ sky130_fd_sc_hd__dfstp_1
X_11813_ net646 _06640_ net451 net323 net1802 vssd1 vssd1 vccd1 vccd1 _01726_ sky130_fd_sc_hd__a32o_1
XANTENNA__11058__A2 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12793_ net1359 vssd1 vssd1 vccd1 vccd1 _00557_ sky130_fd_sc_hd__inv_2
XFILLER_0_96_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_819 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11490__S net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14532_ clknet_leaf_23_wb_clk_i _02296_ _00897_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[886\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_174_3938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11744_ _06565_ net453 net331 net2410 vssd1 vssd1 vccd1 vccd1 _01793_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_174_3949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07131__B1 net1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08365__A net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14463_ clknet_leaf_166_wb_clk_i _02227_ _00828_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[817\]
+ sky130_fd_sc_hd__dfrtp_1
X_11675_ net2581 _06633_ net344 vssd1 vssd1 vccd1 vccd1 _01858_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_12_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08306__S0 net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13414_ net1428 vssd1 vssd1 vccd1 vccd1 _01178_ sky130_fd_sc_hd__inv_2
XFILLER_0_36_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10626_ net1545 team_03_WB.instance_to_wrap.CPU_DAT_O\[3\] net842 vssd1 vssd1 vccd1
+ vccd1 _02502_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_118 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input88_X net88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14394_ clknet_leaf_143_wb_clk_i _02158_ _00759_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[748\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_153_367 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11766__B1 net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10569__B2 _05879_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13345_ net1319 vssd1 vssd1 vccd1 vccd1 _01109_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10557_ net1758 net531 net598 _05861_ vssd1 vssd1 vccd1 vccd1 _02566_ sky130_fd_sc_hd__a22o_1
XFILLER_0_84_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09908__B _05583_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12615__A net1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13276_ net1423 vssd1 vssd1 vccd1 vccd1 _01040_ sky130_fd_sc_hd__inv_2
XFILLER_0_122_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11518__A0 net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10488_ net112 net1027 net905 net1742 vssd1 vssd1 vccd1 vccd1 _02621_ sky130_fd_sc_hd__a22o_1
X_15015_ clknet_leaf_104_wb_clk_i _02735_ _01380_ vssd1 vssd1 vccd1 vccd1 net202 sky130_fd_sc_hd__dfrtp_1
X_12227_ net1589 vssd1 vssd1 vccd1 vccd1 _01430_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__09924__A net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12158_ net1575 vssd1 vssd1 vccd1 vccd1 _02395_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__11665__S net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11109_ net265 net2761 net418 vssd1 vssd1 vccd1 vccd1 _02248_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_1075 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12089_ net639 _06656_ net474 net442 net2102 vssd1 vssd1 vccd1 vccd1 _01458_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_34_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07444__A net1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08698__B1 net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07163__B _03104_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08974__S net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_2056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_752 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_2067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08320_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[568\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[536\]
+ net985 vssd1 vssd1 vccd1 vccd1 _04262_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_375 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08251_ _04187_ _04192_ net871 vssd1 vssd1 vccd1 vccd1 _04193_ sky130_fd_sc_hd__mux2_1
XANTENNA__11413__B _06751_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07673__A1 net1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08870__B1 _04770_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10009__A0 _02888_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07202_ net1170 team_03_WB.instance_to_wrap.core.register_file.registers_state\[210\]
+ net756 team_03_WB.instance_to_wrap.core.register_file.registers_state\[242\] net740
+ vssd1 vssd1 vccd1 vccd1 _03144_ sky130_fd_sc_hd__o221a_1
XFILLER_0_144_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08182_ net935 _04122_ _04123_ vssd1 vssd1 vccd1 vccd1 _04124_ sky130_fd_sc_hd__o21a_1
XFILLER_0_172_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_171_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10029__B net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_395 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11757__B1 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08848__S1 net1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07133_ net1140 _03074_ net719 vssd1 vssd1 vccd1 vccd1 _03075_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_43_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11221__A2 net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07064_ _02998_ _02999_ _03004_ _03005_ net1119 net1139 vssd1 vssd1 vccd1 vccd1 _03006_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__07619__A net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput210 net210 vssd1 vssd1 vccd1 vccd1 gpio_out[13] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_12_Right_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11509__A0 _06505_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput221 net221 vssd1 vssd1 vccd1 vccd1 gpio_out[24] sky130_fd_sc_hd__buf_2
XFILLER_0_112_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_58_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput232 net232 vssd1 vssd1 vccd1 vccd1 gpio_out[35] sky130_fd_sc_hd__buf_2
Xoutput243 net243 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[13] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_58_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput254 net254 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[28] sky130_fd_sc_hd__buf_2
XANTENNA_fanout1027_A net1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10732__A1 _05646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06985__D_N team_03_WB.instance_to_wrap.core.decoder.inst\[14\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout487_A _06680_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07966_ net1193 team_03_WB.instance_to_wrap.core.register_file.registers_state\[176\]
+ net903 net1132 vssd1 vssd1 vccd1 vccd1 _03908_ sky130_fd_sc_hd__a211o_1
XANTENNA__09025__S1 net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09705_ _05646_ vssd1 vssd1 vccd1 vccd1 _05647_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06917_ net1106 team_03_WB.instance_to_wrap.core.register_file.registers_state\[68\]
+ net804 team_03_WB.instance_to_wrap.core.register_file.registers_state\[100\] net750
+ vssd1 vssd1 vccd1 vccd1 _02859_ sky130_fd_sc_hd__a221o_1
XANTENNA__11288__A2 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07897_ net1200 team_03_WB.instance_to_wrap.core.register_file.registers_state\[431\]
+ net877 _02870_ vssd1 vssd1 vccd1 vccd1 _03839_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout275_X net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout654_A net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1396_A net1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10496__B1 net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09636_ net568 _05486_ vssd1 vssd1 vccd1 vccd1 _05578_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_104_2502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06848_ net1241 vssd1 vssd1 vccd1 vccd1 _02791_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_104_2513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_21_Right_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07361__B1 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10986__Y _06564_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_404 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07900__A2 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09567_ _03904_ _04235_ _04816_ vssd1 vssd1 vccd1 vccd1 _05509_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout442_X net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout821_A net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10248__A0 _04294_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1184_X net1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_2860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout919_A net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08518_ _04456_ _04457_ _04459_ _04458_ net916 net859 vssd1 vssd1 vccd1 vccd1 _04460_
+ sky130_fd_sc_hd__mux4_1
X_09498_ _04448_ _04534_ net559 vssd1 vssd1 vccd1 vccd1 _05440_ sky130_fd_sc_hd__mux2_1
XANTENNA__08185__A net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09653__A2 _05587_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10799__A1 team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[30\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11996__A0 _06509_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_147_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08449_ net933 _04389_ _04390_ net854 vssd1 vssd1 vccd1 vccd1 _04391_ sky130_fd_sc_hd__o211a_1
XFILLER_0_53_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08861__B1 net1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11460__A2 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout707_X net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_939 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xwire315 _05611_ vssd1 vssd1 vccd1 vccd1 net315 sky130_fd_sc_hd__buf_2
XFILLER_0_34_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11460_ net514 net642 _06585_ net394 net2227 vssd1 vssd1 vccd1 vccd1 _02034_ sky130_fd_sc_hd__a32o_1
XFILLER_0_18_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_490 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11748__B1 net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10411_ _06002_ _06004_ _06068_ vssd1 vssd1 vccd1 vccd1 _06235_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_45_192 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10507__X _06286_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_326 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08613__B1 net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10654__S net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11391_ net1249 net839 _06545_ net669 vssd1 vssd1 vccd1 vccd1 _06748_ sky130_fd_sc_hd__and4_1
XPHY_EDGE_ROW_30_Right_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13130_ net1284 vssd1 vssd1 vccd1 vccd1 _00894_ sky130_fd_sc_hd__inv_2
X_10342_ team_03_WB.instance_to_wrap.core.pc.current_pc\[24\] _06148_ team_03_WB.instance_to_wrap.core.pc.current_pc\[25\]
+ vssd1 vssd1 vccd1 vccd1 _06178_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_131_540 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13061_ net1348 vssd1 vssd1 vccd1 vccd1 _00825_ sky130_fd_sc_hd__inv_2
X_10273_ _04070_ _06113_ vssd1 vssd1 vccd1 vccd1 _06115_ sky130_fd_sc_hd__xor2_2
XFILLER_0_44_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12012_ _06761_ net475 net361 net2556 vssd1 vssd1 vccd1 vccd1 _01533_ sky130_fd_sc_hd__a22o_1
XFILLER_0_40_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input48_A gpio_in[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1402 net1408 vssd1 vssd1 vccd1 vccd1 net1402 sky130_fd_sc_hd__buf_4
XANTENNA__11920__A0 _06454_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1413 net1436 vssd1 vssd1 vccd1 vccd1 net1413 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_167_3797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1424 net1425 vssd1 vssd1 vccd1 vccd1 net1424 sky130_fd_sc_hd__buf_4
Xclkbuf_leaf_39_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_39_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xfanout1435 net1436 vssd1 vssd1 vccd1 vccd1 net1435 sky130_fd_sc_hd__buf_2
XANTENNA__13266__A net1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout470 net471 vssd1 vssd1 vccd1 vccd1 net470 sky130_fd_sc_hd__buf_2
Xfanout481 _06800_ vssd1 vssd1 vccd1 vccd1 net481 sky130_fd_sc_hd__buf_4
XANTENNA__07264__A team_03_WB.instance_to_wrap.core.decoder.inst\[28\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout492 net517 vssd1 vssd1 vccd1 vccd1 net492 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_45_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13963_ clknet_leaf_38_wb_clk_i _01727_ _00328_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[317\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10487__B1 net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12914_ net1338 vssd1 vssd1 vccd1 vccd1 _00678_ sky130_fd_sc_hd__inv_2
X_13894_ clknet_leaf_27_wb_clk_i _01658_ _00259_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[248\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_115_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_17_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12845_ net1293 vssd1 vssd1 vccd1 vccd1 _00609_ sky130_fd_sc_hd__inv_2
XFILLER_0_115_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_17_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_139_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12776_ net1291 vssd1 vssd1 vccd1 vccd1 _00540_ sky130_fd_sc_hd__inv_2
XANTENNA__11987__A0 _06468_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07104__B1 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08301__C1 net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_14_Left_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_166_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14515_ clknet_leaf_100_wb_clk_i _02279_ _00880_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[869\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_3_0_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11727_ net2153 _06487_ net337 vssd1 vssd1 vccd1 vccd1 _01809_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08852__B1 net1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11451__A2 net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_991 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09919__A _03351_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11658_ net2036 _06479_ net342 vssd1 vssd1 vccd1 vccd1 _01875_ sky130_fd_sc_hd__mux2_1
X_14446_ clknet_leaf_126_wb_clk_i _02210_ _00811_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[800\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10609_ net1828 team_03_WB.instance_to_wrap.CPU_DAT_O\[20\] net840 vssd1 vssd1 vccd1
+ vccd1 _02519_ sky130_fd_sc_hd__mux2_1
XANTENNA__07407__A1 net1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_738 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14377_ clknet_leaf_117_wb_clk_i _02141_ _00742_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[731\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_141_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11589_ net273 net2392 net447 vssd1 vssd1 vccd1 vccd1 _01940_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold907 team_03_WB.instance_to_wrap.core.register_file.registers_state\[921\] vssd1
+ vssd1 vccd1 vccd1 net2400 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13328_ net1325 vssd1 vssd1 vccd1 vccd1 _01092_ sky130_fd_sc_hd__inv_2
Xhold918 team_03_WB.instance_to_wrap.core.register_file.registers_state\[917\] vssd1
+ vssd1 vccd1 vccd1 net2411 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07439__A net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11754__A3 net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold929 team_03_WB.instance_to_wrap.core.register_file.registers_state\[707\] vssd1
+ vssd1 vccd1 vccd1 net2422 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10962__A1 team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[2\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13259_ net1287 vssd1 vssd1 vccd1 vccd1 _01023_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_36_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08907__A1 net1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08368__C1 net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_23_Left_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06918__B1 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08383__A2 net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13176__A net1380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07820_ net1177 team_03_WB.instance_to_wrap.core.register_file.registers_state\[138\]
+ vssd1 vssd1 vccd1 vccd1 _03762_ sky130_fd_sc_hd__or2_1
XFILLER_0_19_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07591__B1 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07018__S0 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07751_ net1098 team_03_WB.instance_to_wrap.core.register_file.registers_state\[364\]
+ net897 vssd1 vssd1 vccd1 vccd1 _03693_ sky130_fd_sc_hd__or3_1
XANTENNA__07605__C net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10478__B1 net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07682_ net1114 _03622_ _03623_ vssd1 vssd1 vccd1 vccd1 _03624_ sky130_fd_sc_hd__or3_1
X_09421_ net1019 net826 team_03_WB.instance_to_wrap.core.decoder.inst\[31\] vssd1
+ vssd1 vccd1 vccd1 _05363_ sky130_fd_sc_hd__o21a_1
XFILLER_0_35_83 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11690__A2 net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08518__S0 net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11424__A _06517_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09352_ _04178_ _05292_ vssd1 vssd1 vccd1 vccd1 _05294_ sky130_fd_sc_hd__nor2_2
XFILLER_0_164_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11978__A0 net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08209__S net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08303_ _04241_ _04244_ net872 vssd1 vssd1 vccd1 vccd1 _04245_ sky130_fd_sc_hd__a21o_1
XFILLER_0_164_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_158_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_142_51 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07646__A1 net1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11143__B net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09283_ _03243_ _05224_ vssd1 vssd1 vccd1 vccd1 _05225_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07340__C net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11442__A2 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08843__B1 net1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_532 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08234_ net1081 _04175_ vssd1 vssd1 vccd1 vccd1 _04176_ sky130_fd_sc_hd__nand2_1
XANTENNA__06952__S net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08165_ _04104_ _04105_ _04106_ net935 net1217 vssd1 vssd1 vccd1 vccd1 _04107_ sky130_fd_sc_hd__a221o_1
XFILLER_0_16_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout402_A _06718_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_160_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_151 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10402__B1 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07116_ net824 _03049_ _03052_ _03057_ vssd1 vssd1 vccd1 vccd1 _03058_ sky130_fd_sc_hd__a22o_2
XFILLER_0_15_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08096_ net1173 team_03_WB.instance_to_wrap.core.register_file.registers_state\[90\]
+ net759 team_03_WB.instance_to_wrap.core.register_file.registers_state\[122\] net725
+ vssd1 vssd1 vccd1 vccd1 _04038_ sky130_fd_sc_hd__o221a_1
XFILLER_0_63_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10953__A1 _06533_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload80 clknet_leaf_27_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload80/X sky130_fd_sc_hd__clkbuf_8
X_07047_ net718 _02982_ _02988_ _02973_ vssd1 vssd1 vccd1 vccd1 _02989_ sky130_fd_sc_hd__a31oi_1
Xclkload91 clknet_leaf_73_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload91/X sky130_fd_sc_hd__clkbuf_8
XANTENNA__08359__C1 net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1409_A net1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09020__B1 net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout771_A net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout392_X net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11902__B1 net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10023__C_N net88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout869_A net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07031__C1 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_3347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_3358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08998_ net1218 _04939_ _04938_ net1210 vssd1 vssd1 vccd1 vccd1 _04940_ sky130_fd_sc_hd__o211a_1
XANTENNA__07084__A net1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07949_ net1088 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1015\]
+ net893 _03890_ net1152 vssd1 vssd1 vccd1 vccd1 _03891_ sky130_fd_sc_hd__o311a_1
XTAP_TAPCELL_ROW_3_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout657_X net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_162_3694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_170_Right_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_123_2911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10960_ _06541_ net2037 net520 vssd1 vssd1 vccd1 vccd1 _02309_ sky130_fd_sc_hd__mux2_1
XANTENNA__07334__B1 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11130__A1 net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09619_ net320 _05550_ _05560_ net321 _05557_ vssd1 vssd1 vccd1 vccd1 _05561_ sky130_fd_sc_hd__a221o_1
XANTENNA__07885__A1 net1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10891_ net313 net309 net316 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[15\]
+ vssd1 vssd1 vccd1 vccd1 _06485_ sky130_fd_sc_hd__o31a_1
XANTENNA__10649__S net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11681__A2 net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout824_X net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12630_ net1257 vssd1 vssd1 vccd1 vccd1 _00394_ sky130_fd_sc_hd__inv_2
XANTENNA_input102_A wbs_we_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_157_wb_clk_i clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_157_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__09087__B1 net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11969__B1 net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_906 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07637__A1 net1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12561_ net1270 vssd1 vssd1 vccd1 vccd1 _00325_ sky130_fd_sc_hd__inv_2
XANTENNA__11053__B net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10641__A0 net1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11512_ _06519_ net2592 net390 vssd1 vssd1 vccd1 vccd1 _01994_ sky130_fd_sc_hd__mux2_1
X_14300_ clknet_leaf_156_wb_clk_i _02064_ _00665_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[654\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_93_596 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12492_ net1311 vssd1 vssd1 vccd1 vccd1 _00256_ sky130_fd_sc_hd__inv_2
XFILLER_0_81_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14231_ clknet_leaf_115_wb_clk_i _01995_ _00596_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[585\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_62_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11443_ net656 _06570_ vssd1 vssd1 vccd1 vccd1 _06761_ sky130_fd_sc_hd__nor2_1
XANTENNA__08598__C1 net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11197__B2 net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11736__A3 net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14162_ clknet_leaf_163_wb_clk_i _01926_ _00527_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[516\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_324 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11374_ net505 net633 _06739_ net400 net1799 vssd1 vssd1 vccd1 vccd1 _02093_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_169_3837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_178 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10944__A1 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_169_3848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13113_ net1357 vssd1 vssd1 vccd1 vccd1 _00877_ sky130_fd_sc_hd__inv_2
XANTENNA__08081__C net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10325_ net282 _06152_ _06161_ net678 vssd1 vssd1 vccd1 vccd1 _06165_ sky130_fd_sc_hd__o31a_1
XANTENNA__07270__C1 net1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14093_ clknet_leaf_185_wb_clk_i _01857_ _00458_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[447\]
+ sky130_fd_sc_hd__dfrtp_1
X_13044_ net1308 vssd1 vssd1 vccd1 vccd1 _00808_ sky130_fd_sc_hd__inv_2
XANTENNA__07546__X _03488_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10256_ _06096_ _06097_ vssd1 vssd1 vccd1 vccd1 _06098_ sky130_fd_sc_hd__nand2_1
XANTENNA__09905__C _05632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1210 net1213 vssd1 vssd1 vccd1 vccd1 net1210 sky130_fd_sc_hd__buf_4
Xfanout1221 net1222 vssd1 vssd1 vccd1 vccd1 net1221 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_56_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1232 net1233 vssd1 vssd1 vccd1 vccd1 net1232 sky130_fd_sc_hd__clkbuf_4
X_10187_ _04591_ team_03_WB.instance_to_wrap.core.pc.current_pc\[6\] net675 vssd1
+ vssd1 vccd1 vccd1 _06029_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_1032 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1243 net1246 vssd1 vssd1 vccd1 vccd1 net1243 sky130_fd_sc_hd__buf_2
Xfanout1254 net1264 vssd1 vssd1 vccd1 vccd1 net1254 sky130_fd_sc_hd__clkbuf_4
Xfanout1265 net1267 vssd1 vssd1 vccd1 vccd1 net1265 sky130_fd_sc_hd__buf_4
XFILLER_0_79_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1276 net1277 vssd1 vssd1 vccd1 vccd1 net1276 sky130_fd_sc_hd__buf_2
Xfanout1287 net1289 vssd1 vssd1 vccd1 vccd1 net1287 sky130_fd_sc_hd__buf_4
X_14995_ clknet_leaf_63_wb_clk_i net43 _01360_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[14\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1298 net1301 vssd1 vssd1 vccd1 vccd1 net1298 sky130_fd_sc_hd__buf_2
XANTENNA__08748__S0 net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13946_ clknet_leaf_146_wb_clk_i _01710_ _00311_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[300\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07325__B1 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07722__A net1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13877_ clknet_leaf_129_wb_clk_i _01641_ _00242_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[231\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10786__C net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_159_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12828_ net1419 vssd1 vssd1 vccd1 vccd1 _00592_ sky130_fd_sc_hd__inv_2
XANTENNA__08825__B1 net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_619 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_928 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12759_ net1386 vssd1 vssd1 vccd1 vccd1 _00523_ sky130_fd_sc_hd__inv_2
XFILLER_0_112_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10632__A0 team_03_WB.instance_to_wrap.core.decoder.inst\[29\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08553__A net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_495 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_890 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14429_ clknet_leaf_166_wb_clk_i _02193_ _00794_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[783\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_142_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08589__C1 net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold704 team_03_WB.instance_to_wrap.core.register_file.registers_state\[336\] vssd1
+ vssd1 vccd1 vccd1 net2197 sky130_fd_sc_hd__dlygate4sd3_1
Xhold715 team_03_WB.instance_to_wrap.core.register_file.registers_state\[676\] vssd1
+ vssd1 vccd1 vccd1 net2208 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10935__A1 net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold726 team_03_WB.instance_to_wrap.core.register_file.registers_state\[809\] vssd1
+ vssd1 vccd1 vccd1 net2219 sky130_fd_sc_hd__dlygate4sd3_1
Xhold737 team_03_WB.instance_to_wrap.core.register_file.registers_state\[371\] vssd1
+ vssd1 vccd1 vccd1 net2230 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_31_Left_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_141_189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09970_ _05889_ net1771 net293 vssd1 vssd1 vccd1 vccd1 _02742_ sky130_fd_sc_hd__mux2_1
Xhold748 team_03_WB.instance_to_wrap.core.register_file.registers_state\[682\] vssd1
+ vssd1 vccd1 vccd1 net2241 sky130_fd_sc_hd__dlygate4sd3_1
Xhold759 net193 vssd1 vssd1 vccd1 vccd1 net2252 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12803__A net1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08921_ net436 net428 net591 vssd1 vssd1 vccd1 vccd1 _04863_ sky130_fd_sc_hd__nor3_1
XANTENNA__14998__Q team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[17\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09002__B1 net1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08852_ net1056 team_03_WB.instance_to_wrap.core.register_file.registers_state\[704\]
+ net1009 team_03_WB.instance_to_wrap.core.register_file.registers_state\[736\] net930
+ vssd1 vssd1 vccd1 vccd1 _04794_ sky130_fd_sc_hd__a221o_1
XANTENNA__11360__A1 net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07564__B1 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08761__C1 net1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07803_ net1097 team_03_WB.instance_to_wrap.core.register_file.registers_state\[75\]
+ net797 team_03_WB.instance_to_wrap.core.register_file.registers_state\[107\] net749
+ vssd1 vssd1 vccd1 vccd1 _03745_ sky130_fd_sc_hd__a221o_1
XFILLER_0_58_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11138__B net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08783_ net1222 _04721_ _04722_ vssd1 vssd1 vccd1 vccd1 _04725_ sky130_fd_sc_hd__nand3_1
XANTENNA__11853__S net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07734_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[909\] net798
+ _03675_ vssd1 vssd1 vccd1 vccd1 _03676_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_140_3244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07316__B1 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_140_3255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_40_Left_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07867__A1 net1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07665_ net1083 net888 team_03_WB.instance_to_wrap.core.register_file.registers_state\[158\]
+ vssd1 vssd1 vccd1 vccd1 _03607_ sky130_fd_sc_hd__o21a_1
XFILLER_0_149_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09404_ _05164_ _05340_ _05345_ vssd1 vssd1 vccd1 vccd1 _05346_ sky130_fd_sc_hd__o21ai_2
XANTENNA__11154__A net1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_49_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_49_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07596_ _03534_ _03537_ net825 vssd1 vssd1 vccd1 vccd1 _03538_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_48_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09335_ _05204_ _05209_ _05213_ vssd1 vssd1 vccd1 vccd1 _05277_ sky130_fd_sc_hd__or3_1
XFILLER_0_36_906 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1261_A net1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1359_A net1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09266_ _05041_ _05206_ vssd1 vssd1 vccd1 vccd1 _05208_ sky130_fd_sc_hd__or2_1
XFILLER_0_29_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11966__A3 net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_827 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08217_ net1233 team_03_WB.instance_to_wrap.core.register_file.registers_state\[465\]
+ net961 team_03_WB.instance_to_wrap.core.register_file.registers_state\[497\] net1211
+ vssd1 vssd1 vccd1 vccd1 _04159_ sky130_fd_sc_hd__o221a_1
XFILLER_0_90_566 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09197_ net557 _05136_ _05138_ net572 vssd1 vssd1 vccd1 vccd1 _05139_ sky130_fd_sc_hd__o211a_1
XFILLER_0_105_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout405_X net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1147_X net1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09993__S net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08148_ net1232 team_03_WB.instance_to_wrap.core.register_file.registers_state\[180\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[148\] net960 net919
+ vssd1 vssd1 vccd1 vccd1 _04090_ sky130_fd_sc_hd__a221o_1
XFILLER_0_120_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_1917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout986_A net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07252__C1 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload180 clknet_leaf_97_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload180/Y sky130_fd_sc_hd__inv_6
X_08079_ net1090 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1014\]
+ net894 _04020_ net1150 vssd1 vssd1 vccd1 vccd1 _04021_ sky130_fd_sc_hd__o311a_1
XANTENNA__12713__A net1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_112_2667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10110_ team_03_WB.instance_to_wrap.core.pc.current_pc\[0\] net660 vssd1 vssd1 vccd1
+ vccd1 _05954_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_8_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11090_ _06479_ net2141 net416 vssd1 vssd1 vccd1 vccd1 _02259_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout774_X net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_164_3734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_164_3745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10041_ net16 net1036 net909 net1806 vssd1 vssd1 vccd1 vccd1 _02690_ sky130_fd_sc_hd__o22a_1
XANTENNA__08978__S0 net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold20 team_03_WB.instance_to_wrap.core.register_file.registers_state\[934\] vssd1
+ vssd1 vccd1 vccd1 net1513 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07555__B1 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold31 team_03_WB.instance_to_wrap.core.register_file.registers_state\[963\] vssd1
+ vssd1 vccd1 vccd1 net1524 sky130_fd_sc_hd__dlygate4sd3_1
Xhold42 team_03_WB.instance_to_wrap.core.register_file.registers_state\[990\] vssd1
+ vssd1 vccd1 vccd1 net1535 sky130_fd_sc_hd__dlygate4sd3_1
Xhold53 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1023\] vssd1
+ vssd1 vccd1 vccd1 net1546 sky130_fd_sc_hd__dlygate4sd3_1
Xhold64 team_03_WB.instance_to_wrap.core.register_file.registers_state\[29\] vssd1
+ vssd1 vccd1 vccd1 net1557 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout941_X net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold75 team_03_WB.instance_to_wrap.core.register_file.registers_state\[12\] vssd1
+ vssd1 vccd1 vccd1 net1568 sky130_fd_sc_hd__dlygate4sd3_1
Xhold86 team_03_WB.instance_to_wrap.core.register_file.registers_state\[993\] vssd1
+ vssd1 vccd1 vccd1 net1579 sky130_fd_sc_hd__dlygate4sd3_1
X_13800_ clknet_leaf_6_wb_clk_i _01564_ _00165_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[154\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold97 team_03_WB.instance_to_wrap.core.register_file.registers_state\[968\] vssd1
+ vssd1 vccd1 vccd1 net1590 sky130_fd_sc_hd__dlygate4sd3_1
X_14780_ clknet_leaf_92_wb_clk_i _02544_ _01145_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_I\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_11992_ net271 net2598 net445 vssd1 vssd1 vccd1 vccd1 _01552_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09847__A2 net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09981__C_N _05082_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07858__A1 net1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10943_ net835 _06527_ vssd1 vssd1 vccd1 vccd1 _06528_ sky130_fd_sc_hd__and2_1
X_13731_ clknet_leaf_35_wb_clk_i _01495_ _00096_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[85\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_28_wb_clk_i_A clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_151_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11064__A net1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10874_ team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[18\] net307 net685 vssd1
+ vssd1 vccd1 vccd1 _06471_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_42_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13662_ clknet_leaf_118_wb_clk_i _01426_ _00027_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_156_738 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12613_ net1353 vssd1 vssd1 vccd1 vccd1 _00377_ sky130_fd_sc_hd__inv_2
XFILLER_0_38_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13593_ net1344 vssd1 vssd1 vccd1 vccd1 _01357_ sky130_fd_sc_hd__inv_2
XANTENNA__08807__B1 net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_894 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12544_ net1397 vssd1 vssd1 vccd1 vccd1 _00308_ sky130_fd_sc_hd__inv_2
XANTENNA__08902__S0 net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07086__A2 net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_235 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12475_ net1362 vssd1 vssd1 vccd1 vccd1 _00239_ sky130_fd_sc_hd__inv_2
XFILLER_0_151_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_1081 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_134 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input70_X net70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14214_ clknet_leaf_117_wb_clk_i _01978_ _00579_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[568\]
+ sky130_fd_sc_hd__dfrtp_1
X_11426_ net295 net2567 net399 vssd1 vssd1 vccd1 vccd1 _02057_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_6 net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_999 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10917__A1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_54_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_54_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__09783__A1 _03459_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14145_ clknet_leaf_177_wb_clk_i _01909_ _00510_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[499\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07243__C1 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11938__S net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11357_ net709 _06468_ net695 vssd1 vssd1 vccd1 vccd1 _06731_ sky130_fd_sc_hd__and3_1
XANTENNA__10842__S net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09916__B _05142_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08820__B net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07794__B1 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10308_ team_03_WB.instance_to_wrap.core.pc.current_pc\[26\] _06148_ _06149_ vssd1
+ vssd1 vccd1 vccd1 _06150_ sky130_fd_sc_hd__and3_1
XANTENNA__09408__S _03064_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08991__C1 net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07717__A net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14076_ clknet_leaf_146_wb_clk_i _01840_ _00441_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[430\]
+ sky130_fd_sc_hd__dfrtp_1
X_11288_ net515 net643 _06711_ net411 net2725 vssd1 vssd1 vccd1 vccd1 _02151_ sky130_fd_sc_hd__a32o_1
X_13027_ net1354 vssd1 vssd1 vccd1 vccd1 _00791_ sky130_fd_sc_hd__inv_2
XANTENNA__11239__A net1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10239_ _06004_ _06069_ _06077_ _06079_ _06075_ vssd1 vssd1 vccd1 vccd1 _06081_ sky130_fd_sc_hd__o41a_1
XANTENNA_clkbuf_leaf_67_wb_clk_i_A clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11342__A1 net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1040 _05904_ vssd1 vssd1 vccd1 vccd1 net1040 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08743__C1 net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1051 net1055 vssd1 vssd1 vccd1 vccd1 net1051 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_174_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1062 net1069 vssd1 vssd1 vccd1 vccd1 net1062 sky130_fd_sc_hd__buf_4
Xfanout1073 net1074 vssd1 vssd1 vccd1 vccd1 net1073 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_83_25 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1084 net1086 vssd1 vssd1 vccd1 vccd1 net1084 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11673__S net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1095 net1096 vssd1 vssd1 vccd1 vccd1 net1095 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_83_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14978_ clknet_leaf_87_wb_clk_i _02730_ _01343_ vssd1 vssd1 vccd1 vccd1 net230 sky130_fd_sc_hd__dfrtp_1
XANTENNA__10797__B _05429_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_159_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13929_ clknet_leaf_75_wb_clk_i _01693_ _00294_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[283\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10853__B1 net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07450_ net1089 net895 team_03_WB.instance_to_wrap.core.register_file.registers_state\[21\]
+ vssd1 vssd1 vccd1 vccd1 _03392_ sky130_fd_sc_hd__o21a_1
XFILLER_0_147_716 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_587 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07381_ net740 _03321_ _03322_ net806 vssd1 vssd1 vccd1 vccd1 _03323_ sky130_fd_sc_hd__a31o_1
XFILLER_0_8_126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11124__D net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09120_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[750\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[718\]
+ net976 vssd1 vssd1 vccd1 vccd1 _05062_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_79_2006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_106_Left_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11948__A3 net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_44_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08274__A1 net1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09051_ net1047 team_03_WB.instance_to_wrap.core.register_file.registers_state\[335\]
+ net998 team_03_WB.instance_to_wrap.core.register_file.registers_state\[367\] net1213
+ vssd1 vssd1 vccd1 vccd1 _04993_ sky130_fd_sc_hd__a221o_1
XFILLER_0_142_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_96_2342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_6_Right_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_96_2353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08002_ _03943_ vssd1 vssd1 vccd1 vccd1 _03944_ sky130_fd_sc_hd__inv_2
XFILLER_0_115_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_170_774 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08026__A1 net1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11140__C net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold501 team_03_WB.instance_to_wrap.core.register_file.registers_state\[751\] vssd1
+ vssd1 vccd1 vccd1 net1994 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_430 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold512 team_03_WB.instance_to_wrap.core.register_file.registers_state\[273\] vssd1
+ vssd1 vccd1 vccd1 net2005 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold523 team_03_WB.instance_to_wrap.core.register_file.registers_state\[130\] vssd1
+ vssd1 vccd1 vccd1 net2016 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11848__S net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09774__B2 _04646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13629__A net1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold534 team_03_WB.instance_to_wrap.core.register_file.registers_state\[644\] vssd1
+ vssd1 vccd1 vccd1 net2027 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_986 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold545 team_03_WB.instance_to_wrap.core.register_file.registers_state\[763\] vssd1
+ vssd1 vccd1 vccd1 net2038 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold556 team_03_WB.instance_to_wrap.core.register_file.registers_state\[186\] vssd1
+ vssd1 vccd1 vccd1 net2049 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold567 team_03_WB.instance_to_wrap.core.register_file.registers_state\[887\] vssd1
+ vssd1 vccd1 vccd1 net2060 sky130_fd_sc_hd__dlygate4sd3_1
Xhold578 team_03_WB.instance_to_wrap.core.register_file.registers_state\[561\] vssd1
+ vssd1 vccd1 vccd1 net2071 sky130_fd_sc_hd__dlygate4sd3_1
X_09953_ _03984_ net661 vssd1 vssd1 vccd1 vccd1 _05881_ sky130_fd_sc_hd__nor2_1
Xhold589 team_03_WB.instance_to_wrap.core.register_file.registers_state\[261\] vssd1
+ vssd1 vccd1 vccd1 net2082 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_115_Left_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_70_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08904_ net1221 _04844_ _04845_ vssd1 vssd1 vccd1 vccd1 _04846_ sky130_fd_sc_hd__o21a_1
X_09884_ _05283_ _05290_ _05599_ net581 vssd1 vssd1 vccd1 vccd1 _05826_ sky130_fd_sc_hd__o31a_1
XFILLER_0_148_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1107_A net1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1201 team_03_WB.instance_to_wrap.core.register_file.registers_state\[537\] vssd1
+ vssd1 vccd1 vccd1 net2694 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_57_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08734__C1 net1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1212 team_03_WB.instance_to_wrap.core.register_file.registers_state\[541\] vssd1
+ vssd1 vccd1 vccd1 net2705 sky130_fd_sc_hd__dlygate4sd3_1
X_08835_ net584 _04775_ vssd1 vssd1 vccd1 vccd1 _04777_ sky130_fd_sc_hd__nor2_4
Xhold1223 team_03_WB.instance_to_wrap.core.register_file.registers_state\[90\] vssd1
+ vssd1 vccd1 vccd1 net2716 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1234 team_03_WB.instance_to_wrap.core.register_file.registers_state\[9\] vssd1
+ vssd1 vccd1 vccd1 net2727 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout567_A _03025_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1245 team_03_WB.instance_to_wrap.core.register_file.registers_state\[860\] vssd1
+ vssd1 vccd1 vccd1 net2738 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11583__S net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1256 team_03_WB.instance_to_wrap.core.register_file.registers_state\[602\] vssd1
+ vssd1 vccd1 vccd1 net2749 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1267 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[9\] vssd1 vssd1 vccd1
+ vccd1 net2760 sky130_fd_sc_hd__dlygate4sd3_1
X_08766_ net1221 _04706_ _04707_ net1076 vssd1 vssd1 vccd1 vccd1 _04708_ sky130_fd_sc_hd__o211a_1
XFILLER_0_169_307 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1278 team_03_WB.instance_to_wrap.core.register_file.registers_state\[776\] vssd1
+ vssd1 vccd1 vccd1 net2771 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_135_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1289 team_03_WB.instance_to_wrap.CPU_DAT_O\[3\] vssd1 vssd1 vccd1 vccd1 net2782
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07362__A net1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07717_ net818 _03656_ _03658_ vssd1 vssd1 vccd1 vccd1 _03659_ sky130_fd_sc_hd__or3_1
X_08697_ net862 _04635_ _04638_ vssd1 vssd1 vccd1 vccd1 _04639_ sky130_fd_sc_hd__o21a_1
XANTENNA__11636__A2 net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout355_X net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout734_A net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1097_X net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09988__S net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07648_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[558\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[526\]
+ net777 vssd1 vssd1 vccd1 vccd1 _03590_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_165_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout522_X net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07579_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[920\] net794
+ net1014 _03520_ vssd1 vssd1 vccd1 vccd1 _03521_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout901_A net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1264_X net1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_24_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09318_ _04808_ _04812_ _04811_ vssd1 vssd1 vccd1 vccd1 _05260_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_24_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_157_3593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07068__A2 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10590_ team_03_WB.instance_to_wrap.core.i_hit _05914_ vssd1 vssd1 vccd1 vccd1 _06300_
+ sky130_fd_sc_hd__and2b_1
XFILLER_0_63_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07301__S net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09249_ _04294_ _05189_ vssd1 vssd1 vccd1 vccd1 _05191_ sky130_fd_sc_hd__nand2_1
XFILLER_0_91_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_2707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_114_2718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12260_ net1356 vssd1 vssd1 vccd1 vccd1 _00024_ sky130_fd_sc_hd__inv_2
XFILLER_0_161_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout891_X net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11211_ _06468_ net2183 net486 vssd1 vssd1 vccd1 vccd1 _02197_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout989_X net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13539__A net1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_101_wb_clk_i_A clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_12191_ net1504 vssd1 vssd1 vccd1 vccd1 _02362_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__07776__B1 net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07537__A net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11142_ net2091 net413 _06647_ net499 vssd1 vssd1 vccd1 vccd1 _02233_ sky130_fd_sc_hd__a22o_1
XANTENNA__11059__A net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11073_ _06614_ net2421 net419 vssd1 vssd1 vccd1 vccd1 _02269_ sky130_fd_sc_hd__mux2_1
X_14901_ clknet_leaf_59_wb_clk_i _02664_ _01266_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.pc.current_pc\[30\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA_input30_A DAT_I[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10024_ _05896_ _05899_ _05900_ _05901_ vssd1 vssd1 vccd1 vccd1 net257 sky130_fd_sc_hd__or4_1
XANTENNA__11493__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08740__A2 net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14832_ clknet_leaf_90_wb_clk_i net1998 _01197_ vssd1 vssd1 vccd1 vccd1 net153 sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_172_wb_clk_i clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_172_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_144_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_99_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_101_wb_clk_i clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_101_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_53_28 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14763_ clknet_leaf_49_wb_clk_i net1752 _01128_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11627__A2 net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11975_ _06405_ net2707 net443 vssd1 vssd1 vccd1 vccd1 _01569_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10835__B1 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13714_ clknet_leaf_118_wb_clk_i _01478_ _00079_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[68\]
+ sky130_fd_sc_hd__dfrtp_1
X_10926_ _06513_ net2266 net521 vssd1 vssd1 vccd1 vccd1 _02315_ sky130_fd_sc_hd__mux2_1
X_14694_ clknet_leaf_64_wb_clk_i _02458_ _01059_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.ADR_I\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_129_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13645_ net1433 vssd1 vssd1 vccd1 vccd1 _01409_ sky130_fd_sc_hd__inv_2
X_10857_ _06380_ _06389_ vssd1 vssd1 vccd1 vccd1 _06456_ sky130_fd_sc_hd__or2_2
XANTENNA__10837__S net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_500 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11522__A _06405_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08256__A1 net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_140_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_54_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13576_ net1426 vssd1 vssd1 vccd1 vccd1 _01340_ sky130_fd_sc_hd__inv_2
X_10788_ team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[31\] team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[31\]
+ net307 vssd1 vssd1 vccd1 vccd1 _06398_ sky130_fd_sc_hd__mux2_1
XFILLER_0_143_229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10063__A1 net2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_59_Right_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08534__C _04475_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11260__B1 net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11241__B net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_1029 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12527_ net1337 vssd1 vssd1 vccd1 vccd1 _00291_ sky130_fd_sc_hd__inv_2
XFILLER_0_41_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09486__X _05428_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09927__A _03638_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12458_ net1285 vssd1 vssd1 vccd1 vccd1 _00222_ sky130_fd_sc_hd__inv_2
XFILLER_0_169_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_10_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11668__S net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11012__B1 net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11409_ net275 net2282 net397 vssd1 vssd1 vccd1 vccd1 _02071_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12389_ net1353 vssd1 vssd1 vccd1 vccd1 _00153_ sky130_fd_sc_hd__inv_2
XFILLER_0_10_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_91_2250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07231__A2 net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14128_ clknet_leaf_158_wb_clk_i _01892_ _00493_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[482\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06950_ net612 _02888_ _02890_ vssd1 vssd1 vccd1 vccd1 _02892_ sky130_fd_sc_hd__o21ai_2
X_14059_ clknet_leaf_37_wb_clk_i _01823_ _00424_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[413\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08977__S net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07519__B1 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_68_Right_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08716__C1 net1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06881_ team_03_WB.instance_to_wrap.core.decoder.inst\[14\] _02820_ vssd1 vssd1 vccd1
+ vccd1 _02823_ sky130_fd_sc_hd__and2_1
XANTENNA__11866__A2 net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08620_ net1223 _04559_ _04560_ vssd1 vssd1 vccd1 vccd1 _04562_ sky130_fd_sc_hd__and3_1
XFILLER_0_55_1108 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08551_ net1232 team_03_WB.instance_to_wrap.core.register_file.registers_state\[222\]
+ net962 team_03_WB.instance_to_wrap.core.register_file.registers_state\[254\] net936
+ vssd1 vssd1 vccd1 vccd1 _04493_ sky130_fd_sc_hd__o221a_1
XANTENNA__11618__A2 net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07502_ net1204 team_03_WB.instance_to_wrap.core.register_file.registers_state\[135\]
+ vssd1 vssd1 vccd1 vccd1 _03444_ sky130_fd_sc_hd__or2_1
XANTENNA__10826__B1 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08482_ net874 _04420_ _04423_ vssd1 vssd1 vccd1 vccd1 _04424_ sky130_fd_sc_hd__or3_1
XANTENNA__08495__A1 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_1000 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07433_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[20\] net764
+ net741 _03374_ vssd1 vssd1 vccd1 vccd1 _03375_ sky130_fd_sc_hd__a211o_1
XFILLER_0_76_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10747__S net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12528__A net1402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_77_Right_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_21_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_21_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08247__A1 net1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07364_ net1083 team_03_WB.instance_to_wrap.core.register_file.registers_state\[956\]
+ net891 net1151 vssd1 vssd1 vccd1 vccd1 _03306_ sky130_fd_sc_hd__o31a_1
XFILLER_0_134_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_135_3143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09103_ net1241 team_03_WB.instance_to_wrap.core.register_file.registers_state\[142\]
+ net976 team_03_WB.instance_to_wrap.core.register_file.registers_state\[174\] net940
+ vssd1 vssd1 vccd1 vccd1 _05045_ sky130_fd_sc_hd__o221a_1
XFILLER_0_45_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_135_3154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_875 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_62 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07455__C1 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07295_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[425\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[393\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[297\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[265\]
+ net784 net1136 vssd1 vssd1 vccd1 vccd1 _03237_ sky130_fd_sc_hd__mux4_1
XFILLER_0_60_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09034_ net944 _04974_ _04975_ net856 vssd1 vssd1 vccd1 vccd1 _04976_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout1057_A net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_152_3490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_142_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11578__S net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold320 _02620_ vssd1 vssd1 vccd1 vccd1 net1813 sky130_fd_sc_hd__dlygate4sd3_1
Xhold331 _02633_ vssd1 vssd1 vccd1 vccd1 net1824 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1224_A net1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold342 team_03_WB.instance_to_wrap.core.register_file.registers_state\[184\] vssd1
+ vssd1 vccd1 vccd1 net1835 sky130_fd_sc_hd__dlygate4sd3_1
Xhold353 net204 vssd1 vssd1 vccd1 vccd1 net1846 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08955__C1 net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold364 team_03_WB.instance_to_wrap.core.register_file.registers_state\[411\] vssd1
+ vssd1 vccd1 vccd1 net1857 sky130_fd_sc_hd__dlygate4sd3_1
Xhold375 team_03_WB.instance_to_wrap.core.register_file.registers_state\[309\] vssd1
+ vssd1 vccd1 vccd1 net1868 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout684_A _03278_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold386 team_03_WB.instance_to_wrap.core.register_file.registers_state\[50\] vssd1
+ vssd1 vccd1 vccd1 net1879 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout800 net801 vssd1 vssd1 vccd1 vccd1 net800 sky130_fd_sc_hd__clkbuf_4
Xhold397 net236 vssd1 vssd1 vccd1 vccd1 net1890 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout811 net816 vssd1 vssd1 vccd1 vccd1 net811 sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_86_Right_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_170 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09936_ _05872_ net1795 net294 vssd1 vssd1 vccd1 vccd1 _02759_ sky130_fd_sc_hd__mux2_1
Xfanout822 net825 vssd1 vssd1 vccd1 vccd1 net822 sky130_fd_sc_hd__buf_4
XANTENNA_fanout1012_X net1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout833 _06387_ vssd1 vssd1 vccd1 vccd1 net833 sky130_fd_sc_hd__buf_4
Xfanout844 net845 vssd1 vssd1 vccd1 vccd1 net844 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06981__A1 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07791__S net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout855 net858 vssd1 vssd1 vccd1 vccd1 net855 sky130_fd_sc_hd__clkbuf_8
Xfanout866 _04083_ vssd1 vssd1 vccd1 vccd1 net866 sky130_fd_sc_hd__buf_6
X_09867_ net320 _05484_ _05495_ net321 _05808_ vssd1 vssd1 vccd1 vccd1 _05809_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout472_X net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout877 net878 vssd1 vssd1 vccd1 vccd1 net877 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout851_A _04096_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1020 team_03_WB.instance_to_wrap.core.register_file.registers_state\[522\] vssd1
+ vssd1 vccd1 vccd1 net2513 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout888 net891 vssd1 vssd1 vccd1 vccd1 net888 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08183__B1 net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout899 net900 vssd1 vssd1 vccd1 vccd1 net899 sky130_fd_sc_hd__buf_2
Xhold1031 team_03_WB.instance_to_wrap.core.register_file.registers_state\[288\] vssd1
+ vssd1 vccd1 vccd1 net2524 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1042 team_03_WB.instance_to_wrap.core.register_file.registers_state\[772\] vssd1
+ vssd1 vccd1 vccd1 net2535 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10070__X _05914_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08818_ net1221 _04756_ _04759_ net1076 vssd1 vssd1 vccd1 vccd1 _04760_ sky130_fd_sc_hd__o211a_1
Xhold1053 team_03_WB.instance_to_wrap.core.register_file.registers_state\[593\] vssd1
+ vssd1 vccd1 vccd1 net2546 sky130_fd_sc_hd__dlygate4sd3_1
X_09798_ net580 _05739_ net353 vssd1 vssd1 vccd1 vccd1 _05740_ sky130_fd_sc_hd__o21a_1
Xhold1064 team_03_WB.instance_to_wrap.core.register_file.registers_state\[216\] vssd1
+ vssd1 vccd1 vccd1 net2557 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1075 team_03_WB.instance_to_wrap.core.register_file.registers_state\[107\] vssd1
+ vssd1 vccd1 vccd1 net2568 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07930__B1 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_2566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1086 team_03_WB.instance_to_wrap.core.register_file.registers_state\[500\] vssd1
+ vssd1 vccd1 vccd1 net2579 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_107_2577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1097 team_03_WB.instance_to_wrap.core.register_file.registers_state\[126\] vssd1
+ vssd1 vccd1 vccd1 net2590 sky130_fd_sc_hd__dlygate4sd3_1
X_08749_ net1221 _04688_ _04689_ vssd1 vssd1 vccd1 vccd1 _04691_ sky130_fd_sc_hd__and3_1
XANTENNA__10230__B net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1381_X net1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout737_X net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10817__A0 net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_159_3633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11760_ _06587_ net462 net332 net2319 vssd1 vssd1 vccd1 vccd1 _01777_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_159_3644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_166_833 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10711_ _02771_ _05499_ net603 vssd1 vssd1 vccd1 vccd1 _06346_ sky130_fd_sc_hd__mux2_1
XANTENNA__07820__A net1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_95_Right_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10657__S net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout904_X net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11691_ _06733_ net379 net338 net2155 vssd1 vssd1 vccd1 vccd1 _01843_ sky130_fd_sc_hd__a22o_1
XFILLER_0_165_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12438__A net1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_153_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13430_ net1432 vssd1 vssd1 vccd1 vccd1 _01194_ sky130_fd_sc_hd__inv_2
X_10642_ team_03_WB.instance_to_wrap.core.decoder.inst\[19\] team_03_WB.instance_to_wrap.CPU_DAT_O\[19\]
+ net845 vssd1 vssd1 vccd1 vccd1 _02486_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_900 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09986__A1 net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13361_ net1325 vssd1 vssd1 vccd1 vccd1 _01125_ sky130_fd_sc_hd__inv_2
XANTENNA__11242__B1 net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_5_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11061__B net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10573_ net1746 net534 net601 net587 vssd1 vssd1 vccd1 vccd1 _02550_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_172_3899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_514 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15100_ net912 vssd1 vssd1 vccd1 vccd1 net259 sky130_fd_sc_hd__clkbuf_1
XANTENNA__11793__A1 _06623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12312_ net1379 vssd1 vssd1 vccd1 vccd1 _00076_ sky130_fd_sc_hd__inv_2
X_13292_ net1322 vssd1 vssd1 vccd1 vccd1 _01056_ sky130_fd_sc_hd__inv_2
XFILLER_0_134_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input78_A wbs_adr_i[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15031_ clknet_leaf_91_wb_clk_i _02751_ _01396_ vssd1 vssd1 vccd1 vccd1 net187 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_146_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12243_ net1665 vssd1 vssd1 vccd1 vccd1 _01414_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07749__B1 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11545__B2 net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07267__A net1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08946__C1 net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12174_ net1512 vssd1 vssd1 vccd1 vccd1 _02379_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11125_ net2243 net412 _06637_ net498 vssd1 vssd1 vccd1 vccd1 _02240_ sky130_fd_sc_hd__a22o_1
XANTENNA__06972__A1 net1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11056_ net2318 net422 _06605_ net510 vssd1 vssd1 vccd1 vccd1 _02277_ sky130_fd_sc_hd__a22o_1
XANTENNA__09913__C _05697_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11076__X _06616_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10007_ _03488_ net2017 net287 vssd1 vssd1 vccd1 vccd1 _02707_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_49 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08098__A net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10520__A2 net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14815_ clknet_leaf_100_wb_clk_i net1726 _01180_ vssd1 vssd1 vccd1 vccd1 net166 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08477__A1 net1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14746_ clknet_leaf_31_wb_clk_i _02510_ _01111_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11958_ net630 _06735_ net461 net364 net2280 vssd1 vssd1 vccd1 vccd1 _01585_ sky130_fd_sc_hd__a32o_1
XFILLER_0_169_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10909_ net297 net2402 net520 vssd1 vssd1 vccd1 vccd1 _02318_ sky130_fd_sc_hd__mux2_1
XANTENNA__07685__C1 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14677_ clknet_leaf_85_wb_clk_i _02441_ _01042_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.ADR_I\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_11889_ net618 _06698_ net451 net371 net2221 vssd1 vssd1 vccd1 vccd1 _01652_ sky130_fd_sc_hd__a32o_1
XFILLER_0_129_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08229__A1 net1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13628_ net1417 vssd1 vssd1 vccd1 vccd1 _01392_ sky130_fd_sc_hd__inv_2
XFILLER_0_172_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11233__A0 net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07437__C1 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13559_ net1428 vssd1 vssd1 vccd1 vccd1 _01323_ sky130_fd_sc_hd__inv_2
XFILLER_0_125_752 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10587__A2 net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07080_ net824 _03021_ net723 vssd1 vssd1 vccd1 vccd1 _03022_ sky130_fd_sc_hd__a21o_1
XFILLER_0_152_571 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07452__A2 net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_130_3040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07448__Y _03390_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_3051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11032__C_N net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_1156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_30 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07982_ net819 _03919_ _03921_ _03923_ net719 vssd1 vssd1 vccd1 vccd1 _03924_ sky130_fd_sc_hd__o41a_1
XANTENNA__12811__A net1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06963__A1 net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09392__A _04382_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09721_ _05216_ _05221_ _05662_ vssd1 vssd1 vccd1 vccd1 _05663_ sky130_fd_sc_hd__or3_1
X_06933_ net1120 _02873_ _02874_ vssd1 vssd1 vccd1 vccd1 _02875_ sky130_fd_sc_hd__a21o_1
XANTENNA__07905__A net1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11427__A net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09652_ _05513_ _05545_ _05550_ net321 _05593_ vssd1 vssd1 vccd1 vccd1 _05594_ sky130_fd_sc_hd__a221o_1
X_06864_ team_03_WB.instance_to_wrap.core.control_logic.instruction\[3\] team_03_WB.instance_to_wrap.core.control_logic.instruction\[2\]
+ team_03_WB.instance_to_wrap.core.control_logic.instruction\[1\] team_03_WB.instance_to_wrap.core.control_logic.instruction\[0\]
+ vssd1 vssd1 vccd1 vccd1 _02806_ sky130_fd_sc_hd__and4bb_1
XANTENNA__10511__A2 net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08603_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[805\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[773\]
+ net993 vssd1 vssd1 vccd1 vccd1 _04545_ sky130_fd_sc_hd__mux2_1
X_09583_ net554 _05095_ _05524_ vssd1 vssd1 vccd1 vccd1 _05525_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_145_62 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11146__B net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11861__S net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout265_A _06528_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08534_ net431 net426 _04475_ vssd1 vssd1 vccd1 vccd1 _04476_ sky130_fd_sc_hd__or3_4
XTAP_TAPCELL_ROW_26_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08468__A1 net1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10985__B net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08465_ net854 _04405_ _04406_ vssd1 vssd1 vccd1 vccd1 _04407_ sky130_fd_sc_hd__or3_1
XFILLER_0_92_403 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_2463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout432_A net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10814__A3 net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_2474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1174_A net1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11162__A net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07416_ net1175 team_03_WB.instance_to_wrap.core.register_file.registers_state\[564\]
+ net880 vssd1 vssd1 vccd1 vccd1 _03358_ sky130_fd_sc_hd__and3_1
XFILLER_0_135_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_154_3530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08396_ net1067 _04335_ _04336_ vssd1 vssd1 vccd1 vccd1 _04338_ sky130_fd_sc_hd__or3_1
XANTENNA__12016__A2 net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_154_3541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07691__A2 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_174_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07347_ net739 _03287_ _03288_ net806 vssd1 vssd1 vccd1 vccd1 _03289_ sky130_fd_sc_hd__a31o_1
XFILLER_0_61_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_163_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1341_A net1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10578__A2 net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout318_X net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07979__B1 _02869_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_150_3449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07278_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[553\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[521\]
+ net784 vssd1 vssd1 vccd1 vccd1 _03220_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout899_A net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09017_ net944 _04958_ vssd1 vssd1 vccd1 vccd1 _04959_ sky130_fd_sc_hd__or2_1
XANTENNA__11101__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1227_X net1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11527__B2 net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold150 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[10\] vssd1 vssd1 vccd1
+ vccd1 net1643 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07087__A net1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold161 team_03_WB.instance_to_wrap.ADR_I\[10\] vssd1 vssd1 vccd1 vccd1 net1654 sky130_fd_sc_hd__dlygate4sd3_1
Xhold172 team_03_WB.instance_to_wrap.core.register_file.registers_state\[4\] vssd1
+ vssd1 vccd1 vccd1 net1665 sky130_fd_sc_hd__dlygate4sd3_1
Xhold183 team_03_WB.instance_to_wrap.ADR_I\[22\] vssd1 vssd1 vccd1 vccd1 net1676 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout687_X net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold194 team_03_WB.instance_to_wrap.core.register_file.registers_state\[954\] vssd1
+ vssd1 vccd1 vccd1 net1687 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07600__C1 net1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout630 net631 vssd1 vssd1 vccd1 vccd1 net630 sky130_fd_sc_hd__clkbuf_4
Xfanout641 _06458_ vssd1 vssd1 vccd1 vccd1 net641 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_109_2606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09919_ _03351_ net661 vssd1 vssd1 vccd1 vccd1 _05861_ sky130_fd_sc_hd__nor2_1
Xfanout652 net659 vssd1 vssd1 vccd1 vccd1 net652 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_109_2617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout663 _05860_ vssd1 vssd1 vccd1 vccd1 net663 sky130_fd_sc_hd__buf_6
Xfanout674 _05948_ vssd1 vssd1 vccd1 vccd1 net674 sky130_fd_sc_hd__buf_2
XANTENNA_fanout854_X net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08156__B1 net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout685 net687 vssd1 vssd1 vccd1 vccd1 net685 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11337__A net1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout696 _06561_ vssd1 vssd1 vccd1 vccd1 net696 sky130_fd_sc_hd__clkbuf_8
X_12930_ net1360 vssd1 vssd1 vccd1 vccd1 _00694_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_126_2953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10502__A2 net1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07903__B1 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12861_ net1388 vssd1 vssd1 vccd1 vccd1 _00625_ sky130_fd_sc_hd__inv_2
XANTENNA__09105__C1 net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14600_ clknet_leaf_10_wb_clk_i _02364_ _00965_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[954\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_96_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11812_ _06639_ net458 net324 net1805 vssd1 vssd1 vccd1 vccd1 _01727_ sky130_fd_sc_hd__a22o_1
X_12792_ net1376 vssd1 vssd1 vccd1 vccd1 _00556_ sky130_fd_sc_hd__inv_2
XANTENNA__10895__B net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07550__A net1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14531_ clknet_leaf_46_wb_clk_i _02295_ _00896_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[885\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11463__B1 net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11743_ net1248 net702 _06803_ vssd1 vssd1 vccd1 vccd1 _06809_ sky130_fd_sc_hd__or3_4
XTAP_TAPCELL_ROW_174_3939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07131__A1 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11072__A net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_154_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14462_ clknet_leaf_119_wb_clk_i _02226_ _00827_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[816\]
+ sky130_fd_sc_hd__dfrtp_1
X_11674_ net2307 _06632_ net345 vssd1 vssd1 vccd1 vccd1 _01859_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_12_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11215__A0 net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13413_ net1433 vssd1 vssd1 vccd1 vccd1 _01177_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_12_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08306__S1 net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10625_ net1631 team_03_WB.instance_to_wrap.CPU_DAT_O\[4\] net842 vssd1 vssd1 vccd1
+ vccd1 _02503_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_503 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14393_ clknet_leaf_155_wb_clk_i _02157_ _00758_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[747\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10569__A2 net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_379 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10556_ team_03_WB.instance_to_wrap.core.ru.state\[5\] _06292_ net1145 vssd1 vssd1
+ vccd1 vccd1 _06299_ sky130_fd_sc_hd__and3b_4
X_13344_ net1342 vssd1 vssd1 vccd1 vccd1 _01108_ sky130_fd_sc_hd__inv_2
XANTENNA__08631__A1 net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10487_ net1688 net1027 net905 net1642 vssd1 vssd1 vccd1 vccd1 _02622_ sky130_fd_sc_hd__a22o_1
X_13275_ net1404 vssd1 vssd1 vccd1 vccd1 _01039_ sky130_fd_sc_hd__inv_2
XFILLER_0_122_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09764__X _05706_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15014_ clknet_leaf_101_wb_clk_i _02734_ _01379_ vssd1 vssd1 vccd1 vccd1 net201 sky130_fd_sc_hd__dfrtp_1
X_12226_ net1598 vssd1 vssd1 vccd1 vccd1 _01431_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__07428__C net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12157_ net1531 vssd1 vssd1 vccd1 vccd1 _02396_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__10741__A2 net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11108_ _06629_ net2677 net419 vssd1 vssd1 vccd1 vccd1 _02249_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12088_ _06788_ net462 net439 net1928 vssd1 vssd1 vccd1 vccd1 _01459_ sky130_fd_sc_hd__a22o_1
XANTENNA__08320__S net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_34_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11247__A net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11039_ net490 net646 _06595_ net420 net2112 vssd1 vssd1 vccd1 vccd1 _02284_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_34_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08698__A1 net1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13462__A net1328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_2057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_764 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_82_2068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14729_ clknet_leaf_49_wb_clk_i _02493_ _01094_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.decoder.inst\[26\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__11454__B1 net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08250_ net1218 _04190_ _04191_ vssd1 vssd1 vccd1 vccd1 _04192_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_172_600 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_173 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11206__A0 _06434_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07201_ net1170 team_03_WB.instance_to_wrap.core.register_file.registers_state\[82\]
+ net756 team_03_WB.instance_to_wrap.core.register_file.registers_state\[114\] net725
+ vssd1 vssd1 vccd1 vccd1 _03143_ sky130_fd_sc_hd__o221a_1
XFILLER_0_171_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_171_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08181_ net1230 team_03_WB.instance_to_wrap.core.register_file.registers_state\[179\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[147\] net959 net918
+ vssd1 vssd1 vccd1 vccd1 _04123_ sky130_fd_sc_hd__a221o_1
XFILLER_0_131_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_171_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12806__A net1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11757__A1 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_9_wb_clk_i clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_9_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_54_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07132_ net1118 _03068_ _03069_ _03070_ _03073_ vssd1 vssd1 vccd1 vccd1 _03074_ sky130_fd_sc_hd__a32o_1
XFILLER_0_171_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07063_ _03000_ _03001_ net749 vssd1 vssd1 vccd1 vccd1 _03005_ sky130_fd_sc_hd__mux2_1
XANTENNA__07976__A3 net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput200 net200 vssd1 vssd1 vccd1 vccd1 gpio_oeb[35] sky130_fd_sc_hd__buf_2
Xoutput211 net211 vssd1 vssd1 vccd1 vccd1 gpio_out[14] sky130_fd_sc_hd__clkbuf_4
Xoutput222 net222 vssd1 vssd1 vccd1 vccd1 gpio_out[25] sky130_fd_sc_hd__buf_2
XFILLER_0_11_731 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput233 net233 vssd1 vssd1 vccd1 vccd1 gpio_out[5] sky130_fd_sc_hd__buf_2
XFILLER_0_112_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_58_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput244 net244 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[15] sky130_fd_sc_hd__buf_2
XFILLER_0_112_276 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput255 net255 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[2] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_151_Right_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11856__S net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10193__B1 _02893_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07194__X _03136_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07965_ net1107 net903 team_03_WB.instance_to_wrap.core.register_file.registers_state\[144\]
+ vssd1 vssd1 vccd1 vccd1 _03907_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout382_A net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09704_ net582 _05636_ _05637_ _05645_ vssd1 vssd1 vccd1 vccd1 _05646_ sky130_fd_sc_hd__a31o_4
XANTENNA__11157__A net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06916_ _02855_ _02857_ net808 vssd1 vssd1 vccd1 vccd1 _02858_ sky130_fd_sc_hd__o21a_1
X_07896_ _03835_ _03837_ net1117 vssd1 vssd1 vccd1 vccd1 _03838_ sky130_fd_sc_hd__a21o_1
X_09635_ net569 _05487_ _05576_ vssd1 vssd1 vccd1 vccd1 _05577_ sky130_fd_sc_hd__a21boi_2
XANTENNA__11693__B1 net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_2503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06847_ net1222 vssd1 vssd1 vccd1 vccd1 _02790_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_104_2514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07361__A1 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1291_A net1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10996__A net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout268_X net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout647_A net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08737__Y _04679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11591__S net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1389_A net1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_416 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09638__B1 net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09566_ net580 _04477_ _05125_ _05507_ vssd1 vssd1 vccd1 vccd1 _05508_ sky130_fd_sc_hd__a31o_1
XFILLER_0_78_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09102__A2 net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_2861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08517_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[1023\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[991\]
+ net952 vssd1 vssd1 vccd1 vccd1 _04459_ sky130_fd_sc_hd__mux2_1
XANTENNA__11445__B1 net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09497_ net564 net554 _04478_ vssd1 vssd1 vccd1 vccd1 _05439_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout814_A net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1177_X net1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10000__S net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08448_ net1045 team_03_WB.instance_to_wrap.core.register_file.registers_state\[668\]
+ net996 team_03_WB.instance_to_wrap.core.register_file.registers_state\[700\] net917
+ vssd1 vssd1 vccd1 vccd1 _04390_ sky130_fd_sc_hd__a221o_1
XFILLER_0_81_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_148_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08379_ _04317_ _04318_ _04320_ _04319_ net937 net866 vssd1 vssd1 vccd1 vccd1 _04321_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_46_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10410_ _06002_ _06004_ _06068_ vssd1 vssd1 vccd1 vccd1 _06234_ sky130_fd_sc_hd__or3_1
XANTENNA__09297__A _04619_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11390_ net507 net635 _06747_ net402 net1966 vssd1 vssd1 vccd1 vccd1 _02085_ sky130_fd_sc_hd__a32o_1
XFILLER_0_150_338 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10341_ team_03_WB.instance_to_wrap.core.pc.current_pc\[26\] _06177_ net679 vssd1
+ vssd1 vccd1 vccd1 _02660_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13060_ net1367 vssd1 vssd1 vccd1 vccd1 _00824_ sky130_fd_sc_hd__inv_2
X_10272_ _04070_ _06113_ vssd1 vssd1 vccd1 vccd1 _06114_ sky130_fd_sc_hd__and2b_1
XFILLER_0_143_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12011_ net619 _06569_ net452 net359 net2150 vssd1 vssd1 vccd1 vccd1 _01534_ sky130_fd_sc_hd__a32o_1
XANTENNA__07816__Y _03758_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1403 net1408 vssd1 vssd1 vccd1 vccd1 net1403 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_167_3798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1414 net1418 vssd1 vssd1 vccd1 vccd1 net1414 sky130_fd_sc_hd__buf_4
Xfanout1425 net1426 vssd1 vssd1 vccd1 vccd1 net1425 sky130_fd_sc_hd__buf_2
Xfanout1436 net1437 vssd1 vssd1 vccd1 vccd1 net1436 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08129__A0 _04069_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout460 net463 vssd1 vssd1 vccd1 vccd1 net460 sky130_fd_sc_hd__buf_4
Xfanout471 net472 vssd1 vssd1 vccd1 vccd1 net471 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07264__B net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout482 _06779_ vssd1 vssd1 vccd1 vccd1 net482 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_6_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout493 net496 vssd1 vssd1 vccd1 vccd1 net493 sky130_fd_sc_hd__clkbuf_4
X_13962_ clknet_leaf_2_wb_clk_i _01726_ _00327_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[316\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09182__D _03104_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_79_wb_clk_i clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_79_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_12913_ net1277 vssd1 vssd1 vccd1 vccd1 _00677_ sky130_fd_sc_hd__inv_2
XFILLER_0_88_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11684__B1 net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13893_ clknet_leaf_11_wb_clk_i _01657_ _00258_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[247\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12844_ net1314 vssd1 vssd1 vccd1 vccd1 _00608_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_17_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_17_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12775_ net1363 vssd1 vssd1 vccd1 vccd1 _00539_ sky130_fd_sc_hd__inv_2
XANTENNA__08301__B1 net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14514_ clknet_leaf_164_wb_clk_i _02278_ _00879_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[868\]
+ sky130_fd_sc_hd__dfrtp_1
X_11726_ net2494 _06483_ net336 vssd1 vssd1 vccd1 vccd1 _01810_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_847 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14445_ clknet_leaf_190_wb_clk_i _02209_ _00810_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[799\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09919__B net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11657_ net2729 _06621_ net342 vssd1 vssd1 vccd1 vccd1 _01876_ sky130_fd_sc_hd__mux2_1
XANTENNA__11739__A1 net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_171 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10608_ net1619 team_03_WB.instance_to_wrap.CPU_DAT_O\[21\] net840 vssd1 vssd1 vccd1
+ vccd1 _02520_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14376_ clknet_leaf_10_wb_clk_i _02140_ _00741_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[730\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09801__B1 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11588_ _06468_ net2214 net447 vssd1 vssd1 vccd1 vccd1 _01941_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_141_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_675 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13327_ net1317 vssd1 vssd1 vccd1 vccd1 _01091_ sky130_fd_sc_hd__inv_2
Xhold908 team_03_WB.instance_to_wrap.core.register_file.registers_state\[117\] vssd1
+ vssd1 vccd1 vccd1 net2401 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10146__A _03109_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold919 team_03_WB.instance_to_wrap.core.register_file.registers_state\[344\] vssd1
+ vssd1 vccd1 vccd1 net2412 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10539_ net136 net1034 net1026 net1818 vssd1 vssd1 vccd1 vccd1 _02571_ sky130_fd_sc_hd__a22o_1
XFILLER_0_110_703 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09494__X _05436_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09935__A _04069_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13258_ net1284 vssd1 vssd1 vccd1 vccd1 _01022_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_36_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08368__B1 net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_36_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_47 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13457__A net1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12209_ net1513 vssd1 vssd1 vccd1 vccd1 _02344_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__12361__A net1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13189_ net1348 vssd1 vssd1 vccd1 vccd1 _00953_ sky130_fd_sc_hd__inv_2
XANTENNA__06918__A1 net1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10714__A2 net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07040__B1 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08383__A3 _04323_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07750_ _03688_ _03691_ net809 _03687_ vssd1 vssd1 vccd1 vccd1 _03692_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__07018__S1 net1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07681_ net1174 team_03_WB.instance_to_wrap.core.register_file.registers_state\[606\]
+ net761 team_03_WB.instance_to_wrap.core.register_file.registers_state\[638\] net727
+ vssd1 vssd1 vccd1 vccd1 _03623_ sky130_fd_sc_hd__o221a_1
XFILLER_0_56_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07343__A1 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09420_ _02782_ _02804_ net664 _05342_ vssd1 vssd1 vccd1 vccd1 _05362_ sky130_fd_sc_hd__o22a_1
XFILLER_0_35_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_149_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09351_ _04178_ _05292_ vssd1 vssd1 vccd1 vccd1 _05293_ sky130_fd_sc_hd__nand2_1
XANTENNA__08518__S1 net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11424__B _06751_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_712 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08302_ net855 _04242_ _04243_ vssd1 vssd1 vccd1 vccd1 _04244_ sky130_fd_sc_hd__or3_1
X_09282_ _03208_ _05146_ _02937_ vssd1 vssd1 vccd1 vccd1 _05224_ sky130_fd_sc_hd__o21a_1
XFILLER_0_118_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_63 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_918 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_650 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08233_ net1217 _04174_ _04173_ vssd1 vssd1 vccd1 vccd1 _04175_ sky130_fd_sc_hd__o21ai_1
XANTENNA__10650__A1 team_03_WB.instance_to_wrap.CPU_DAT_O\[11\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10755__S net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11440__A net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10982__C net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08164_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[692\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[660\]
+ net959 vssd1 vssd1 vccd1 vccd1 _04106_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08225__S net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10402__A1 net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07115_ net815 _03054_ _03056_ net818 vssd1 vssd1 vccd1 vccd1 _03057_ sky130_fd_sc_hd__o31a_1
XFILLER_0_42_163 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07949__A3 net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07803__C1 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08095_ _04034_ _04036_ net811 vssd1 vssd1 vccd1 vccd1 _04037_ sky130_fd_sc_hd__a21o_1
XFILLER_0_141_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkload70 clknet_leaf_50_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload70/X sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout1137_A _02785_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07046_ _02986_ _02987_ net824 vssd1 vssd1 vccd1 vccd1 _02988_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_30_347 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload81 clknet_leaf_28_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload81/X sky130_fd_sc_hd__clkbuf_4
Xclkload92 clknet_leaf_60_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload92/Y sky130_fd_sc_hd__inv_8
XANTENNA__08359__B1 net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_149_3440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11586__S net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13367__A net1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09020__A1 net1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1304_A net1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09056__S net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11902__A1 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_3348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_145_3359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08997_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[938\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[906\]
+ net955 vssd1 vssd1 vccd1 vccd1 _04939_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout764_A net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout385_X net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07582__A1 net1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07948_ net1181 team_03_WB.instance_to_wrap.core.register_file.registers_state\[983\]
+ vssd1 vssd1 vccd1 vccd1 _03890_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_3_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_162_3695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout931_A net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout552_X net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07334__A1 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07879_ net724 _03806_ _03812_ _03820_ vssd1 vssd1 vccd1 vccd1 _03821_ sky130_fd_sc_hd__a22oi_4
XANTENNA_clkbuf_leaf_18_wb_clk_i_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11130__A2 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07371__Y _03313_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09618_ net564 _05469_ _05558_ _05559_ vssd1 vssd1 vccd1 vccd1 _05560_ sky130_fd_sc_hd__a22o_1
XFILLER_0_168_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10890_ net693 _05646_ net585 vssd1 vssd1 vccd1 vccd1 _06484_ sky130_fd_sc_hd__o21a_1
XFILLER_0_78_550 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11418__A0 net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09549_ _03529_ _04267_ net664 _05490_ vssd1 vssd1 vccd1 vccd1 _05491_ sky130_fd_sc_hd__a22o_1
XANTENNA__09087__A1 net1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout817_X net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11969__A1 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12560_ net1403 vssd1 vssd1 vccd1 vccd1 _00324_ sky130_fd_sc_hd__inv_2
XANTENNA__12091__B1 net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11053__C _06536_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_203 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11511_ _06628_ net2691 net391 vssd1 vssd1 vccd1 vccd1 _01995_ sky130_fd_sc_hd__mux2_1
X_12491_ net1282 vssd1 vssd1 vccd1 vccd1 _00255_ sky130_fd_sc_hd__inv_2
XFILLER_0_110_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14230_ clknet_leaf_151_wb_clk_i _01994_ _00595_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[584\]
+ sky130_fd_sc_hd__dfrtp_1
X_11442_ net491 net619 _06569_ net392 net2209 vssd1 vssd1 vccd1 vccd1 _02046_ sky130_fd_sc_hd__a32o_1
Xclkbuf_leaf_126_wb_clk_i clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_126_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_163_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08598__B1 net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11197__A2 net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14161_ clknet_leaf_143_wb_clk_i _01925_ _00526_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[515\]
+ sky130_fd_sc_hd__dfrtp_1
X_11373_ net710 _06504_ net698 vssd1 vssd1 vccd1 vccd1 _06739_ sky130_fd_sc_hd__and3_1
XFILLER_0_104_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_169_3838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10944__A2 net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_169_3849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10324_ _06162_ _06163_ net283 vssd1 vssd1 vccd1 vccd1 _06164_ sky130_fd_sc_hd__a21bo_1
X_13112_ net1380 vssd1 vssd1 vccd1 vccd1 _00876_ sky130_fd_sc_hd__inv_2
XANTENNA_input60_A gpio_in[35] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14092_ clknet_leaf_16_wb_clk_i _01856_ _00457_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[446\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_131_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11496__S net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10255_ _03901_ _06095_ vssd1 vssd1 vccd1 vccd1 _06097_ sky130_fd_sc_hd__or2_1
X_13043_ net1267 vssd1 vssd1 vccd1 vccd1 _00807_ sky130_fd_sc_hd__inv_2
XANTENNA__09011__A1 net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_57_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout1200 net1201 vssd1 vssd1 vccd1 vccd1 net1200 sky130_fd_sc_hd__clkbuf_4
Xfanout1211 net1213 vssd1 vssd1 vccd1 vccd1 net1211 sky130_fd_sc_hd__buf_2
X_10186_ _06026_ _06027_ vssd1 vssd1 vccd1 vccd1 _06028_ sky130_fd_sc_hd__nor2_1
Xfanout1222 net1224 vssd1 vssd1 vccd1 vccd1 net1222 sky130_fd_sc_hd__buf_4
XANTENNA__07706__C net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1233 net1238 vssd1 vssd1 vccd1 vccd1 net1233 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_79_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1244 net1245 vssd1 vssd1 vccd1 vccd1 net1244 sky130_fd_sc_hd__clkbuf_4
Xfanout1255 net1264 vssd1 vssd1 vccd1 vccd1 net1255 sky130_fd_sc_hd__buf_4
Xfanout1266 net1267 vssd1 vssd1 vccd1 vccd1 net1266 sky130_fd_sc_hd__buf_2
Xfanout1277 net1278 vssd1 vssd1 vccd1 vccd1 net1277 sky130_fd_sc_hd__clkbuf_2
X_14994_ clknet_leaf_10_wb_clk_i net42 _01359_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[13\]
+ sky130_fd_sc_hd__dfrtp_2
Xfanout290 _05891_ vssd1 vssd1 vccd1 vccd1 net290 sky130_fd_sc_hd__buf_4
Xfanout1288 net1302 vssd1 vssd1 vccd1 vccd1 net1288 sky130_fd_sc_hd__buf_4
Xfanout1299 net1300 vssd1 vssd1 vccd1 vccd1 net1299 sky130_fd_sc_hd__buf_4
XANTENNA__08117__A3 net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08748__S1 net1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13945_ clknet_leaf_169_wb_clk_i _01709_ _00310_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[299\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09865__A3 net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07876__A2 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13876_ clknet_leaf_133_wb_clk_i _01640_ _00241_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[230\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11409__A0 net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12827_ net1296 vssd1 vssd1 vccd1 vccd1 _00591_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12082__B1 net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12758_ net1258 vssd1 vssd1 vccd1 vccd1 _00522_ sky130_fd_sc_hd__inv_2
XANTENNA__08834__A net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11709_ _06459_ _06803_ vssd1 vssd1 vccd1 vccd1 _06807_ sky130_fd_sc_hd__nor2_1
X_12689_ net1273 vssd1 vssd1 vccd1 vccd1 _00453_ sky130_fd_sc_hd__inv_2
XFILLER_0_71_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06931__S0 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14428_ clknet_leaf_151_wb_clk_i _02192_ _00793_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[782\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_96_wb_clk_i_A clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold705 team_03_WB.instance_to_wrap.core.register_file.registers_state\[873\] vssd1
+ vssd1 vccd1 vccd1 net2198 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14359_ clknet_leaf_115_wb_clk_i _02123_ _00724_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[713\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10396__B1 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08684__S0 net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold716 team_03_WB.instance_to_wrap.core.register_file.registers_state\[636\] vssd1
+ vssd1 vccd1 vccd1 net2209 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10935__A2 _05846_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold727 team_03_WB.instance_to_wrap.core.register_file.registers_state\[507\] vssd1
+ vssd1 vccd1 vccd1 net2220 sky130_fd_sc_hd__dlygate4sd3_1
Xhold738 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[11\] vssd1 vssd1 vccd1
+ vccd1 net2231 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold749 team_03_WB.instance_to_wrap.core.register_file.registers_state\[97\] vssd1
+ vssd1 vccd1 vccd1 net2242 sky130_fd_sc_hd__dlygate4sd3_1
X_08920_ net591 vssd1 vssd1 vccd1 vccd1 _04862_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13187__A net1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11896__B1 net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08851_ _04791_ _04792_ net869 vssd1 vssd1 vccd1 vccd1 _04793_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_51_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11360__A2 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08761__B1 net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07802_ _03741_ _03743_ net809 vssd1 vssd1 vccd1 vccd1 _03744_ sky130_fd_sc_hd__o21a_1
XANTENNA__11138__C net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08782_ net1066 _04723_ vssd1 vssd1 vccd1 vccd1 _04724_ sky130_fd_sc_hd__nand2_1
XFILLER_0_97_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07913__A net1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07733_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[941\] net778
+ net1014 vssd1 vssd1 vccd1 vccd1 _03675_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_140_3245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_3256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11435__A net1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07664_ net1174 team_03_WB.instance_to_wrap.core.register_file.registers_state\[62\]
+ net880 vssd1 vssd1 vccd1 vccd1 _03606_ sky130_fd_sc_hd__and3_1
X_09403_ _05343_ _05344_ vssd1 vssd1 vccd1 vccd1 _05345_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_48_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_49_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11154__B net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09069__A1 net1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07595_ net808 _03535_ _03536_ vssd1 vssd1 vccd1 vccd1 _03537_ sky130_fd_sc_hd__or3_1
XFILLER_0_153_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout345_A _06805_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1087_A net1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09334_ _05235_ _05275_ _05213_ vssd1 vssd1 vccd1 vccd1 _05276_ sky130_fd_sc_hd__a21o_1
XFILLER_0_34_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_158_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08277__C1 net1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_164_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_842 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10623__A1 team_03_WB.instance_to_wrap.CPU_DAT_O\[6\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_62_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09265_ _05041_ _05206_ vssd1 vssd1 vccd1 vccd1 _05207_ sky130_fd_sc_hd__and2_1
XANTENNA__11820__B1 net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_173_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout512_A net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1254_A net1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11170__A net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_839 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08216_ net1232 team_03_WB.instance_to_wrap.core.register_file.registers_state\[337\]
+ net961 team_03_WB.instance_to_wrap.core.register_file.registers_state\[369\] net1074
+ vssd1 vssd1 vccd1 vccd1 _04158_ sky130_fd_sc_hd__o221a_1
XFILLER_0_145_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09196_ net545 _04771_ _05137_ net561 vssd1 vssd1 vccd1 vccd1 _05138_ sky130_fd_sc_hd__a211o_1
XFILLER_0_16_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_160_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08147_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[52\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[20\]
+ net960 vssd1 vssd1 vccd1 vccd1 _04089_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout300_X net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_2760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1421_A net1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_1918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07252__B1 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkload170 clknet_leaf_86_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload170/Y sky130_fd_sc_hd__inv_8
X_08078_ net1186 team_03_WB.instance_to_wrap.core.register_file.registers_state\[982\]
+ vssd1 vssd1 vccd1 vccd1 _04020_ sky130_fd_sc_hd__or2_1
XFILLER_0_101_511 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload181 clknet_leaf_98_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload181/Y sky130_fd_sc_hd__clkinv_8
XFILLER_0_3_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout881_A net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_112_2668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07029_ _02968_ _02970_ net748 vssd1 vssd1 vccd1 vccd1 _02971_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout979_A net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_2679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_892 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_164_3735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10040_ net17 net1036 net910 net1961 vssd1 vssd1 vccd1 vccd1 _02691_ sky130_fd_sc_hd__o22a_1
XFILLER_0_11_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_164_3746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08978__S1 net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11887__B1 net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold10 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1008\] vssd1
+ vssd1 vccd1 vccd1 net1503 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07555__A1 net1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold21 team_03_WB.instance_to_wrap.core.register_file.registers_state\[959\] vssd1
+ vssd1 vccd1 vccd1 net1514 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout767_X net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold32 team_03_WB.instance_to_wrap.core.register_file.registers_state\[933\] vssd1
+ vssd1 vccd1 vccd1 net1525 sky130_fd_sc_hd__dlygate4sd3_1
Xhold43 team_03_WB.instance_to_wrap.core.register_file.registers_state\[987\] vssd1
+ vssd1 vccd1 vccd1 net1536 sky130_fd_sc_hd__dlygate4sd3_1
Xhold54 team_03_WB.instance_to_wrap.core.register_file.registers_state\[981\] vssd1
+ vssd1 vccd1 vccd1 net1547 sky130_fd_sc_hd__dlygate4sd3_1
Xhold65 team_03_WB.instance_to_wrap.core.register_file.registers_state\[996\] vssd1
+ vssd1 vccd1 vccd1 net1558 sky130_fd_sc_hd__dlygate4sd3_1
Xhold76 team_03_WB.instance_to_wrap.core.register_file.registers_state\[928\] vssd1
+ vssd1 vccd1 vccd1 net1569 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11639__B1 net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold87 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1003\] vssd1
+ vssd1 vccd1 vccd1 net1580 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout934_X net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold98 team_03_WB.instance_to_wrap.core.register_file.registers_state\[23\] vssd1
+ vssd1 vccd1 vccd1 net1591 sky130_fd_sc_hd__dlygate4sd3_1
X_11991_ net299 net2537 net446 vssd1 vssd1 vccd1 vccd1 _01553_ sky130_fd_sc_hd__mux2_1
XANTENNA__11345__A net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13730_ clknet_leaf_174_wb_clk_i _01494_ _00095_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[84\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10942_ _06524_ _06525_ _06526_ _06399_ vssd1 vssd1 vccd1 vccd1 _06527_ sky130_fd_sc_hd__o211a_4
XFILLER_0_129_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10862__A1 net1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13661_ clknet_leaf_27_wb_clk_i _01425_ _00026_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_10873_ team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[18\] net305 vssd1
+ vssd1 vccd1 vccd1 _06470_ sky130_fd_sc_hd__nand2_1
XFILLER_0_156_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12064__A0 _06519_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12612_ net1382 vssd1 vssd1 vccd1 vccd1 _00376_ sky130_fd_sc_hd__inv_2
XFILLER_0_109_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08807__A1 net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_130_wb_clk_i_A clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_13592_ net1304 vssd1 vssd1 vccd1 vccd1 _01356_ sky130_fd_sc_hd__inv_2
XFILLER_0_137_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12543_ net1350 vssd1 vssd1 vccd1 vccd1 _00307_ sky130_fd_sc_hd__inv_2
XANTENNA__08902__S1 net1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11811__B1 net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_164_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11080__A net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12474_ net1377 vssd1 vssd1 vccd1 vccd1 _00238_ sky130_fd_sc_hd__inv_2
XFILLER_0_123_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14213_ clknet_leaf_37_wb_clk_i _01977_ _00578_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[567\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_149_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_146 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11425_ net2704 net398 _06755_ net503 vssd1 vssd1 vccd1 vccd1 _02058_ sky130_fd_sc_hd__a22o_1
XFILLER_0_22_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_7 team_03_WB.instance_to_wrap.core.decoder.inst\[12\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__10917__A2 _05686_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14144_ clknet_leaf_190_wb_clk_i _01908_ _00509_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[498\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07243__B1 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09783__A2 _04619_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11356_ net495 net624 _06730_ net400 net1827 vssd1 vssd1 vccd1 vccd1 _02102_ sky130_fd_sc_hd__a32o_1
XFILLER_0_50_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09916__C _05799_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07794__A1 net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08991__B1 net995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10307_ team_03_WB.instance_to_wrap.core.pc.current_pc\[25\] team_03_WB.instance_to_wrap.core.pc.current_pc\[24\]
+ vssd1 vssd1 vccd1 vccd1 _06149_ sky130_fd_sc_hd__and2_1
X_14075_ clknet_leaf_159_wb_clk_i _01839_ _00440_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[429\]
+ sky130_fd_sc_hd__dfrtp_1
X_11287_ net715 net269 net831 vssd1 vssd1 vccd1 vccd1 _06711_ sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_94_wb_clk_i clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_94_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_13026_ net1287 vssd1 vssd1 vccd1 vccd1 _00790_ sky130_fd_sc_hd__inv_2
X_10238_ _03602_ _06073_ _06078_ vssd1 vssd1 vccd1 vccd1 _06080_ sky130_fd_sc_hd__or3_1
XANTENNA_clkbuf_4_0__f_wb_clk_i_A clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11239__B net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11878__B1 net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1030 net1035 vssd1 vssd1 vccd1 vccd1 net1030 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07546__A1 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11342__A2 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08743__B1 net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1041 _02871_ vssd1 vssd1 vccd1 vccd1 net1041 sky130_fd_sc_hd__buf_8
Xclkbuf_leaf_23_wb_clk_i clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_23_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_10169_ _04893_ net675 vssd1 vssd1 vccd1 vccd1 _06011_ sky130_fd_sc_hd__or2_1
Xfanout1052 net1055 vssd1 vssd1 vccd1 vccd1 net1052 sky130_fd_sc_hd__clkbuf_4
Xfanout1063 net1064 vssd1 vssd1 vccd1 vccd1 net1063 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08829__A _04080_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1074 _02789_ vssd1 vssd1 vccd1 vccd1 net1074 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_83_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1085 net1086 vssd1 vssd1 vccd1 vccd1 net1085 sky130_fd_sc_hd__clkbuf_4
Xfanout1096 net1105 vssd1 vssd1 vccd1 vccd1 net1096 sky130_fd_sc_hd__clkbuf_4
X_14977_ clknet_leaf_88_wb_clk_i _02729_ _01342_ vssd1 vssd1 vccd1 vccd1 net229 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11255__A net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13928_ clknet_leaf_6_wb_clk_i _01692_ _00293_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[282\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_16_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_1025 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10853__A1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13859_ clknet_leaf_34_wb_clk_i _01623_ _00224_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[213\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08835__Y _04777_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12055__A0 _06479_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07380_ net1171 team_03_WB.instance_to_wrap.core.register_file.registers_state\[223\]
+ vssd1 vssd1 vccd1 vccd1 _03322_ sky130_fd_sc_hd__or2_1
XFILLER_0_8_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10605__A1 team_03_WB.instance_to_wrap.CPU_DAT_O\[24\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_79_2007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09471__A1 net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_923 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09050_ net861 _04990_ _04991_ _04989_ vssd1 vssd1 vccd1 vccd1 _04992_ sky130_fd_sc_hd__a31o_1
XANTENNA__07482__B1 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_96_2343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_96_2354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08001_ net1219 net1015 _03107_ vssd1 vssd1 vccd1 vccd1 _03943_ sky130_fd_sc_hd__a21o_1
XANTENNA__11140__D net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_142_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold502 team_03_WB.instance_to_wrap.core.register_file.registers_state\[265\] vssd1
+ vssd1 vccd1 vccd1 net1995 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_170_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold513 team_03_WB.instance_to_wrap.core.register_file.registers_state\[409\] vssd1
+ vssd1 vccd1 vccd1 net2006 sky130_fd_sc_hd__dlygate4sd3_1
Xhold524 net207 vssd1 vssd1 vccd1 vccd1 net2017 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold535 team_03_WB.instance_to_wrap.core.register_file.registers_state\[304\] vssd1
+ vssd1 vccd1 vccd1 net2028 sky130_fd_sc_hd__dlygate4sd3_1
Xhold546 team_03_WB.instance_to_wrap.core.register_file.registers_state\[910\] vssd1
+ vssd1 vccd1 vccd1 net2039 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold557 team_03_WB.instance_to_wrap.core.register_file.registers_state\[255\] vssd1
+ vssd1 vccd1 vccd1 net2050 sky130_fd_sc_hd__dlygate4sd3_1
Xhold568 team_03_WB.instance_to_wrap.core.register_file.registers_state\[114\] vssd1
+ vssd1 vccd1 vccd1 net2061 sky130_fd_sc_hd__dlygate4sd3_1
X_09952_ _05880_ net1741 net292 vssd1 vssd1 vccd1 vccd1 _02751_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold579 team_03_WB.instance_to_wrap.core.register_file.registers_state\[884\] vssd1
+ vssd1 vccd1 vccd1 net2072 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10334__A net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08903_ net1065 _04842_ _04843_ vssd1 vssd1 vccd1 vccd1 _04845_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_70_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11869__A0 net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09883_ _05283_ _05599_ _05290_ vssd1 vssd1 vccd1 vccd1 _05825_ sky130_fd_sc_hd__o21ai_1
XANTENNA__09082__S0 net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11864__S net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout295_A _06523_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1202 team_03_WB.instance_to_wrap.core.register_file.registers_state\[835\] vssd1
+ vssd1 vccd1 vccd1 net2695 sky130_fd_sc_hd__dlygate4sd3_1
X_08834_ net583 _02953_ vssd1 vssd1 vccd1 vccd1 _04776_ sky130_fd_sc_hd__and2_1
Xhold1213 team_03_WB.instance_to_wrap.core.register_file.registers_state\[717\] vssd1
+ vssd1 vccd1 vccd1 net2706 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10541__B1 net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1224 team_03_WB.instance_to_wrap.core.register_file.registers_state\[72\] vssd1
+ vssd1 vccd1 vccd1 net2717 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1002_A net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1235 team_03_WB.instance_to_wrap.core.register_file.registers_state\[604\] vssd1
+ vssd1 vccd1 vccd1 net2728 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11884__A3 net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07643__A net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1246 team_03_WB.instance_to_wrap.core.register_file.registers_state\[582\] vssd1
+ vssd1 vccd1 vccd1 net2739 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1257 team_03_WB.instance_to_wrap.core.register_file.registers_state\[730\] vssd1
+ vssd1 vccd1 vccd1 net2750 sky130_fd_sc_hd__dlygate4sd3_1
X_08765_ net1052 team_03_WB.instance_to_wrap.core.register_file.registers_state\[835\]
+ net1004 team_03_WB.instance_to_wrap.core.register_file.registers_state\[867\] net1065
+ vssd1 vssd1 vccd1 vccd1 _04707_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout462_A net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1268 team_03_WB.instance_to_wrap.core.register_file.registers_state\[838\] vssd1
+ vssd1 vccd1 vccd1 net2761 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1279 team_03_WB.instance_to_wrap.CPU_DAT_O\[4\] vssd1 vssd1 vccd1 vccd1 net2772
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11165__A net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07716_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[269\] net800
+ _02871_ _03657_ vssd1 vssd1 vccd1 vccd1 _03658_ sky130_fd_sc_hd__o211a_1
X_08696_ net857 _04636_ _04637_ vssd1 vssd1 vccd1 vccd1 _04638_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_68_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_68_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07647_ net730 _03587_ _03588_ net1164 vssd1 vssd1 vccd1 vccd1 _03589_ sky130_fd_sc_hd__o211ai_1
XANTENNA_fanout727_A net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout348_X net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08474__A _04080_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07578_ net1092 team_03_WB.instance_to_wrap.core.register_file.registers_state\[952\]
+ net895 vssd1 vssd1 vccd1 vccd1 _03520_ sky130_fd_sc_hd__or3_1
XFILLER_0_137_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_153_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09317_ net592 _05258_ vssd1 vssd1 vccd1 vccd1 _05259_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_24_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_118_2800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_157_3594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout515_X net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_940 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09857__X _05799_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09248_ _04294_ _05189_ vssd1 vssd1 vccd1 vccd1 _05190_ sky130_fd_sc_hd__nor2_1
XANTENNA__07473__B1 net1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_114_2708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_2719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08017__A2 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09179_ net552 _04807_ net540 net582 vssd1 vssd1 vccd1 vccd1 _05121_ sky130_fd_sc_hd__o22a_1
XANTENNA__08648__S0 net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_274 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07225__B1 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11210_ net274 net2367 net486 vssd1 vssd1 vccd1 vccd1 _02198_ sky130_fd_sc_hd__mux2_1
X_12190_ net1499 vssd1 vssd1 vccd1 vccd1 _02363_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__07818__A net1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11021__B2 net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08422__C1 net1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09736__C net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout884_X net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08973__B1 net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11141_ net649 _06646_ vssd1 vssd1 vccd1 vccd1 _06647_ sky130_fd_sc_hd__and2_1
XFILLER_0_102_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_352 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07029__S net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11072_ net834 _06422_ vssd1 vssd1 vccd1 vccd1 _06614_ sky130_fd_sc_hd__and2_2
XANTENNA__11059__B net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput100 wbs_dat_i[0] vssd1 vssd1 vccd1 vccd1 net100 sky130_fd_sc_hd__clkbuf_1
XANTENNA__07256__C net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14900_ clknet_leaf_58_wb_clk_i _02663_ _01265_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.pc.current_pc\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08725__B1 net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10023_ net91 net90 net88 net87 vssd1 vssd1 vccd1 vccd1 _05901_ sky130_fd_sc_hd__or4bb_1
XANTENNA__13555__A net1435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10532__B1 net1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input23_A DAT_I[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14831_ clknet_leaf_94_wb_clk_i net1717 _01196_ vssd1 vssd1 vccd1 vccd1 net152 sky130_fd_sc_hd__dfrtp_1
XANTENNA__08001__X _03943_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14762_ clknet_leaf_61_wb_clk_i _02526_ _01127_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_11974_ _06447_ _06751_ _06394_ vssd1 vssd1 vccd1 vccd1 _06816_ sky130_fd_sc_hd__or3b_1
X_13713_ clknet_leaf_139_wb_clk_i _01477_ _00078_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[67\]
+ sky130_fd_sc_hd__dfrtp_1
X_10925_ net690 _06511_ _06512_ _06510_ vssd1 vssd1 vccd1 vccd1 _06513_ sky130_fd_sc_hd__o31a_2
X_14693_ clknet_leaf_59_wb_clk_i _02457_ _01058_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.ADR_I\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07700__A1 net1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13644_ net1405 vssd1 vssd1 vccd1 vccd1 _01408_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_141_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_141_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__12037__B1 net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10856_ _06380_ _06389_ vssd1 vssd1 vccd1 vccd1 _06455_ sky130_fd_sc_hd__nor2_2
XFILLER_0_73_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11522__B net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13575_ net1432 vssd1 vssd1 vccd1 vccd1 _01339_ sky130_fd_sc_hd__inv_2
X_10787_ net313 net309 net316 vssd1 vssd1 vccd1 vccd1 _06397_ sky130_fd_sc_hd__or3_1
XFILLER_0_87_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10063__A2 net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11260__A1 net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12526_ net1274 vssd1 vssd1 vccd1 vccd1 _00290_ sky130_fd_sc_hd__inv_2
XANTENNA__11241__C net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08661__C1 net1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09927__B net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12457_ net1254 vssd1 vssd1 vccd1 vccd1 _00221_ sky130_fd_sc_hd__inv_2
XFILLER_0_48_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11012__A1 net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11408_ net300 net2624 net397 vssd1 vssd1 vccd1 vccd1 _02072_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_10_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12388_ net1356 vssd1 vssd1 vccd1 vccd1 _00152_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_91_2240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14127_ clknet_leaf_135_wb_clk_i _01891_ _00492_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[481\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_91_2251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11339_ net1247 net836 net279 net668 vssd1 vssd1 vccd1 vccd1 _06722_ sky130_fd_sc_hd__and4_1
XANTENNA__09943__A _04029_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14058_ clknet_leaf_2_wb_clk_i _01822_ _00423_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[412\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_123_1085 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07519__A1 net1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08716__B1 net999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13465__A net1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13009_ net1268 vssd1 vssd1 vccd1 vccd1 _00773_ sky130_fd_sc_hd__inv_2
XANTENNA__09662__B _04207_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06880_ _02808_ _02817_ _02820_ team_03_WB.instance_to_wrap.core.decoder.inst\[31\]
+ vssd1 vssd1 vccd1 vccd1 _02822_ sky130_fd_sc_hd__and4bb_1
XANTENNA__10523__B1 net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07463__A net1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08550_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[190\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[158\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[62\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[30\]
+ net955 net917 vssd1 vssd1 vccd1 vccd1 _04492_ sky130_fd_sc_hd__mux4_1
X_07501_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[7\] net803
+ net735 _03442_ vssd1 vssd1 vccd1 vccd1 _03443_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_46_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08481_ _04421_ _04422_ net864 vssd1 vssd1 vccd1 vccd1 _04423_ sky130_fd_sc_hd__o21a_1
XFILLER_0_43_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_46_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07432_ net1177 team_03_WB.instance_to_wrap.core.register_file.registers_state\[52\]
+ net880 vssd1 vssd1 vccd1 vccd1 _03374_ sky130_fd_sc_hd__and3_1
XANTENNA__12028__B1 net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_536 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08294__A _04235_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_238 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_63_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07363_ net1146 _03297_ _03298_ net1160 vssd1 vssd1 vccd1 vccd1 _03305_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_63_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_3144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09102_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[14\] net1001
+ net924 _05043_ vssd1 vssd1 vccd1 vccd1 _05044_ sky130_fd_sc_hd__o211a_1
XANTENNA__10054__A2 net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07455__B1 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08798__A3 net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_3155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07294_ net1202 team_03_WB.instance_to_wrap.core.register_file.registers_state\[457\]
+ vssd1 vssd1 vccd1 vccd1 _03236_ sky130_fd_sc_hd__or2_1
XFILLER_0_73_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_150_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11859__S net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09033_ net1059 team_03_WB.instance_to_wrap.core.register_file.registers_state\[656\]
+ net1013 team_03_WB.instance_to_wrap.core.register_file.registers_state\[688\] net928
+ vssd1 vssd1 vccd1 vccd1 _04975_ sky130_fd_sc_hd__a221o_1
XFILLER_0_4_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_152_3491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout308_A _06396_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold310 team_03_WB.instance_to_wrap.ADR_I\[15\] vssd1 vssd1 vccd1 vccd1 net1803 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08404__C1 net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold321 team_03_WB.instance_to_wrap.core.register_file.registers_state\[960\] vssd1
+ vssd1 vccd1 vccd1 net1814 sky130_fd_sc_hd__dlygate4sd3_1
Xhold332 team_03_WB.instance_to_wrap.core.register_file.registers_state\[307\] vssd1
+ vssd1 vccd1 vccd1 net1825 sky130_fd_sc_hd__dlygate4sd3_1
Xhold343 team_03_WB.instance_to_wrap.core.register_file.registers_state\[315\] vssd1
+ vssd1 vccd1 vccd1 net1836 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold354 team_03_WB.instance_to_wrap.core.register_file.registers_state\[880\] vssd1
+ vssd1 vccd1 vccd1 net1847 sky130_fd_sc_hd__dlygate4sd3_1
Xhold365 team_03_WB.instance_to_wrap.core.register_file.registers_state\[35\] vssd1
+ vssd1 vccd1 vccd1 net1858 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06966__C1 net1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold376 team_03_WB.instance_to_wrap.core.register_file.registers_state\[425\] vssd1
+ vssd1 vccd1 vccd1 net1869 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1217_A net1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold387 team_03_WB.instance_to_wrap.core.register_file.registers_state\[413\] vssd1
+ vssd1 vccd1 vccd1 net1880 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1014 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout801 net805 vssd1 vssd1 vccd1 vccd1 net801 sky130_fd_sc_hd__clkbuf_4
Xhold398 team_03_WB.instance_to_wrap.core.register_file.registers_state\[412\] vssd1
+ vssd1 vccd1 vccd1 net1891 sky130_fd_sc_hd__dlygate4sd3_1
X_09935_ _04069_ net663 vssd1 vssd1 vccd1 vccd1 _05872_ sky130_fd_sc_hd__nor2_2
Xfanout812 net816 vssd1 vssd1 vccd1 vccd1 net812 sky130_fd_sc_hd__buf_4
XFILLER_0_110_182 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout823 net824 vssd1 vssd1 vccd1 vccd1 net823 sky130_fd_sc_hd__buf_4
Xfanout834 _06387_ vssd1 vssd1 vccd1 vccd1 net834 sky130_fd_sc_hd__clkbuf_8
XANTENNA__10999__A net1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11594__S net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout845 _06303_ vssd1 vssd1 vccd1 vccd1 net845 sky130_fd_sc_hd__buf_4
XANTENNA__06981__A2 _02921_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout298_X net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1069 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout856 net858 vssd1 vssd1 vccd1 vccd1 net856 sky130_fd_sc_hd__buf_4
X_09866_ _04824_ _05126_ _05371_ _05806_ _05807_ vssd1 vssd1 vccd1 vccd1 _05808_ sky130_fd_sc_hd__a311o_1
Xfanout867 net870 vssd1 vssd1 vccd1 vccd1 net867 sky130_fd_sc_hd__buf_8
XANTENNA__10514__B1 net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout878 net879 vssd1 vssd1 vccd1 vccd1 net878 sky130_fd_sc_hd__buf_2
Xhold1010 team_03_WB.instance_to_wrap.core.register_file.registers_state\[330\] vssd1
+ vssd1 vccd1 vccd1 net2503 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1021 team_03_WB.instance_to_wrap.core.register_file.registers_state\[623\] vssd1
+ vssd1 vccd1 vccd1 net2514 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout889 net891 vssd1 vssd1 vccd1 vccd1 net889 sky130_fd_sc_hd__clkbuf_4
Xhold1032 team_03_WB.instance_to_wrap.core.register_file.registers_state\[539\] vssd1
+ vssd1 vccd1 vccd1 net2525 sky130_fd_sc_hd__dlygate4sd3_1
X_08817_ net1055 team_03_WB.instance_to_wrap.core.register_file.registers_state\[833\]
+ net1005 team_03_WB.instance_to_wrap.core.register_file.registers_state\[865\] net1065
+ vssd1 vssd1 vccd1 vccd1 _04759_ sky130_fd_sc_hd__a221o_1
Xhold1043 team_03_WB.instance_to_wrap.core.register_file.registers_state\[158\] vssd1
+ vssd1 vccd1 vccd1 net2536 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout844_A net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09797_ _05110_ _05119_ _05130_ _05113_ net562 net570 vssd1 vssd1 vccd1 vccd1 _05739_
+ sky130_fd_sc_hd__mux4_1
Xhold1054 team_03_WB.instance_to_wrap.core.register_file.registers_state\[851\] vssd1
+ vssd1 vccd1 vccd1 net2547 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1065 team_03_WB.instance_to_wrap.core.register_file.registers_state\[210\] vssd1
+ vssd1 vccd1 vccd1 net2558 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07930__A1 net1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1076 team_03_WB.instance_to_wrap.core.register_file.registers_state\[864\] vssd1
+ vssd1 vccd1 vccd1 net2569 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10003__S net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_2567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08748_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[419\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[387\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[291\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[259\]
+ net980 net1076 vssd1 vssd1 vccd1 vccd1 _04690_ sky130_fd_sc_hd__mux4_1
Xhold1087 team_03_WB.instance_to_wrap.core.register_file.registers_state\[911\] vssd1
+ vssd1 vccd1 vccd1 net2580 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_107_2578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1098 team_03_WB.instance_to_wrap.core.register_file.registers_state\[608\] vssd1
+ vssd1 vccd1 vccd1 net2591 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_159_3634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_3_2_0_wb_clk_i_X clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_159_3645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08679_ net435 net430 _04620_ net550 vssd1 vssd1 vccd1 vccd1 _04621_ sky130_fd_sc_hd__o31a_1
XANTENNA_fanout632_X net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10938__S net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07143__C1 net1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10710_ net523 _06344_ _06345_ net528 net1617 vssd1 vssd1 vccd1 vccd1 _02459_ sky130_fd_sc_hd__a32o_1
XANTENNA__12019__B1 net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08408__S net992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11690_ _06732_ net379 net338 net1871 vssd1 vssd1 vccd1 vccd1 _01844_ sky130_fd_sc_hd__a22o_1
X_10641_ net1185 net1964 net844 vssd1 vssd1 vccd1 vccd1 _02487_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_761 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_912 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11242__A1 net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13360_ net1325 vssd1 vssd1 vccd1 vccd1 _01124_ sky130_fd_sc_hd__inv_2
XANTENNA__07446__B1 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11061__C net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10572_ net1684 net534 net601 _05882_ vssd1 vssd1 vccd1 vccd1 _02551_ sky130_fd_sc_hd__a22o_1
XANTENNA__08643__C1 net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_165_Right_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07997__A1 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12311_ net1390 vssd1 vssd1 vccd1 vccd1 _00075_ sky130_fd_sc_hd__inv_2
X_13291_ net1322 vssd1 vssd1 vccd1 vccd1 _01055_ sky130_fd_sc_hd__inv_2
XFILLER_0_161_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15030_ clknet_leaf_101_wb_clk_i _02750_ _01395_ vssd1 vssd1 vccd1 vccd1 net186 sky130_fd_sc_hd__dfrtp_1
X_12242_ net2652 vssd1 vssd1 vccd1 vccd1 _01415_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__07548__A _03489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_959 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07749__A1 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11545__A2 net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12173_ net1602 vssd1 vssd1 vccd1 vccd1 _02380_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11124_ net280 net649 net704 net696 vssd1 vssd1 vccd1 vccd1 _06637_ sky130_fd_sc_hd__and4_1
X_11055_ net655 net705 _06541_ net829 vssd1 vssd1 vccd1 vccd1 _06605_ sky130_fd_sc_hd__and4_1
XANTENNA__10505__B1 net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09913__D _05686_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08174__A1 net1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07283__A net1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10006_ _03458_ net1962 net288 vssd1 vssd1 vccd1 vccd1 _02708_ sky130_fd_sc_hd__mux2_1
XANTENNA__07921__A1 net1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14814_ clknet_leaf_96_wb_clk_i net1662 _01179_ vssd1 vssd1 vccd1 vccd1 net165 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_98_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14745_ clknet_leaf_48_wb_clk_i _02509_ _01110_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_28_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11957_ net641 _06734_ net474 net366 net2443 vssd1 vssd1 vccd1 vccd1 _01586_ sky130_fd_sc_hd__a32o_1
XFILLER_0_80_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10908_ net686 _06497_ _06498_ _06496_ vssd1 vssd1 vccd1 vccd1 _06499_ sky130_fd_sc_hd__o31a_4
X_14676_ clknet_leaf_85_wb_clk_i _02440_ _01041_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.ADR_I\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09774__A1_N net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11888_ net623 _06697_ net454 net371 net2115 vssd1 vssd1 vccd1 vccd1 _01653_ sky130_fd_sc_hd__a32o_1
XFILLER_0_67_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13627_ net1415 vssd1 vssd1 vccd1 vccd1 _01391_ sky130_fd_sc_hd__inv_2
X_10839_ team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[22\] _05865_ net318 _06403_
+ net686 vssd1 vssd1 vccd1 vccd1 _06440_ sky130_fd_sc_hd__a41o_1
XANTENNA__10149__A _03138_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12025__A3 net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10036__A2 net1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07437__B1 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13558_ net1420 vssd1 vssd1 vccd1 vccd1 _01322_ sky130_fd_sc_hd__inv_2
XFILLER_0_27_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_132_Right_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07988__A1 net1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12509_ net1383 vssd1 vssd1 vccd1 vccd1 _00273_ sky130_fd_sc_hd__inv_2
XFILLER_0_81_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_140_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13489_ net1341 vssd1 vssd1 vccd1 vccd1 _01253_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_734 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_751 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_3041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_130_3052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_39_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_42 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07981_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[272\] net804
+ _02871_ _03922_ vssd1 vssd1 vccd1 vccd1 _03923_ sky130_fd_sc_hd__o211a_1
X_09720_ _05217_ _05227_ _05660_ vssd1 vssd1 vccd1 vccd1 _05662_ sky130_fd_sc_hd__and3_1
X_06932_ _02865_ _02866_ _02868_ net1136 net1166 vssd1 vssd1 vccd1 vccd1 _02874_ sky130_fd_sc_hd__o221a_1
XFILLER_0_129_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08165__B2 net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09651_ _05592_ vssd1 vssd1 vccd1 vccd1 _05593_ sky130_fd_sc_hd__inv_2
XANTENNA__09901__A2 _05841_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11427__B net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06863_ team_03_WB.instance_to_wrap.core.control_logic.instruction\[2\] team_03_WB.instance_to_wrap.core.control_logic.instruction\[1\]
+ team_03_WB.instance_to_wrap.core.control_logic.instruction\[0\] vssd1 vssd1 vccd1
+ vccd1 _02805_ sky130_fd_sc_hd__nand3b_1
XANTENNA__07912__A1 net1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08602_ net930 _04542_ _04543_ net865 vssd1 vssd1 vccd1 vccd1 _04544_ sky130_fd_sc_hd__a211o_1
X_09582_ net547 _04417_ _05103_ net553 vssd1 vssd1 vccd1 vccd1 _05524_ sky130_fd_sc_hd__a211o_1
XANTENNA__11146__C net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1086 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_26_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08533_ _04461_ _04474_ net849 vssd1 vssd1 vccd1 vccd1 _04475_ sky130_fd_sc_hd__mux2_8
XTAP_TAPCELL_ROW_65_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09665__A1 _02804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_166_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11443__A net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_171 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_3_7_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_7_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_08464_ net1227 team_03_WB.instance_to_wrap.core.register_file.registers_state\[220\]
+ net953 team_03_WB.instance_to_wrap.core.register_file.registers_state\[252\] net933
+ vssd1 vssd1 vccd1 vccd1 _04406_ sky130_fd_sc_hd__o221a_1
XFILLER_0_49_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11472__B2 net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_2464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_102_2475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11162__B net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07415_ net1084 net889 team_03_WB.instance_to_wrap.core.register_file.registers_state\[532\]
+ vssd1 vssd1 vccd1 vccd1 _03357_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_154_3531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08395_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[441\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[409\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[313\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[281\]
+ net991 net1079 vssd1 vssd1 vccd1 vccd1 _04337_ sky130_fd_sc_hd__mux4_1
XFILLER_0_107_208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout425_A net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_154_3542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1167_A net1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_169_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07346_ net1171 team_03_WB.instance_to_wrap.core.register_file.registers_state\[220\]
+ vssd1 vssd1 vccd1 vccd1 _03288_ sky130_fd_sc_hd__or2_1
XFILLER_0_18_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11589__S net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11775__A2 net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07277_ net1201 team_03_WB.instance_to_wrap.core.register_file.registers_state\[713\]
+ net782 team_03_WB.instance_to_wrap.core.register_file.registers_state\[745\] net751
+ vssd1 vssd1 vccd1 vccd1 _03219_ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout1334_A net1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09016_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[48\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[16\]
+ net984 vssd1 vssd1 vccd1 vccd1 _04958_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11527__A2 net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout794_A net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold140 team_03_WB.instance_to_wrap.ADR_I\[27\] vssd1 vssd1 vccd1 vccd1 net1633 sky130_fd_sc_hd__dlygate4sd3_1
Xhold151 team_03_WB.instance_to_wrap.CPU_DAT_I\[5\] vssd1 vssd1 vccd1 vccd1 net1644
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold162 _02613_ vssd1 vssd1 vccd1 vccd1 net1655 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10735__B1 net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1122_X net1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold173 team_03_WB.instance_to_wrap.CPU_DAT_I\[2\] vssd1 vssd1 vccd1 vccd1 net1666
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold184 team_03_WB.instance_to_wrap.ADR_I\[26\] vssd1 vssd1 vccd1 vccd1 net1677 sky130_fd_sc_hd__dlygate4sd3_1
Xhold195 net113 vssd1 vssd1 vccd1 vccd1 net1688 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout582_X net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout961_A net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout620 net621 vssd1 vssd1 vccd1 vccd1 net620 sky130_fd_sc_hd__clkbuf_4
Xfanout631 _06458_ vssd1 vssd1 vccd1 vccd1 net631 sky130_fd_sc_hd__clkbuf_4
X_09918_ _02829_ _02837_ vssd1 vssd1 vccd1 vccd1 _05860_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_109_2607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout642 net645 vssd1 vssd1 vccd1 vccd1 net642 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10081__X _05925_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout653 net655 vssd1 vssd1 vccd1 vccd1 net653 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_109_2618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout664 net666 vssd1 vssd1 vccd1 vccd1 net664 sky130_fd_sc_hd__buf_2
XANTENNA__08156__A1 net1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout675 _05948_ vssd1 vssd1 vccd1 vccd1 net675 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07307__S net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout686 net687 vssd1 vssd1 vccd1 vccd1 net686 sky130_fd_sc_hd__clkbuf_4
X_09849_ _04834_ _05520_ _05786_ _05790_ vssd1 vssd1 vccd1 vccd1 _05791_ sky130_fd_sc_hd__o211a_1
Xfanout697 net698 vssd1 vssd1 vccd1 vccd1 net697 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11337__B net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout847_X net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07903__A1 net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12860_ net1419 vssd1 vssd1 vccd1 vccd1 _00624_ sky130_fd_sc_hd__inv_2
XANTENNA__09522__S net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09105__B1 net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11811_ _06637_ net460 net323 net1929 vssd1 vssd1 vccd1 vccd1 _01728_ sky130_fd_sc_hd__a22o_1
XFILLER_0_68_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12791_ net1386 vssd1 vssd1 vccd1 vccd1 _00555_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_1_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11353__A _06446_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14530_ clknet_leaf_177_wb_clk_i _02294_ _00895_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[884\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_166_620 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11463__A1 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11742_ net1924 net266 net336 vssd1 vssd1 vccd1 vccd1 _01794_ sky130_fd_sc_hd__mux2_1
XANTENNA__08864__C1 net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1040 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11072__B _06422_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14461_ clknet_leaf_165_wb_clk_i _02225_ _00826_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[815\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11673_ net2177 net263 net344 vssd1 vssd1 vccd1 vccd1 _01860_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_139 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13412_ net1427 vssd1 vssd1 vccd1 vccd1 _01176_ sky130_fd_sc_hd__inv_2
XFILLER_0_113_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10624_ net2121 team_03_WB.instance_to_wrap.CPU_DAT_O\[5\] net842 vssd1 vssd1 vccd1
+ vccd1 _02504_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_12_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input90_A wbs_adr_i[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14392_ clknet_leaf_186_wb_clk_i _02156_ _00757_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[746\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_133_Left_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_515 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11499__S net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11766__A2 net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13343_ net1335 vssd1 vssd1 vccd1 vccd1 _01107_ sky130_fd_sc_hd__inv_2
XFILLER_0_36_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10555_ _02765_ _06296_ _06297_ vssd1 vssd1 vccd1 vccd1 _06298_ sky130_fd_sc_hd__or3_4
XANTENNA__08092__B1 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13274_ net1423 vssd1 vssd1 vccd1 vccd1 _01038_ sky130_fd_sc_hd__inv_2
XFILLER_0_11_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10486_ net115 net1027 net905 net1564 vssd1 vssd1 vccd1 vccd1 _02623_ sky130_fd_sc_hd__a22o_1
X_15013_ clknet_leaf_102_wb_clk_i _02733_ _01378_ vssd1 vssd1 vccd1 vccd1 net174 sky130_fd_sc_hd__dfrtp_1
X_12225_ net1555 vssd1 vssd1 vccd1 vccd1 _01432_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__09041__C1 net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09493__A net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12156_ net1536 vssd1 vssd1 vccd1 vccd1 _02397_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__06910__A net1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11107_ net834 _06523_ vssd1 vssd1 vccd1 vccd1 _06629_ sky130_fd_sc_hd__and2_1
X_12087_ net618 _06653_ net451 net439 net1879 vssd1 vssd1 vccd1 vccd1 _01460_ sky130_fd_sc_hd__a32o_1
XPHY_EDGE_ROW_142_Left_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09344__B1 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11038_ net1044 net836 net270 net670 vssd1 vssd1 vccd1 vccd1 _06595_ sky130_fd_sc_hd__and4_1
XANTENNA__11247__B net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11151__B1 net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07355__C1 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09432__S net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09647__A1 net1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12989_ net1389 vssd1 vssd1 vccd1 vccd1 _00753_ sky130_fd_sc_hd__inv_2
XANTENNA__11263__A net1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_2058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11454__A1 net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_2069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14728_ clknet_leaf_49_wb_clk_i _02492_ _01093_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.decoder.inst\[25\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__07122__A2 _03059_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_156_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_815 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14659_ clknet_leaf_47_wb_clk_i _02423_ _01024_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1013\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_60_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_60_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_151_Left_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07200_ _03140_ _03141_ net740 vssd1 vssd1 vccd1 vccd1 _03142_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08180_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[51\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[19\]
+ net959 vssd1 vssd1 vccd1 vccd1 _04122_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07131_ net752 _03072_ net1166 vssd1 vssd1 vccd1 vccd1 _03073_ sky130_fd_sc_hd__o21a_1
XFILLER_0_125_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11202__S net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_520 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07062_ net733 _03003_ _03002_ vssd1 vssd1 vccd1 vccd1 _03004_ sky130_fd_sc_hd__o21a_1
Xoutput201 net201 vssd1 vssd1 vccd1 vccd1 gpio_oeb[5] sky130_fd_sc_hd__buf_2
XFILLER_0_3_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput212 net212 vssd1 vssd1 vccd1 vccd1 gpio_out[15] sky130_fd_sc_hd__buf_2
Xoutput223 net223 vssd1 vssd1 vccd1 vccd1 gpio_out[26] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_11_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_58_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput234 net234 vssd1 vssd1 vccd1 vccd1 gpio_out[6] sky130_fd_sc_hd__buf_2
Xoutput245 net245 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[16] sky130_fd_sc_hd__buf_2
XANTENNA__10717__B1 net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12822__A net1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput256 net256 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[30] sky130_fd_sc_hd__buf_2
XANTENNA__11390__B1 net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07594__C1 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_160_Left_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11438__A net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07964_ net1193 team_03_WB.instance_to_wrap.core.register_file.registers_state\[48\]
+ net886 vssd1 vssd1 vccd1 vccd1 _03906_ sky130_fd_sc_hd__and3_1
XFILLER_0_4_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_147_3390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09703_ net351 _05385_ _05644_ vssd1 vssd1 vccd1 vccd1 _05645_ sky130_fd_sc_hd__a21o_1
XANTENNA__09690__X _05632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11157__B net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06915_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[4\] net804
+ net734 _02856_ vssd1 vssd1 vccd1 vccd1 _02857_ sky130_fd_sc_hd__o211a_1
XANTENNA__09886__A1 _04816_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07895_ net1187 team_03_WB.instance_to_wrap.core.register_file.registers_state\[495\]
+ net877 _03836_ net1130 vssd1 vssd1 vccd1 vccd1 _03837_ sky130_fd_sc_hd__a311o_1
XANTENNA__11872__S net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout375_A _06812_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09634_ net567 _05493_ vssd1 vssd1 vccd1 vccd1 _05576_ sky130_fd_sc_hd__nand2_1
XANTENNA__07922__Y _03864_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10496__A2 net1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06846_ net1214 vssd1 vssd1 vccd1 vccd1 _02789_ sky130_fd_sc_hd__inv_2
XANTENNA__07897__B1 _02870_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_2504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10996__B net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_2515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07005__A_N _02945_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09565_ net573 _05506_ vssd1 vssd1 vccd1 vccd1 _05507_ sky130_fd_sc_hd__and2_1
XANTENNA__09638__A1 net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout542_A net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11173__A net1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_2851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08516_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[895\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[863\]
+ net952 vssd1 vssd1 vccd1 vccd1 _04458_ sky130_fd_sc_hd__mux2_1
XANTENNA__11445__A1 net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_2862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09496_ _05436_ _05437_ net574 vssd1 vssd1 vccd1 vccd1 _05438_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08846__C1 net1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08447_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[572\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[540\]
+ net953 vssd1 vssd1 vccd1 vccd1 _04389_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout330_X net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_234 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1072_X net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout807_A net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08482__A net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08378_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[886\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[854\]
+ net970 vssd1 vssd1 vccd1 vccd1 _04320_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11748__A2 net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07329_ net1087 team_03_WB.instance_to_wrap.core.register_file.registers_state\[509\]
+ net893 vssd1 vssd1 vccd1 vccd1 _03271_ sky130_fd_sc_hd__or3_1
XFILLER_0_33_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11112__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07098__A net1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10340_ _06175_ _06176_ net283 vssd1 vssd1 vccd1 vccd1 _06177_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07821__B1 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout797_X net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10271_ _04383_ team_03_WB.instance_to_wrap.core.pc.current_pc\[26\] net673 vssd1
+ vssd1 vccd1 vccd1 _06113_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_1130 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09023__C1 net1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12010_ _06760_ net458 net360 net2213 vssd1 vssd1 vccd1 vccd1 _01535_ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_47_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout964_X net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1404 net1408 vssd1 vssd1 vccd1 vccd1 net1404 sky130_fd_sc_hd__buf_4
XANTENNA__14720__Q team_03_WB.instance_to_wrap.core.decoder.inst\[17\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_167_3799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1415 net1417 vssd1 vssd1 vccd1 vccd1 net1415 sky130_fd_sc_hd__buf_4
Xfanout1426 net1436 vssd1 vssd1 vccd1 vccd1 net1426 sky130_fd_sc_hd__buf_2
Xfanout1437 net1438 vssd1 vssd1 vccd1 vccd1 net1437 sky130_fd_sc_hd__clkbuf_4
Xfanout450 _06801_ vssd1 vssd1 vccd1 vccd1 net450 sky130_fd_sc_hd__buf_4
Xfanout461 net462 vssd1 vssd1 vccd1 vccd1 net461 sky130_fd_sc_hd__buf_4
Xfanout472 net481 vssd1 vssd1 vccd1 vccd1 net472 sky130_fd_sc_hd__buf_2
X_13961_ clknet_leaf_76_wb_clk_i _01725_ _00326_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[315\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout483 _06779_ vssd1 vssd1 vccd1 vccd1 net483 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_6_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout494 net496 vssd1 vssd1 vccd1 vccd1 net494 sky130_fd_sc_hd__clkbuf_2
XANTENNA__11782__S net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12912_ net1412 vssd1 vssd1 vccd1 vccd1 _00676_ sky130_fd_sc_hd__inv_2
X_13892_ clknet_leaf_29_wb_clk_i _01656_ _00257_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[246\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_159_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12843_ net1282 vssd1 vssd1 vccd1 vccd1 _00607_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_17_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08837__C1 _04778_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12774_ net1300 vssd1 vssd1 vccd1 vccd1 _00538_ sky130_fd_sc_hd__inv_2
XFILLER_0_84_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08301__A1 net1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14513_ clknet_leaf_140_wb_clk_i _02277_ _00878_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[867\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_48_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_48_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_11725_ net596 _06479_ net456 _06808_ net1949 vssd1 vssd1 vccd1 vccd1 _01811_ sky130_fd_sc_hd__a32o_1
XFILLER_0_83_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_859 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14444_ clknet_leaf_14_wb_clk_i _02208_ _00809_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[798\]
+ sky130_fd_sc_hd__dfrtp_1
X_11656_ net2600 _06469_ net343 vssd1 vssd1 vccd1 vccd1 _01877_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_656 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06905__A net1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10607_ net2648 net1806 net840 vssd1 vssd1 vccd1 vccd1 _02521_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_86_wb_clk_i_A clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_14375_ clknet_leaf_108_wb_clk_i _02139_ _00740_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[729\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_36_183 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11587_ net274 net2472 net447 vssd1 vssd1 vccd1 vccd1 _01942_ sky130_fd_sc_hd__mux2_1
X_13326_ net1317 vssd1 vssd1 vccd1 vccd1 _01090_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_239 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10538_ net147 net1034 net1026 net1614 vssd1 vssd1 vccd1 vccd1 _02572_ sky130_fd_sc_hd__a22o_1
Xhold909 team_03_WB.instance_to_wrap.core.register_file.registers_state\[908\] vssd1
+ vssd1 vccd1 vccd1 net2402 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_49_1074 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_687 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13257_ net1255 vssd1 vssd1 vccd1 vccd1 _01021_ sky130_fd_sc_hd__inv_2
XANTENNA__09935__B net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10469_ _02765_ team_03_WB.instance_to_wrap.BUSY_O vssd1 vssd1 vccd1 vccd1 _06281_
+ sky130_fd_sc_hd__nor2_1
XANTENNA__12642__A net1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08368__A1 net1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12208_ net1533 vssd1 vssd1 vccd1 vccd1 _02345_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__08331__S net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13188_ net1367 vssd1 vssd1 vccd1 vccd1 _00952_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11372__B1 net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07576__C1 net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12139_ net1584 vssd1 vssd1 vccd1 vccd1 _02414_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_53_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09951__A _03169_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07591__A2 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09868__A1 net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07328__C1 net1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_84_2109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07680_ net1174 team_03_WB.instance_to_wrap.core.register_file.registers_state\[734\]
+ net761 team_03_WB.instance_to_wrap.core.register_file.registers_state\[766\] net743
+ vssd1 vssd1 vccd1 vccd1 _03622_ sky130_fd_sc_hd__o221a_1
XFILLER_0_126_98 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09350_ _03989_ _05149_ vssd1 vssd1 vccd1 vccd1 _05292_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_75_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08301_ net1236 team_03_WB.instance_to_wrap.core.register_file.registers_state\[216\]
+ net972 team_03_WB.instance_to_wrap.core.register_file.registers_state\[248\] net939
+ vssd1 vssd1 vccd1 vccd1 _04243_ sky130_fd_sc_hd__o221a_1
X_09281_ net609 _05145_ vssd1 vssd1 vccd1 vccd1 _05223_ sky130_fd_sc_hd__nor2_1
XFILLER_0_117_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08232_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[689\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[657\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[561\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[529\]
+ net960 net919 vssd1 vssd1 vccd1 vccd1 _04174_ sky130_fd_sc_hd__mux4_1
XFILLER_0_172_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_662 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07410__S net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10982__D net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08163_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[564\] net959
+ net918 vssd1 vssd1 vccd1 vccd1 _04105_ sky130_fd_sc_hd__o21a_1
XFILLER_0_160_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_1028 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07114_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[161\] net778
+ net748 _03055_ vssd1 vssd1 vccd1 vccd1 _03056_ sky130_fd_sc_hd__o211a_1
XANTENNA__07803__B1 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_740 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08094_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[154\] net760
+ net725 _04035_ vssd1 vssd1 vccd1 vccd1 _04036_ sky130_fd_sc_hd__a211o_1
XFILLER_0_30_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11867__S net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload60 clknet_leaf_39_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload60/Y sky130_fd_sc_hd__clkinv_4
Xclkload71 clknet_leaf_51_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload71/Y sky130_fd_sc_hd__clkinv_2
X_07045_ net1134 _02984_ _02983_ net1165 vssd1 vssd1 vccd1 vccd1 _02987_ sky130_fd_sc_hd__o211a_1
XFILLER_0_42_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_1960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09845__B net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload82 clknet_leaf_29_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload82/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_141_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_149_3430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload93 clknet_leaf_62_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload93/Y sky130_fd_sc_hd__inv_6
XFILLER_0_113_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08359__A1 net1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_149_3441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout492_A net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07031__A1 team_03_WB.instance_to_wrap.core.decoder.inst\[23\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11168__A net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15089__1475 vssd1 vssd1 vccd1 vccd1 _15089__1475/HI net1475 sky130_fd_sc_hd__conb_1
X_08996_ net1045 team_03_WB.instance_to_wrap.core.register_file.registers_state\[970\]
+ net995 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1002\] net1062
+ vssd1 vssd1 vccd1 vccd1 _04938_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_145_3349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11115__A0 net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07084__C net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07947_ net1182 team_03_WB.instance_to_wrap.core.register_file.registers_state\[855\]
+ vssd1 vssd1 vccd1 vccd1 _03889_ sky130_fd_sc_hd__or2_1
XFILLER_0_138_1113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout280_X net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout378_X net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout757_A net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_162_3696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11666__A1 _06628_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07878_ net823 _03815_ _03819_ net719 vssd1 vssd1 vccd1 vccd1 _03820_ sky130_fd_sc_hd__o31a_1
XFILLER_0_98_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08531__A1 net1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09617_ net553 _05365_ net568 vssd1 vssd1 vccd1 vccd1 _05559_ sky130_fd_sc_hd__o21a_1
X_06829_ team_03_WB.instance_to_wrap.core.pc.current_pc\[20\] vssd1 vssd1 vccd1 vccd1
+ _02772_ sky130_fd_sc_hd__inv_2
XFILLER_0_74_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout924_A net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09548_ _03529_ _04267_ net538 vssd1 vssd1 vccd1 vccd1 _05490_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_78_562 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_120_wb_clk_i_A clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12091__A1 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09479_ net564 _05420_ vssd1 vssd1 vccd1 vccd1 _05421_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout712_X net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_459 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11053__D net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11510_ _06627_ net2609 net388 vssd1 vssd1 vccd1 vccd1 _01996_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12490_ net1284 vssd1 vssd1 vccd1 vccd1 _00254_ sky130_fd_sc_hd__inv_2
XFILLER_0_47_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_163_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14715__Q team_03_WB.instance_to_wrap.core.decoder.inst\[12\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11441_ net2578 net395 _06760_ net499 vssd1 vssd1 vccd1 vccd1 _02047_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09876__B1_N net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08598__A1 net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14160_ clknet_leaf_161_wb_clk_i _01924_ _00525_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[514\]
+ sky130_fd_sc_hd__dfrtp_1
X_11372_ net507 net635 _06738_ net402 net2137 vssd1 vssd1 vccd1 vccd1 _02094_ sky130_fd_sc_hd__a32o_1
XANTENNA_clkbuf_leaf_3_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11777__S net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13111_ net1392 vssd1 vssd1 vccd1 vccd1 _00875_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_169_3839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10323_ _05968_ _05970_ _06127_ vssd1 vssd1 vccd1 vccd1 _06163_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07270__A1 net1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10944__A3 net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14091_ clknet_leaf_38_wb_clk_i _01855_ _00456_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[445\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_166_wb_clk_i clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_166_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_input53_A gpio_in[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13042_ net1397 vssd1 vssd1 vccd1 vccd1 _00806_ sky130_fd_sc_hd__inv_2
X_10254_ _03901_ _06095_ vssd1 vssd1 vccd1 vccd1 _06096_ sky130_fd_sc_hd__nand2_1
XANTENNA__08004__X _03946_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11354__B1 net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11078__A net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07022__A1 net1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1201 net1202 vssd1 vssd1 vccd1 vccd1 net1201 sky130_fd_sc_hd__clkbuf_4
Xfanout1212 net1213 vssd1 vssd1 vccd1 vccd1 net1212 sky130_fd_sc_hd__buf_4
X_10185_ _03430_ _06025_ vssd1 vssd1 vccd1 vccd1 _06027_ sky130_fd_sc_hd__nor2_1
Xfanout1223 net1224 vssd1 vssd1 vccd1 vccd1 net1223 sky130_fd_sc_hd__buf_4
XFILLER_0_56_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09193__D net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07990__S net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1234 net1235 vssd1 vssd1 vccd1 vccd1 net1234 sky130_fd_sc_hd__clkbuf_4
Xfanout1245 net1246 vssd1 vssd1 vccd1 vccd1 net1245 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11106__A0 _06519_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1256 net1264 vssd1 vssd1 vccd1 vccd1 net1256 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_31_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1267 net1278 vssd1 vssd1 vccd1 vccd1 net1267 sky130_fd_sc_hd__buf_4
Xfanout1278 net1438 vssd1 vssd1 vccd1 vccd1 net1278 sky130_fd_sc_hd__buf_2
X_14993_ clknet_leaf_10_wb_clk_i net41 _01358_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[12\]
+ sky130_fd_sc_hd__dfrtp_2
Xfanout280 _06409_ vssd1 vssd1 vccd1 vccd1 net280 sky130_fd_sc_hd__buf_2
Xfanout291 net294 vssd1 vssd1 vccd1 vccd1 net291 sky130_fd_sc_hd__clkbuf_4
XANTENNA__13293__A net1328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1289 net1302 vssd1 vssd1 vccd1 vccd1 net1289 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_89_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13944_ clknet_leaf_4_wb_clk_i _01708_ _00309_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[298\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08522__A1 net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07722__C net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13875_ clknet_leaf_105_wb_clk_i _01639_ _00240_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[229\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_158_203 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12826_ net1378 vssd1 vssd1 vccd1 vccd1 _00590_ sky130_fd_sc_hd__inv_2
XFILLER_0_69_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_258 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_735 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12757_ net1291 vssd1 vssd1 vccd1 vccd1 _00521_ sky130_fd_sc_hd__inv_2
XFILLER_0_84_543 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11708_ _06750_ net386 net340 net2433 vssd1 vssd1 vccd1 vccd1 _01826_ sky130_fd_sc_hd__a22o_1
X_12688_ net1412 vssd1 vssd1 vccd1 vccd1 _00452_ sky130_fd_sc_hd__inv_2
XFILLER_0_25_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08038__B1 net1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14427_ clknet_leaf_121_wb_clk_i _02191_ _00792_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[781\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06931__S1 net1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11639_ _06713_ net384 net348 net2132 vssd1 vssd1 vccd1 vccd1 _01893_ sky130_fd_sc_hd__a22o_1
XANTENNA__10157__A _03943_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08589__A1 net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_141_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14358_ clknet_leaf_152_wb_clk_i _02122_ _00723_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[712\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_170_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10396__A1 net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08850__A net1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11593__A0 net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold706 team_03_WB.instance_to_wrap.core.register_file.registers_state\[250\] vssd1
+ vssd1 vccd1 vccd1 net2199 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08684__S1 net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold717 team_03_WB.instance_to_wrap.core.register_file.registers_state\[473\] vssd1
+ vssd1 vccd1 vccd1 net2210 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10935__A3 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13309_ net1334 vssd1 vssd1 vccd1 vccd1 _01073_ sky130_fd_sc_hd__inv_2
XANTENNA__07261__A1 net1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold728 team_03_WB.instance_to_wrap.core.register_file.registers_state\[242\] vssd1
+ vssd1 vccd1 vccd1 net2221 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07737__Y _03679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14289_ clknet_leaf_143_wb_clk_i _02053_ _00654_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[643\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold739 team_03_WB.instance_to_wrap.core.register_file.registers_state\[897\] vssd1
+ vssd1 vccd1 vccd1 net2232 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_55_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09157__S net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10148__A1 _04207_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08850_ net1223 _04788_ _04789_ vssd1 vssd1 vccd1 vccd1 _04792_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_51_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11896__A1 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08761__A1 net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07801_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[171\] net775
+ net746 _03742_ vssd1 vssd1 vccd1 vccd1 _03743_ sky130_fd_sc_hd__o211a_1
X_08781_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[418\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[386\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[290\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[258\]
+ net977 net1080 vssd1 vssd1 vccd1 vccd1 _04723_ sky130_fd_sc_hd__mux4_1
XANTENNA__11138__D net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07732_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[781\] net800
+ _03673_ vssd1 vssd1 vccd1 vccd1 _03674_ sky130_fd_sc_hd__o21ai_1
XANTENNA__08297__A net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_95 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_140_3246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_3257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07663_ net1083 net888 team_03_WB.instance_to_wrap.core.register_file.registers_state\[30\]
+ vssd1 vssd1 vccd1 vccd1 _03605_ sky130_fd_sc_hd__o21a_1
X_09402_ _03641_ _05162_ net607 vssd1 vssd1 vccd1 vccd1 _05344_ sky130_fd_sc_hd__a21o_1
XFILLER_0_88_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11154__C _06478_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07594_ net1203 team_03_WB.instance_to_wrap.core.register_file.registers_state\[217\]
+ net786 team_03_WB.instance_to_wrap.core.register_file.registers_state\[249\] net752
+ vssd1 vssd1 vccd1 vccd1 _03536_ sky130_fd_sc_hd__o221a_1
XFILLER_0_149_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_61 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09333_ _05240_ _05274_ _05271_ vssd1 vssd1 vccd1 vccd1 _05275_ sky130_fd_sc_hd__or3b_2
XFILLER_0_47_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_3_7_0_wb_clk_i_X clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08277__B1 net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout338_A _06806_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_145_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09264_ _03682_ _05205_ vssd1 vssd1 vccd1 vccd1 _05206_ sky130_fd_sc_hd__xnor2_1
XANTENNA__11820__A1 net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_854 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_145_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11170__B _06503_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08215_ net855 _04155_ _04156_ _04154_ vssd1 vssd1 vccd1 vccd1 _04157_ sky130_fd_sc_hd__o31a_1
XANTENNA__08029__B1 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09195_ net544 _04825_ vssd1 vssd1 vccd1 vccd1 _05137_ sky130_fd_sc_hd__nor2_1
XANTENNA__10067__A net1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout505_A net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_145_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1247_A net1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_199 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08146_ _02799_ _02801_ _02810_ _02812_ net1073 vssd1 vssd1 vccd1 vccd1 _04088_ sky130_fd_sc_hd__a221o_2
XTAP_TAPCELL_ROW_116_2750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_2761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08760__A net1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11584__A0 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07788__C1 net1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_1908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11597__S net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_1919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07252__A1 net1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload160 clknet_leaf_103_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload160/X sky130_fd_sc_hd__clkbuf_8
X_08077_ net1090 team_03_WB.instance_to_wrap.core.register_file.registers_state\[886\]
+ net894 _04018_ net1130 vssd1 vssd1 vccd1 vccd1 _04019_ sky130_fd_sc_hd__o311a_1
Xclkload171 clknet_leaf_87_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload171/X sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout1035_X net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload182 clknet_leaf_100_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload182/Y sky130_fd_sc_hd__clkinv_2
XFILLER_0_101_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07028_ net1196 team_03_WB.instance_to_wrap.core.register_file.registers_state\[739\]
+ net884 _02969_ vssd1 vssd1 vccd1 vccd1 _02970_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_112_2669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout874_A net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout495_X net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11336__B1 net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_164_3736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10006__S net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11887__A1 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_164_3747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1202_X net1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold11 team_03_WB.instance_to_wrap.core.register_file.registers_state\[952\] vssd1
+ vssd1 vccd1 vccd1 net1504 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08752__A1 net1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold22 team_03_WB.instance_to_wrap.core.register_file.registers_state\[955\] vssd1
+ vssd1 vccd1 vccd1 net1515 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08752__B2 net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold33 team_03_WB.instance_to_wrap.ADR_I\[12\] vssd1 vssd1 vccd1 vccd1 net1526 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout662_X net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08979_ net869 _04920_ _04915_ vssd1 vssd1 vccd1 vccd1 _04921_ sky130_fd_sc_hd__o21ai_1
Xhold44 team_03_WB.instance_to_wrap.core.register_file.registers_state\[956\] vssd1
+ vssd1 vccd1 vccd1 net1537 sky130_fd_sc_hd__dlygate4sd3_1
Xhold55 team_03_WB.instance_to_wrap.core.register_file.registers_state\[962\] vssd1
+ vssd1 vccd1 vccd1 net1548 sky130_fd_sc_hd__dlygate4sd3_1
Xhold66 team_03_WB.instance_to_wrap.core.register_file.registers_state\[979\] vssd1
+ vssd1 vccd1 vccd1 net1559 sky130_fd_sc_hd__dlygate4sd3_1
Xhold77 team_03_WB.instance_to_wrap.core.register_file.registers_state\[999\] vssd1
+ vssd1 vccd1 vccd1 net1570 sky130_fd_sc_hd__dlygate4sd3_1
Xhold88 team_03_WB.instance_to_wrap.core.register_file.registers_state\[995\] vssd1
+ vssd1 vccd1 vccd1 net1581 sky130_fd_sc_hd__dlygate4sd3_1
X_11990_ net272 net2657 net444 vssd1 vssd1 vccd1 vccd1 _01554_ sky130_fd_sc_hd__mux2_1
Xhold99 team_03_WB.instance_to_wrap.core.register_file.registers_state\[967\] vssd1
+ vssd1 vccd1 vccd1 net1592 sky130_fd_sc_hd__dlygate4sd3_1
X_10941_ net689 net319 vssd1 vssd1 vccd1 vccd1 _06526_ sky130_fd_sc_hd__nand2_1
XANTENNA__11345__B net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout927_X net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_819 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13660_ clknet_leaf_148_wb_clk_i _01424_ _00025_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11064__C net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10872_ net494 net596 _06469_ net518 net1975 vssd1 vssd1 vccd1 vccd1 _02325_ sky130_fd_sc_hd__a32o_1
XFILLER_0_168_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12611_ net1374 vssd1 vssd1 vccd1 vccd1 _00375_ sky130_fd_sc_hd__inv_2
XFILLER_0_94_830 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13591_ net1343 vssd1 vssd1 vccd1 vccd1 _01355_ sky130_fd_sc_hd__inv_2
XFILLER_0_149_770 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11361__A net1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12542_ net1387 vssd1 vssd1 vccd1 vccd1 _00306_ sky130_fd_sc_hd__inv_2
XFILLER_0_137_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_442 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11080__B net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12473_ net1355 vssd1 vssd1 vccd1 vccd1 _00237_ sky130_fd_sc_hd__inv_2
X_14212_ clknet_leaf_29_wb_clk_i _01976_ _00577_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[566\]
+ sky130_fd_sc_hd__dfrtp_1
X_11424_ _06517_ _06751_ vssd1 vssd1 vccd1 vccd1 _06755_ sky130_fd_sc_hd__nor2_1
XFILLER_0_50_911 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07779__C1 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_495 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_8 net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13288__A net1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07243__A1 net1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14143_ clknet_leaf_170_wb_clk_i _01907_ _00508_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[497\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11355_ net274 net709 net695 vssd1 vssd1 vccd1 vccd1 _06730_ sky130_fd_sc_hd__and3_1
XANTENNA__11300__S net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10306_ team_03_WB.instance_to_wrap.core.pc.current_pc\[23\] team_03_WB.instance_to_wrap.core.pc.current_pc\[22\]
+ _06146_ vssd1 vssd1 vccd1 vccd1 _06148_ sky130_fd_sc_hd__and3_2
XFILLER_0_21_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08991__A1 net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14074_ clknet_leaf_145_wb_clk_i _01838_ _00439_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[428\]
+ sky130_fd_sc_hd__dfrtp_1
X_11286_ net509 net636 _06710_ net410 net2245 vssd1 vssd1 vccd1 vccd1 _02152_ sky130_fd_sc_hd__a32o_1
XANTENNA__11327__A0 net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13025_ net1261 vssd1 vssd1 vccd1 vccd1 _00789_ sky130_fd_sc_hd__inv_2
X_10237_ _03602_ _06078_ vssd1 vssd1 vccd1 vccd1 _06079_ sky130_fd_sc_hd__xnor2_1
XANTENNA__11878__A1 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12920__A net1376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11239__C _06413_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1020 net1022 vssd1 vssd1 vccd1 vccd1 net1020 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08743__A1 net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1031 net1032 vssd1 vssd1 vccd1 vccd1 net1031 sky130_fd_sc_hd__clkbuf_4
Xfanout1042 net1043 vssd1 vssd1 vccd1 vccd1 net1042 sky130_fd_sc_hd__clkbuf_4
X_10168_ team_03_WB.instance_to_wrap.core.pc.current_pc\[11\] net675 vssd1 vssd1 vccd1
+ vccd1 _06010_ sky130_fd_sc_hd__nand2_1
Xfanout1053 net1054 vssd1 vssd1 vccd1 vccd1 net1053 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_174_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11095__X _06624_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1064 net1069 vssd1 vssd1 vccd1 vccd1 net1064 sky130_fd_sc_hd__buf_4
XANTENNA__07951__C1 net1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08829__B _04770_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1075 net1080 vssd1 vssd1 vccd1 vccd1 net1075 sky130_fd_sc_hd__buf_4
XANTENNA__11536__A net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1086 net1093 vssd1 vssd1 vccd1 vccd1 net1086 sky130_fd_sc_hd__clkbuf_4
Xfanout1097 net1105 vssd1 vssd1 vccd1 vccd1 net1097 sky130_fd_sc_hd__clkbuf_4
X_14976_ clknet_leaf_88_wb_clk_i _02728_ _01341_ vssd1 vssd1 vccd1 vccd1 net228 sky130_fd_sc_hd__dfrtp_2
X_10099_ _02832_ net312 _05942_ vssd1 vssd1 vccd1 vccd1 _05943_ sky130_fd_sc_hd__or3b_1
XFILLER_0_117_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_63_wb_clk_i clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_63_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_117_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11255__B net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13927_ clknet_leaf_111_wb_clk_i _01691_ _00292_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[281\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07703__C1 net1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10853__A2 _05623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13858_ clknet_leaf_174_wb_clk_i _01622_ _00223_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[212\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12809_ net1254 vssd1 vssd1 vccd1 vccd1 _00573_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13789_ clknet_leaf_28_wb_clk_i _01553_ _00154_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[143\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11271__A net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09012__Y _04954_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_716 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11802__A1 net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_2008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15088__1474 vssd1 vssd1 vccd1 vccd1 _15088__1474/HI net1474 sky130_fd_sc_hd__conb_1
XFILLER_0_123_77 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09471__A2 net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_44_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07482__A1 net1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08000_ _03934_ _03941_ _03925_ vssd1 vssd1 vccd1 vccd1 _03942_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_96_2344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_96_2355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_142_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11566__B1 net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold503 team_03_WB.instance_to_wrap.core.register_file.registers_state\[428\] vssd1
+ vssd1 vccd1 vccd1 net1996 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold514 team_03_WB.instance_to_wrap.core.register_file.registers_state\[674\] vssd1
+ vssd1 vccd1 vccd1 net2007 sky130_fd_sc_hd__dlygate4sd3_1
Xhold525 team_03_WB.instance_to_wrap.core.register_file.registers_state\[285\] vssd1
+ vssd1 vccd1 vccd1 net2018 sky130_fd_sc_hd__dlygate4sd3_1
Xhold536 team_03_WB.instance_to_wrap.core.register_file.registers_state\[280\] vssd1
+ vssd1 vccd1 vccd1 net2029 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11210__S net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold547 team_03_WB.instance_to_wrap.core.register_file.registers_state\[679\] vssd1
+ vssd1 vccd1 vccd1 net2040 sky130_fd_sc_hd__dlygate4sd3_1
X_09951_ _03169_ net662 vssd1 vssd1 vccd1 vccd1 _05880_ sky130_fd_sc_hd__nor2_1
Xhold558 team_03_WB.instance_to_wrap.core.register_file.registers_state\[424\] vssd1
+ vssd1 vccd1 vccd1 net2051 sky130_fd_sc_hd__dlygate4sd3_1
Xhold569 team_03_WB.instance_to_wrap.core.register_file.registers_state\[759\] vssd1
+ vssd1 vccd1 vccd1 net2062 sky130_fd_sc_hd__dlygate4sd3_1
X_08902_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[428\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[396\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[300\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[268\]
+ net981 net1076 vssd1 vssd1 vccd1 vccd1 _04844_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_70_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09882_ _05596_ _05633_ _05823_ net315 vssd1 vssd1 vccd1 vccd1 _05824_ sky130_fd_sc_hd__or4b_1
XFILLER_0_110_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09082__S1 net1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07483__X _03425_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08734__A1 net1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08833_ _02953_ net573 vssd1 vssd1 vccd1 vccd1 _04775_ sky130_fd_sc_hd__nand2_2
Xhold1203 team_03_WB.instance_to_wrap.core.register_file.registers_state\[461\] vssd1
+ vssd1 vccd1 vccd1 net2696 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1214 team_03_WB.instance_to_wrap.core.register_file.registers_state\[159\] vssd1
+ vssd1 vccd1 vccd1 net2707 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1225 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[23\] vssd1 vssd1
+ vccd1 vccd1 net2718 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout288_A net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08739__B net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07942__C1 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1236 team_03_WB.instance_to_wrap.core.register_file.registers_state\[466\] vssd1
+ vssd1 vccd1 vccd1 net2729 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11446__A net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1247 team_03_WB.instance_to_wrap.core.register_file.registers_state\[195\] vssd1
+ vssd1 vccd1 vccd1 net2740 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12041__S net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08764_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[803\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[771\]
+ net980 vssd1 vssd1 vccd1 vccd1 _04706_ sky130_fd_sc_hd__mux2_1
Xhold1258 team_03_WB.instance_to_wrap.core.register_file.registers_state\[87\] vssd1
+ vssd1 vccd1 vccd1 net2751 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1269 team_03_WB.instance_to_wrap.core.register_file.registers_state\[215\] vssd1
+ vssd1 vccd1 vccd1 net2762 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07715_ net1104 team_03_WB.instance_to_wrap.core.register_file.registers_state\[301\]
+ net899 vssd1 vssd1 vccd1 vccd1 _03657_ sky130_fd_sc_hd__or3_1
X_08695_ net1241 team_03_WB.instance_to_wrap.core.register_file.registers_state\[200\]
+ net958 team_03_WB.instance_to_wrap.core.register_file.registers_state\[232\] net935
+ vssd1 vssd1 vccd1 vccd1 _04637_ sky130_fd_sc_hd__o221a_1
XFILLER_0_68_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout455_A net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1197_A net1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07646_ net1094 team_03_WB.instance_to_wrap.core.register_file.registers_state\[590\]
+ net796 team_03_WB.instance_to_wrap.core.register_file.registers_state\[622\] net746
+ vssd1 vssd1 vccd1 vccd1 _03588_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_68_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_146_Right_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10844__A2 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07577_ net1130 _03515_ _03516_ _03518_ vssd1 vssd1 vccd1 vccd1 _03519_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout622_A net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08474__B _04415_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1364_A net1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11181__A net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09316_ net572 _05257_ vssd1 vssd1 vccd1 vccd1 _05258_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10057__B1 net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09998__A0 net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_157_3595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_2801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09247_ _03428_ _05188_ vssd1 vssd1 vccd1 vccd1 _05189_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_35_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_173_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout410_X net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1152_X net1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_412 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout508_X net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_2709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07658__X _03600_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09178_ _05110_ _05113_ _05117_ _05119_ net555 net567 vssd1 vssd1 vccd1 vccd1 _05120_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout991_A net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08648__S1 net1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08921__C net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08129_ _04069_ _04070_ net610 vssd1 vssd1 vccd1 vccd1 _04071_ sky130_fd_sc_hd__mux2_2
XFILLER_0_121_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07225__A1 net1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11021__A2 net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_286 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08973__A1 net1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11140_ net1044 net837 net301 net668 vssd1 vssd1 vccd1 vccd1 _06646_ sky130_fd_sc_hd__and4_1
XFILLER_0_101_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09864__A2_N net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11309__A0 _06619_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout877_X net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11908__X _06814_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11071_ _06613_ net2738 net416 vssd1 vssd1 vccd1 vccd1 _02270_ sky130_fd_sc_hd__mux2_1
XANTENNA__11059__C net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput101 wbs_stb_i vssd1 vssd1 vccd1 vccd1 net101 sky130_fd_sc_hd__clkbuf_1
XANTENNA__08725__A1 net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10022_ net84 net83 net86 net85 vssd1 vssd1 vccd1 vccd1 _05900_ sky130_fd_sc_hd__or4_1
XFILLER_0_76_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14830_ clknet_leaf_84_wb_clk_i net1596 _01195_ vssd1 vssd1 vccd1 vccd1 net151 sky130_fd_sc_hd__dfrtp_1
XANTENNA_input16_A DAT_I[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14761_ clknet_leaf_49_wb_clk_i _02525_ _01126_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_11973_ net642 _06750_ net477 net365 net2166 vssd1 vssd1 vccd1 vccd1 _01570_ sky130_fd_sc_hd__a32o_1
XANTENNA__11790__S net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11643__X _06805_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10924_ team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[9\] net312 _05845_ net318
+ vssd1 vssd1 vccd1 vccd1 _06512_ sky130_fd_sc_hd__and4_1
X_13712_ clknet_leaf_157_wb_clk_i _01476_ _00077_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[66\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14692_ clknet_leaf_59_wb_clk_i _02456_ _01057_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.ADR_I\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_113_Right_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07700__A2 net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_375 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12037__A1 net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13643_ net1424 vssd1 vssd1 vccd1 vccd1 _01407_ sky130_fd_sc_hd__inv_2
X_10855_ net833 net274 vssd1 vssd1 vccd1 vccd1 _06454_ sky130_fd_sc_hd__and2_2
XFILLER_0_116_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10048__B1 net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11091__A net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13574_ net1432 vssd1 vssd1 vccd1 vccd1 _01338_ sky130_fd_sc_hd__inv_2
XFILLER_0_94_682 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10786_ net311 net310 net317 vssd1 vssd1 vccd1 vccd1 _06396_ sky130_fd_sc_hd__and3_2
XANTENNA__11522__C net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12525_ net1311 vssd1 vssd1 vccd1 vccd1 _00289_ sky130_fd_sc_hd__inv_2
XFILLER_0_147_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_181_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_181_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__11241__D net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08661__B1 net1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_423 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_922 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12456_ net1290 vssd1 vssd1 vccd1 vccd1 _00220_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_1019 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08604__S net992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_110_wb_clk_i clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_110_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_2_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_151_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11407_ net301 net2330 net396 vssd1 vssd1 vccd1 vccd1 _02073_ sky130_fd_sc_hd__mux2_1
XANTENNA__11012__A2 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12387_ net1371 vssd1 vssd1 vccd1 vccd1 _00151_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14126_ clknet_leaf_131_wb_clk_i _01890_ _00491_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[480\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_91_2241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11338_ net499 net627 _06721_ net401 net1980 vssd1 vssd1 vccd1 vccd1 _02111_ sky130_fd_sc_hd__a32o_1
XFILLER_0_22_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_91_2252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14057_ clknet_leaf_75_wb_clk_i _01821_ _00422_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[411\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09943__B net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11269_ net713 net271 net831 vssd1 vssd1 vccd1 vccd1 _06702_ sky130_fd_sc_hd__and3_1
XFILLER_0_24_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08716__A1 net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09435__S net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_37 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13008_ net1410 vssd1 vssd1 vccd1 vccd1 _00772_ sky130_fd_sc_hd__inv_2
XANTENNA__10170__A _03758_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14959_ clknet_leaf_83_wb_clk_i _02711_ _01324_ vssd1 vssd1 vccd1 vccd1 net211 sky130_fd_sc_hd__dfrtp_1
XANTENNA__10287__A0 _04475_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07500_ net1109 team_03_WB.instance_to_wrap.core.register_file.registers_state\[39\]
+ net901 vssd1 vssd1 vccd1 vccd1 _03442_ sky130_fd_sc_hd__or3_1
XFILLER_0_159_320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10826__A2 _06429_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08480_ net1242 team_03_WB.instance_to_wrap.core.register_file.registers_state\[731\]
+ net987 team_03_WB.instance_to_wrap.core.register_file.registers_state\[763\] net945
+ vssd1 vssd1 vccd1 vccd1 _04422_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_46_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07431_ net1147 _03362_ _03372_ vssd1 vssd1 vccd1 vccd1 _03373_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_147_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_159_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_147_548 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11205__S net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07362_ net1138 _03301_ _03302_ vssd1 vssd1 vccd1 vccd1 _03304_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_63_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_21_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08101__C1 net1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_170 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_28_Left_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_21_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09101_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[46\] net976
+ vssd1 vssd1 vccd1 vccd1 _05043_ sky130_fd_sc_hd__or2_1
XFILLER_0_31_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_165_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_135_3145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07455__A1 net1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_3156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07293_ net1108 team_03_WB.instance_to_wrap.core.register_file.registers_state\[489\]
+ net902 vssd1 vssd1 vccd1 vccd1 _03235_ sky130_fd_sc_hd__or3_1
XFILLER_0_5_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09032_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[560\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[528\]
+ net984 vssd1 vssd1 vccd1 vccd1 _04974_ sky130_fd_sc_hd__mux2_1
XFILLER_0_142_231 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_152_3492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold300 team_03_WB.instance_to_wrap.core.register_file.registers_state\[60\] vssd1
+ vssd1 vccd1 vccd1 net1793 sky130_fd_sc_hd__dlygate4sd3_1
Xhold311 _02618_ vssd1 vssd1 vccd1 vccd1 net1804 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold322 team_03_WB.instance_to_wrap.core.register_file.registers_state\[3\] vssd1
+ vssd1 vccd1 vccd1 net1815 sky130_fd_sc_hd__dlygate4sd3_1
Xhold333 net222 vssd1 vssd1 vccd1 vccd1 net1826 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08955__A1 net1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold344 team_03_WB.instance_to_wrap.CPU_DAT_I\[26\] vssd1 vssd1 vccd1 vccd1 net1837
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08955__B2 net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold355 team_03_WB.instance_to_wrap.ADR_I\[30\] vssd1 vssd1 vccd1 vccd1 net1848 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold366 team_03_WB.instance_to_wrap.core.register_file.registers_state\[47\] vssd1
+ vssd1 vccd1 vccd1 net1859 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06966__B1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10064__B team_03_WB.instance_to_wrap.core.decoder.inst\[10\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold377 team_03_WB.instance_to_wrap.core.register_file.registers_state\[386\] vssd1
+ vssd1 vccd1 vccd1 net1870 sky130_fd_sc_hd__dlygate4sd3_1
Xhold388 team_03_WB.instance_to_wrap.core.register_file.registers_state\[805\] vssd1
+ vssd1 vccd1 vccd1 net1881 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout802 net805 vssd1 vssd1 vccd1 vccd1 net802 sky130_fd_sc_hd__clkbuf_4
X_09934_ _05871_ net1883 net293 vssd1 vssd1 vccd1 vccd1 _02760_ sky130_fd_sc_hd__mux2_1
Xhold399 team_03_WB.instance_to_wrap.core.register_file.registers_state\[387\] vssd1
+ vssd1 vccd1 vccd1 net1892 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1026 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06969__S net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout813 net816 vssd1 vssd1 vccd1 vccd1 net813 sky130_fd_sc_hd__buf_4
XANTENNA_fanout1112_A net1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout824 net825 vssd1 vssd1 vccd1 vccd1 net824 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_110_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_37_Left_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout835 _06387_ vssd1 vssd1 vccd1 vccd1 net835 sky130_fd_sc_hd__clkbuf_2
XANTENNA__10999__B net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout846 net847 vssd1 vssd1 vccd1 vccd1 net846 sky130_fd_sc_hd__buf_4
XANTENNA__07654__A net1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09865_ _03947_ net535 net590 _03944_ _02804_ vssd1 vssd1 vccd1 vccd1 _05807_ sky130_fd_sc_hd__o32ai_2
Xfanout857 net858 vssd1 vssd1 vccd1 vccd1 net857 sky130_fd_sc_hd__clkbuf_8
XANTENNA_input8_A DAT_I[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1000 team_03_WB.instance_to_wrap.core.register_file.registers_state\[855\] vssd1
+ vssd1 vccd1 vccd1 net2493 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout572_A _03024_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout868 net870 vssd1 vssd1 vccd1 vccd1 net868 sky130_fd_sc_hd__buf_4
Xfanout879 net887 vssd1 vssd1 vccd1 vccd1 net879 sky130_fd_sc_hd__buf_2
Xhold1011 team_03_WB.instance_to_wrap.core.register_file.registers_state\[528\] vssd1
+ vssd1 vccd1 vccd1 net2504 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11176__A net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1022 team_03_WB.instance_to_wrap.core.register_file.registers_state\[490\] vssd1
+ vssd1 vccd1 vccd1 net2515 sky130_fd_sc_hd__dlygate4sd3_1
X_08816_ net1221 _04755_ vssd1 vssd1 vccd1 vccd1 _04758_ sky130_fd_sc_hd__or2_1
Xhold1033 team_03_WB.instance_to_wrap.core.register_file.registers_state\[512\] vssd1
+ vssd1 vccd1 vccd1 net2526 sky130_fd_sc_hd__dlygate4sd3_1
X_09796_ _05113_ _05130_ net555 vssd1 vssd1 vccd1 vccd1 _05738_ sky130_fd_sc_hd__mux2_1
Xhold1044 team_03_WB.instance_to_wrap.core.register_file.registers_state\[143\] vssd1
+ vssd1 vccd1 vccd1 net2537 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1055 team_03_WB.instance_to_wrap.core.register_file.registers_state\[202\] vssd1
+ vssd1 vccd1 vccd1 net2548 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1066 team_03_WB.instance_to_wrap.core.register_file.registers_state\[84\] vssd1
+ vssd1 vccd1 vccd1 net2559 sky130_fd_sc_hd__dlygate4sd3_1
X_08747_ net1052 team_03_WB.instance_to_wrap.core.register_file.registers_state\[451\]
+ net1005 team_03_WB.instance_to_wrap.core.register_file.registers_state\[483\] net1076
+ vssd1 vssd1 vccd1 vccd1 _04689_ sky130_fd_sc_hd__a221o_1
Xhold1077 team_03_WB.instance_to_wrap.core.register_file.registers_state\[729\] vssd1
+ vssd1 vccd1 vccd1 net2570 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_107_2568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout360_X net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1088 team_03_WB.instance_to_wrap.core.register_file.registers_state\[448\] vssd1
+ vssd1 vccd1 vccd1 net2581 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1099 team_03_WB.instance_to_wrap.core.register_file.registers_state\[584\] vssd1
+ vssd1 vccd1 vccd1 net2592 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_107_2579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout837_A _06386_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout458_X net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09132__B2 _05073_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_936 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08678_ _04619_ vssd1 vssd1 vccd1 vccd1 _04620_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_159_3635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07143__B1 net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_159_3646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08340__C1 net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_165_301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07629_ net1192 team_03_WB.instance_to_wrap.core.register_file.registers_state\[142\]
+ net881 net1154 vssd1 vssd1 vccd1 vccd1 _03571_ sky130_fd_sc_hd__o211a_1
XANTENNA__12019__A1 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout625_X net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11115__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1367_X net1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_46_Left_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10640_ net1162 net2736 net844 vssd1 vssd1 vccd1 vccd1 _02488_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_165_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_924 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10571_ net1711 net534 net601 _05881_ vssd1 vssd1 vccd1 vccd1 _02552_ sky130_fd_sc_hd__a22o_1
XANTENNA__11242__A2 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11061__D net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12310_ net1280 vssd1 vssd1 vccd1 vccd1 _00074_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07829__A net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13290_ net1327 vssd1 vssd1 vccd1 vccd1 _01054_ sky130_fd_sc_hd__inv_2
XFILLER_0_134_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_184 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout994_X net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09199__A1 _05073_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09199__B2 _04777_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12241_ net1777 vssd1 vssd1 vccd1 vccd1 _01416_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__10255__A _03901_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08946__A1 net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12172_ net1605 vssd1 vssd1 vccd1 vccd1 _02381_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__08946__B2 net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07267__C net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11950__B1 net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11785__S net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11123_ net2659 net412 _06636_ net492 vssd1 vssd1 vccd1 vccd1 _02241_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_55_Left_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11054_ net511 net656 _06604_ net422 net2009 vssd1 vssd1 vccd1 vccd1 _02278_ sky130_fd_sc_hd__a32o_1
X_15087__1473 vssd1 vssd1 vccd1 vccd1 _15087__1473/HI net1473 sky130_fd_sc_hd__conb_1
XANTENNA__10505__A1 net114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11702__B1 net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10005_ _05890_ net2491 net287 vssd1 vssd1 vccd1 vccd1 _02709_ sky130_fd_sc_hd__mux2_1
X_14813_ clknet_leaf_94_wb_clk_i net1623 _01178_ vssd1 vssd1 vccd1 vccd1 net164 sky130_fd_sc_hd__dfrtp_1
XANTENNA_input19_X net19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14744_ clknet_leaf_49_wb_clk_i _02508_ _01109_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_114_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_28_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_104 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11956_ net624 _06733_ net455 net363 net2224 vssd1 vssd1 vccd1 vccd1 _01587_ sky130_fd_sc_hd__a32o_1
XANTENNA__06908__A net1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10907_ team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[12\] net311 net310 net317
+ vssd1 vssd1 vccd1 vccd1 _06498_ sky130_fd_sc_hd__and4_1
XANTENNA__07685__A1 net1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14675_ clknet_leaf_87_wb_clk_i _02439_ _01040_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.ADR_I\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_11887_ net622 _06696_ net455 net371 net2253 vssd1 vssd1 vccd1 vccd1 _01654_ sky130_fd_sc_hd__a32o_1
XANTENNA__07685__B2 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10838_ net313 net309 net316 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[22\]
+ vssd1 vssd1 vccd1 vccd1 _06439_ sky130_fd_sc_hd__o31a_1
X_13626_ net1415 vssd1 vssd1 vccd1 vccd1 _01390_ sky130_fd_sc_hd__inv_2
XFILLER_0_156_367 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10149__B _05990_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11769__B1 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07437__A1 net1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10769_ net525 _06378_ _06379_ net530 net1599 vssd1 vssd1 vccd1 vccd1 _02434_ sky130_fd_sc_hd__a32o_1
X_13557_ net1432 vssd1 vssd1 vccd1 vccd1 _01321_ sky130_fd_sc_hd__inv_2
XFILLER_0_13_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12508_ net1409 vssd1 vssd1 vccd1 vccd1 _00272_ sky130_fd_sc_hd__inv_2
X_13488_ net1344 vssd1 vssd1 vccd1 vccd1 _01252_ sky130_fd_sc_hd__inv_2
XFILLER_0_152_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08334__S net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_59 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12439_ net1390 vssd1 vssd1 vccd1 vccd1 _00203_ sky130_fd_sc_hd__inv_2
XANTENNA__10165__A _03724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_3042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_763 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_130_3053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06930__X _02872_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_39_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07070__C1 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14109_ clknet_leaf_25_wb_clk_i _01873_ _00474_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[463\]
+ sky130_fd_sc_hd__dfrtp_1
X_15089_ net1475 vssd1 vssd1 vccd1 vccd1 la_data_out[25] sky130_fd_sc_hd__buf_2
XANTENNA__09673__B _05570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07980_ net1106 team_03_WB.instance_to_wrap.core.register_file.registers_state\[304\]
+ net901 vssd1 vssd1 vccd1 vccd1 _03922_ sky130_fd_sc_hd__or3_1
XFILLER_0_129_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06931_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[420\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[388\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[292\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[260\]
+ net781 net1136 vssd1 vssd1 vccd1 vccd1 _02873_ sky130_fd_sc_hd__mux4_1
XANTENNA__07905__C net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09650_ _05356_ _05547_ _05589_ _05591_ vssd1 vssd1 vccd1 vccd1 _05592_ sky130_fd_sc_hd__o211a_1
XANTENNA__08796__S0 net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06862_ _02799_ _02801_ vssd1 vssd1 vccd1 vccd1 _02804_ sky130_fd_sc_hd__nand2_8
XFILLER_0_98_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11427__C _06463_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08601_ net1059 team_03_WB.instance_to_wrap.core.register_file.registers_state\[677\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[645\] net1011 net946
+ vssd1 vssd1 vccd1 vccd1 _04543_ sky130_fd_sc_hd__o221a_1
XFILLER_0_59_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09581_ _05521_ _05522_ net576 vssd1 vssd1 vccd1 vccd1 _05523_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_1098 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08532_ _04468_ _04473_ net871 vssd1 vssd1 vccd1 vccd1 _04474_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_26_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_65_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08463_ net1227 team_03_WB.instance_to_wrap.core.register_file.registers_state\[92\]
+ net953 team_03_WB.instance_to_wrap.core.register_file.registers_state\[124\] net917
+ vssd1 vssd1 vccd1 vccd1 _04405_ sky130_fd_sc_hd__o221a_1
XFILLER_0_93_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11472__A2 net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_102_2465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07414_ net726 _03353_ _03354_ net1115 vssd1 vssd1 vccd1 vccd1 _03356_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_102_2476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11162__C net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_833 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08394_ net1244 team_03_WB.instance_to_wrap.core.register_file.registers_state\[473\]
+ net991 team_03_WB.instance_to_wrap.core.register_file.registers_state\[505\] net1216
+ vssd1 vssd1 vccd1 vccd1 _04336_ sky130_fd_sc_hd__o221a_1
XFILLER_0_169_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_154_3532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_154_3543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07345_ net1083 team_03_WB.instance_to_wrap.core.register_file.registers_state\[252\]
+ net891 vssd1 vssd1 vccd1 vccd1 _03287_ sky130_fd_sc_hd__or3_1
XFILLER_0_46_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_174_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1062_A net1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout418_A _06610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07979__A2 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09200__Y _05142_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07276_ net1201 team_03_WB.instance_to_wrap.core.register_file.registers_state\[585\]
+ net784 team_03_WB.instance_to_wrap.core.register_file.registers_state\[617\] net734
+ vssd1 vssd1 vccd1 vccd1 _03218_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_171_3890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09015_ _04895_ _04956_ net558 vssd1 vssd1 vccd1 vccd1 _04957_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1327_A net1328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08389__C1 net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold130 _02577_ vssd1 vssd1 vccd1 vccd1 net1623 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold141 net122 vssd1 vssd1 vccd1 vccd1 net1634 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_37_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__07087__C net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold152 _02576_ vssd1 vssd1 vccd1 vccd1 net1645 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11932__A0 _06519_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold163 team_03_WB.instance_to_wrap.CPU_DAT_I\[19\] vssd1 vssd1 vccd1 vccd1 net1656
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout787_A net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold174 _02573_ vssd1 vssd1 vccd1 vccd1 net1667 sky130_fd_sc_hd__dlygate4sd3_1
Xhold185 _02629_ vssd1 vssd1 vccd1 vccd1 net1678 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07600__A1 net1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12290__A net1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout610 net611 vssd1 vssd1 vccd1 vccd1 net610 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_111_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1115_X net1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold196 net183 vssd1 vssd1 vccd1 vccd1 net1689 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout621 net631 vssd1 vssd1 vccd1 vccd1 net621 sky130_fd_sc_hd__clkbuf_2
X_09917_ _05082_ _05852_ _05858_ vssd1 vssd1 vccd1 vccd1 _05859_ sky130_fd_sc_hd__or3_1
Xfanout632 net634 vssd1 vssd1 vccd1 vccd1 net632 sky130_fd_sc_hd__clkbuf_4
Xfanout643 net644 vssd1 vssd1 vccd1 vccd1 net643 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_109_2608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_2619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout654 net655 vssd1 vssd1 vccd1 vccd1 net654 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout954_A net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout665 net666 vssd1 vssd1 vccd1 vccd1 net665 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__10499__B1 net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout676 _05948_ vssd1 vssd1 vccd1 vccd1 net676 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_77_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout687 _02840_ vssd1 vssd1 vccd1 vccd1 net687 sky130_fd_sc_hd__clkbuf_4
X_09848_ net537 _05787_ _05789_ vssd1 vssd1 vccd1 vccd1 _05790_ sky130_fd_sc_hd__o21a_1
XANTENNA__11337__C _06413_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07364__B1 net1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout698 net700 vssd1 vssd1 vccd1 vccd1 net698 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_38_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_126_2955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10949__S net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout742_X net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09779_ _04649_ _04956_ net562 vssd1 vssd1 vccd1 vccd1 _05721_ sky130_fd_sc_hd__mux2_1
XANTENNA__09105__A1 net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11810_ _06636_ net451 net323 net2357 vssd1 vssd1 vccd1 vccd1 _01729_ sky130_fd_sc_hd__a22o_1
X_12790_ net1280 vssd1 vssd1 vccd1 vccd1 _00554_ sky130_fd_sc_hd__inv_2
XFILLER_0_96_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14718__Q team_03_WB.instance_to_wrap.core.decoder.inst\[15\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11353__B net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11741_ net1989 net267 net336 vssd1 vssd1 vccd1 vccd1 _01795_ sky130_fd_sc_hd__mux2_1
XANTENNA__07667__A1 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11463__A2 net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07550__C net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11672_ net2663 _06631_ net345 vssd1 vssd1 vccd1 vccd1 _01861_ sky130_fd_sc_hd__mux2_1
X_14460_ clknet_leaf_150_wb_clk_i _02224_ _00825_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[814\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_153_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_166_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10623_ net1560 team_03_WB.instance_to_wrap.CPU_DAT_O\[6\] net842 vssd1 vssd1 vccd1
+ vccd1 _02505_ sky130_fd_sc_hd__mux2_1
XANTENNA__07419__A1 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13411_ net1416 vssd1 vssd1 vccd1 vccd1 _01175_ sky130_fd_sc_hd__inv_2
XFILLER_0_107_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14391_ clknet_leaf_113_wb_clk_i _02155_ _00756_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[745\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_4_12__f_wb_clk_i_A clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_76_wb_clk_i_A clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_994 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13342_ net1342 vssd1 vssd1 vccd1 vccd1 _01106_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10554_ team_03_WB.instance_to_wrap.BUSY_O team_03_WB.instance_to_wrap.core.ru.state\[5\]
+ net606 net1145 vssd1 vssd1 vccd1 vccd1 _06297_ sky130_fd_sc_hd__a22o_1
XANTENNA_input83_A wbs_adr_i[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1057 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10974__A1 net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13273_ net1423 vssd1 vssd1 vccd1 vccd1 _01037_ sky130_fd_sc_hd__inv_2
XFILLER_0_121_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10485_ net1902 net1027 net905 team_03_WB.instance_to_wrap.ADR_I\[21\] vssd1 vssd1
+ vccd1 vccd1 _02624_ sky130_fd_sc_hd__a22o_1
XFILLER_0_134_595 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08919__A1 net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07846__X _03788_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15012_ clknet_leaf_10_wb_clk_i net60 _01377_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[31\]
+ sky130_fd_sc_hd__dfrtp_2
X_12224_ net1591 vssd1 vssd1 vccd1 vccd1 _01433_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__10726__A1 net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11923__A0 _06479_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13296__A net1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12155_ net1632 vssd1 vssd1 vccd1 vccd1 _02398_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_102_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06910__B net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07294__A net1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11106_ _06519_ net2484 net418 vssd1 vssd1 vccd1 vccd1 _02250_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12086_ net622 _06652_ net454 net439 net1817 vssd1 vssd1 vccd1 vccd1 _01461_ sky130_fd_sc_hd__a32o_1
X_11037_ net2404 net422 _06594_ net503 vssd1 vssd1 vccd1 vccd1 _02285_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_34_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11151__A1 net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08677__X _04619_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11247__C net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07355__B1 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08552__C1 net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06909__Y _02851_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11544__A net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08329__S net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07107__B1 net1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09647__A2 _02804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12100__B1 net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12988_ net1418 vssd1 vssd1 vccd1 vccd1 _00752_ sky130_fd_sc_hd__inv_2
XANTENNA__08304__C1 net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11263__B net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_2059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14727_ clknet_leaf_48_wb_clk_i _02491_ _01092_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.decoder.inst\[24\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_59_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11454__A2 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07658__B2 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11939_ _06632_ net2775 net369 vssd1 vssd1 vccd1 vccd1 _01603_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_107 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09949__A _03136_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14658_ clknet_leaf_176_wb_clk_i _02422_ _01023_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1012\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_60_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_145_827 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13609_ net1340 vssd1 vssd1 vccd1 vccd1 _01373_ sky130_fd_sc_hd__inv_2
XFILLER_0_145_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14589_ clknet_leaf_165_wb_clk_i _02353_ _00954_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[943\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_54_151 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07130_ net1198 team_03_WB.instance_to_wrap.core.register_file.registers_state\[608\]
+ net885 _03071_ vssd1 vssd1 vccd1 vccd1 _03072_ sky130_fd_sc_hd__a31o_1
XANTENNA__07469__A net1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11757__A3 net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_wire588_A _05068_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_153_882 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07061_ net1097 team_03_WB.instance_to_wrap.core.register_file.registers_state\[706\]
+ net797 team_03_WB.instance_to_wrap.core.register_file.registers_state\[738\] vssd1
+ vssd1 vccd1 vccd1 _03003_ sky130_fd_sc_hd__a22o_1
XANTENNA__07830__A1 net1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09955__Y _05882_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08999__S net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_908 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput202 net202 vssd1 vssd1 vccd1 vccd1 gpio_oeb[6] sky130_fd_sc_hd__buf_2
Xoutput213 net213 vssd1 vssd1 vccd1 vccd1 gpio_out[16] sky130_fd_sc_hd__buf_2
XFILLER_0_3_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput224 net224 vssd1 vssd1 vccd1 vccd1 gpio_out[27] sky130_fd_sc_hd__clkbuf_4
XANTENNA__10717__A1 net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput235 net235 vssd1 vssd1 vccd1 vccd1 gpio_out[7] sky130_fd_sc_hd__buf_2
XFILLER_0_2_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_58_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput246 net246 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[18] sky130_fd_sc_hd__buf_2
Xoutput257 net914 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[31] sky130_fd_sc_hd__buf_2
XANTENNA__09583__A1 net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11390__A1 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07594__B1 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08791__C1 net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11438__B net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07963_ net1107 net903 team_03_WB.instance_to_wrap.core.register_file.registers_state\[16\]
+ vssd1 vssd1 vccd1 vccd1 _03905_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_147_3391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09702_ _05073_ _05506_ _05638_ _04777_ _05643_ vssd1 vssd1 vccd1 vccd1 _05644_ sky130_fd_sc_hd__a221o_1
XFILLER_0_4_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06914_ net1106 team_03_WB.instance_to_wrap.core.register_file.registers_state\[36\]
+ net903 vssd1 vssd1 vccd1 vccd1 _02856_ sky130_fd_sc_hd__or3_1
X_07894_ net1091 team_03_WB.instance_to_wrap.core.register_file.registers_state\[463\]
+ vssd1 vssd1 vccd1 vccd1 _03836_ sky130_fd_sc_hd__and2_1
XANTENNA__11157__C net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08543__C1 net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11142__B2 net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07932__A net1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09633_ net584 _04775_ _05570_ _05573_ _05574_ vssd1 vssd1 vccd1 vccd1 _05575_ sky130_fd_sc_hd__o311a_1
X_06845_ net1208 vssd1 vssd1 vccd1 vccd1 _02788_ sky130_fd_sc_hd__inv_2
XANTENNA__07897__A1 net1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11693__A2 net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout270_A _06509_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_2505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout368_A _06814_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_2516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09564_ _04269_ _04386_ _04448_ _04534_ net559 net564 vssd1 vssd1 vccd1 vccd1 _05506_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_clkbuf_4_8__f_wb_clk_i_A clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08515_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[831\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[799\]
+ net952 vssd1 vssd1 vccd1 vccd1 _04457_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_110_wb_clk_i_A clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11173__B net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09495_ _05377_ _05381_ net567 vssd1 vssd1 vccd1 vccd1 _05437_ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_121_2852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11445__A2 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08846__B1 net1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_2863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_714 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout535_A net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1277_A net1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09859__A _05730_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08446_ net1228 team_03_WB.instance_to_wrap.core.register_file.registers_state\[604\]
+ net953 team_03_WB.instance_to_wrap.core.register_file.registers_state\[636\] net917
+ vssd1 vssd1 vccd1 vccd1 _04388_ sky130_fd_sc_hd__o221a_1
XFILLER_0_148_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_173_3930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08763__A net1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_162_112 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08377_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[1014\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[982\]
+ net970 vssd1 vssd1 vccd1 vccd1 _04319_ sky130_fd_sc_hd__mux2_1
XFILLER_0_147_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout323_X net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1065_X net1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15086__1472 vssd1 vssd1 vccd1 vccd1 _15086__1472/HI net1472 sky130_fd_sc_hd__conb_1
XFILLER_0_33_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07379__A net1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07328_ net1182 team_03_WB.instance_to_wrap.core.register_file.registers_state\[349\]
+ net768 team_03_WB.instance_to_wrap.core.register_file.registers_state\[381\] net1128
+ vssd1 vssd1 vccd1 vccd1 _03270_ sky130_fd_sc_hd__o221a_1
XANTENNA__08074__A1 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09810__A2 _04565_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07259_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[424\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[392\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[296\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[264\]
+ net774 net1131 vssd1 vssd1 vccd1 vccd1 _03201_ sky130_fd_sc_hd__mux4_1
XFILLER_0_5_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10009__S net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1232_X net1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09594__A net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10270_ _05975_ _06111_ vssd1 vssd1 vccd1 vccd1 _06112_ sky130_fd_sc_hd__and2_1
XANTENNA__09023__B1 net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11905__B1 net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09574__A1 net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11188__X _06675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1405 net1408 vssd1 vssd1 vccd1 vccd1 net1405 sky130_fd_sc_hd__buf_2
Xfanout1416 net1417 vssd1 vssd1 vccd1 vccd1 net1416 sky130_fd_sc_hd__buf_4
Xfanout1427 net1429 vssd1 vssd1 vccd1 vccd1 net1427 sky130_fd_sc_hd__buf_4
XANTENNA__08003__A net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout440 _06819_ vssd1 vssd1 vccd1 vccd1 net440 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout957_X net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1438 net66 vssd1 vssd1 vccd1 vccd1 net1438 sky130_fd_sc_hd__buf_4
Xfanout451 net453 vssd1 vssd1 vccd1 vccd1 net451 sky130_fd_sc_hd__buf_4
Xfanout462 net463 vssd1 vssd1 vccd1 vccd1 net462 sky130_fd_sc_hd__buf_4
X_13960_ clknet_leaf_13_wb_clk_i _01724_ _00325_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[314\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout473 net476 vssd1 vssd1 vccd1 vccd1 net473 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07337__B1 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout484 _06779_ vssd1 vssd1 vccd1 vccd1 net484 sky130_fd_sc_hd__clkbuf_8
XANTENNA__11133__B2 net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout495 net496 vssd1 vssd1 vccd1 vccd1 net495 sky130_fd_sc_hd__clkbuf_4
X_12911_ net1394 vssd1 vssd1 vccd1 vccd1 _00675_ sky130_fd_sc_hd__inv_2
XANTENNA__07888__A1 net1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11684__A2 net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13891_ clknet_leaf_35_wb_clk_i _01655_ _00256_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[245\]
+ sky130_fd_sc_hd__dfrtp_1
X_12842_ net1283 vssd1 vssd1 vccd1 vccd1 _00606_ sky130_fd_sc_hd__inv_2
XFILLER_0_150_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_17_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_1016 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12773_ net1351 vssd1 vssd1 vccd1 vccd1 _00537_ sky130_fd_sc_hd__inv_2
XANTENNA__10644__A0 net1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14512_ clknet_leaf_156_wb_clk_i _02276_ _00877_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[866\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08932__S0 net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11724_ net1952 net273 net335 vssd1 vssd1 vccd1 vccd1 _01812_ sky130_fd_sc_hd__mux2_1
X_14443_ clknet_leaf_45_wb_clk_i _02207_ _00808_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[797\]
+ sky130_fd_sc_hd__dfrtp_1
X_11655_ net2630 _06454_ net342 vssd1 vssd1 vccd1 vccd1 _01878_ sky130_fd_sc_hd__mux2_1
XANTENNA__06905__B net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11303__S net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_668 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_88_wb_clk_i clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_88_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_10606_ net2718 net1961 net840 vssd1 vssd1 vccd1 vccd1 _02522_ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11586_ net275 net2477 net448 vssd1 vssd1 vccd1 vccd1 _01943_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07499__S0 net1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14374_ clknet_leaf_27_wb_clk_i _02138_ _00739_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[728\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_153_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10947__A1 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13325_ net1318 vssd1 vssd1 vccd1 vccd1 _01089_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_17_wb_clk_i clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_17_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_10537_ net158 net1034 net1026 net1666 vssd1 vssd1 vccd1 vccd1 _02573_ sky130_fd_sc_hd__a22o_1
XANTENNA__07812__B2 net1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1086 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10468_ team_03_WB.instance_to_wrap.core.pc.current_pc\[2\] _06280_ net683 vssd1
+ vssd1 vccd1 vccd1 _02636_ sky130_fd_sc_hd__mux2_1
X_13256_ net1298 vssd1 vssd1 vccd1 vccd1 _01020_ sky130_fd_sc_hd__inv_2
XANTENNA__06921__A team_03_WB.instance_to_wrap.core.decoder.inst\[24\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12207_ net1511 vssd1 vssd1 vccd1 vccd1 _02346_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_36_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13187_ net1354 vssd1 vssd1 vccd1 vccd1 _00951_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_36_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10399_ _06004_ _06069_ _06079_ _06078_ _03602_ vssd1 vssd1 vccd1 vccd1 _06225_ sky130_fd_sc_hd__o32a_1
XANTENNA__11372__A1 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07228__S net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09009__A net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12138_ net1577 vssd1 vssd1 vccd1 vccd1 _02415_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_53_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09951__B net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12069_ _06631_ net2700 net357 vssd1 vssd1 vccd1 vccd1 _01477_ sky130_fd_sc_hd__mux2_1
XANTENNA__07328__B1 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09443__S net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_1085 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07752__A net1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07879__A1 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10635__A0 team_03_WB.instance_to_wrap.core.decoder.inst\[26\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08300_ net1242 team_03_WB.instance_to_wrap.core.register_file.registers_state\[88\]
+ net972 team_03_WB.instance_to_wrap.core.register_file.registers_state\[120\] net921
+ vssd1 vssd1 vccd1 vccd1 _04242_ sky130_fd_sc_hd__o221a_1
X_09280_ _05217_ _05221_ vssd1 vssd1 vccd1 vccd1 _05222_ sky130_fd_sc_hd__nand2_1
XFILLER_0_129_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08583__A net1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08231_ net1061 _04171_ _04172_ vssd1 vssd1 vccd1 vccd1 _04173_ sky130_fd_sc_hd__or3_1
XFILLER_0_129_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08162_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[532\] net995
+ vssd1 vssd1 vccd1 vccd1 _04104_ sky130_fd_sc_hd__or2_1
XFILLER_0_15_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07113_ net1195 team_03_WB.instance_to_wrap.core.register_file.registers_state\[129\]
+ vssd1 vssd1 vccd1 vccd1 _03055_ sky130_fd_sc_hd__or2_1
XFILLER_0_42_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07803__A1 net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08093_ net1173 team_03_WB.instance_to_wrap.core.register_file.registers_state\[186\]
+ vssd1 vssd1 vccd1 vccd1 _04035_ sky130_fd_sc_hd__and2_1
XFILLER_0_141_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07486__X _03428_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_752 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload50 clknet_leaf_170_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload50/Y sky130_fd_sc_hd__clkinv_2
XANTENNA_clkbuf_4_11__f_wb_clk_i_X clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_07044_ net1118 _02985_ vssd1 vssd1 vccd1 vccd1 _02986_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_77_1950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_1961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload61 clknet_leaf_41_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload61/Y sky130_fd_sc_hd__clkinv_2
Xclkload72 clknet_leaf_52_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload72/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_2_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload83 clknet_leaf_30_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload83/X sky130_fd_sc_hd__clkbuf_8
Xclkload94 clknet_leaf_63_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload94/Y sky130_fd_sc_hd__clkinv_2
XTAP_TAPCELL_ROW_149_3431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_749 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_149_3442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12044__S net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1025_A _06286_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08995_ _04935_ _04936_ net867 vssd1 vssd1 vccd1 vccd1 _04937_ sky130_fd_sc_hd__a21o_1
XFILLER_0_103_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_167_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout485_A _06779_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_10_Left_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09861__B _05686_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07946_ net1088 team_03_WB.instance_to_wrap.core.register_file.registers_state\[887\]
+ net893 vssd1 vssd1 vccd1 vccd1 _03888_ sky130_fd_sc_hd__or3_1
XANTENNA__08758__A net1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_3_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07877_ net751 _03816_ _03818_ net808 vssd1 vssd1 vccd1 vccd1 _03819_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_162_3697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_123_2903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout652_A net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1394_A net1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11184__A net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1135 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09616_ net559 _05357_ vssd1 vssd1 vccd1 vccd1 _05558_ sky130_fd_sc_hd__or2_1
X_06828_ team_03_WB.instance_to_wrap.core.pc.current_pc\[24\] vssd1 vssd1 vccd1 vccd1
+ _02771_ sky130_fd_sc_hd__inv_2
XFILLER_0_92_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09547_ net563 _05486_ _05488_ vssd1 vssd1 vccd1 vccd1 _05489_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout440_X net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout538_X net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout917_A net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11969__A3 net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09478_ net542 _04476_ _05101_ net560 vssd1 vssd1 vccd1 vccd1 _05420_ sky130_fd_sc_hd__a211o_1
XFILLER_0_109_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_484 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08429_ _04369_ _04370_ net1220 vssd1 vssd1 vccd1 vccd1 _04371_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout705_X net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_739 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11440_ net652 _06567_ vssd1 vssd1 vccd1 vccd1 _06760_ sky130_fd_sc_hd__nor2_1
Xclkload0 clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload0/X sky130_fd_sc_hd__clkbuf_8
XANTENNA__09101__B net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_151_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_150_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11371_ net712 net297 net697 vssd1 vssd1 vccd1 vccd1 _06738_ sky130_fd_sc_hd__and3_1
XANTENNA__12743__A net1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10322_ _05968_ _05970_ _06127_ vssd1 vssd1 vccd1 vccd1 _06162_ sky130_fd_sc_hd__or3_1
XANTENNA__09528__S net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13110_ net1258 vssd1 vssd1 vccd1 vccd1 _00874_ sky130_fd_sc_hd__inv_2
X_14090_ clknet_leaf_3_wb_clk_i _01854_ _00455_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[444\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_132_885 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14731__Q team_03_WB.instance_to_wrap.core.decoder.inst\[28\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11359__A net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13041_ net1270 vssd1 vssd1 vccd1 vccd1 _00805_ sky130_fd_sc_hd__inv_2
X_10253_ _04235_ team_03_WB.instance_to_wrap.core.pc.current_pc\[23\] net672 vssd1
+ vssd1 vccd1 vccd1 _06095_ sky130_fd_sc_hd__mux2_1
XANTENNA__11354__A1 net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07558__B1 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11078__B _06434_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07022__A2 net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input46_A gpio_in[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10184_ _03430_ _06025_ vssd1 vssd1 vccd1 vccd1 _06026_ sky130_fd_sc_hd__and2_1
Xfanout1202 net1206 vssd1 vssd1 vccd1 vccd1 net1202 sky130_fd_sc_hd__clkbuf_4
Xfanout1213 team_03_WB.instance_to_wrap.core.decoder.inst\[17\] vssd1 vssd1 vccd1
+ vccd1 net1213 sky130_fd_sc_hd__buf_4
Xfanout1224 net1225 vssd1 vssd1 vccd1 vccd1 net1224 sky130_fd_sc_hd__buf_4
XANTENNA__11793__S net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1235 net1238 vssd1 vssd1 vccd1 vccd1 net1235 sky130_fd_sc_hd__clkbuf_4
Xfanout1246 team_03_WB.instance_to_wrap.core.decoder.inst\[15\] vssd1 vssd1 vccd1
+ vccd1 net1246 sky130_fd_sc_hd__buf_4
XANTENNA__09771__B _04646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14992_ clknet_leaf_66_wb_clk_i net40 _01357_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[11\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1257 net1259 vssd1 vssd1 vccd1 vccd1 net1257 sky130_fd_sc_hd__buf_4
Xclkbuf_leaf_135_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_135_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_31_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout270 _06509_ vssd1 vssd1 vccd1 vccd1 net270 sky130_fd_sc_hd__buf_2
Xfanout1268 net1270 vssd1 vssd1 vccd1 vccd1 net1268 sky130_fd_sc_hd__buf_4
XFILLER_0_79_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout281 _06405_ vssd1 vssd1 vccd1 vccd1 net281 sky130_fd_sc_hd__buf_2
Xfanout1279 net1280 vssd1 vssd1 vccd1 vccd1 net1279 sky130_fd_sc_hd__buf_4
Xfanout292 net293 vssd1 vssd1 vccd1 vccd1 net292 sky130_fd_sc_hd__buf_4
X_13943_ clknet_leaf_78_wb_clk_i _01707_ _00308_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[297\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_159_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13874_ clknet_leaf_164_wb_clk_i _01638_ _00239_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[228\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_159_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07730__B1 net1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_158_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12825_ net1351 vssd1 vssd1 vccd1 vccd1 _00589_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12918__A net1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_1028 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12082__A2 net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12756_ net1305 vssd1 vssd1 vccd1 vccd1 _00520_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_7__f_wb_clk_i_X clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_57_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_155_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11707_ _06749_ net383 net340 net1861 vssd1 vssd1 vccd1 vccd1 _01827_ sky130_fd_sc_hd__a22o_1
XANTENNA__11290__B1 net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12687_ net1337 vssd1 vssd1 vccd1 vccd1 _00451_ sky130_fd_sc_hd__inv_2
XFILLER_0_127_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14426_ clknet_leaf_147_wb_clk_i _02190_ _00791_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[780\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08038__A1 net1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11638_ _06712_ net385 net348 net2523 vssd1 vssd1 vccd1 vccd1 _01894_ sky130_fd_sc_hd__a22o_1
XFILLER_0_86_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_806 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14357_ clknet_leaf_105_wb_clk_i _02121_ _00722_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[711\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11569_ net505 net633 _06677_ net484 net1850 vssd1 vssd1 vccd1 vccd1 _01956_ sky130_fd_sc_hd__a32o_1
XFILLER_0_13_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold707 team_03_WB.instance_to_wrap.core.register_file.registers_state\[923\] vssd1
+ vssd1 vccd1 vccd1 net2200 sky130_fd_sc_hd__dlygate4sd3_1
X_13308_ net1326 vssd1 vssd1 vccd1 vccd1 _01072_ sky130_fd_sc_hd__inv_2
XANTENNA__07747__A net1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold718 team_03_WB.instance_to_wrap.core.register_file.registers_state\[271\] vssd1
+ vssd1 vccd1 vccd1 net2211 sky130_fd_sc_hd__dlygate4sd3_1
Xhold729 team_03_WB.instance_to_wrap.core.register_file.registers_state\[770\] vssd1
+ vssd1 vccd1 vccd1 net2222 sky130_fd_sc_hd__dlygate4sd3_1
X_14288_ clknet_leaf_161_wb_clk_i _02052_ _00653_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[642\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_150_682 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11269__A net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13239_ net1391 vssd1 vssd1 vccd1 vccd1 _01003_ sky130_fd_sc_hd__inv_2
XFILLER_0_21_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08746__C1 net1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_51_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07800_ net1193 team_03_WB.instance_to_wrap.core.register_file.registers_state\[139\]
+ vssd1 vssd1 vccd1 vccd1 _03742_ sky130_fd_sc_hd__or2_1
X_08780_ net1050 team_03_WB.instance_to_wrap.core.register_file.registers_state\[450\]
+ net1002 team_03_WB.instance_to_wrap.core.register_file.registers_state\[482\] net1075
+ vssd1 vssd1 vccd1 vccd1 _04722_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_127_Right_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07731_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[813\] net778
+ net1041 vssd1 vssd1 vccd1 vccd1 _03673_ sky130_fd_sc_hd__o21a_1
X_15085__1471 vssd1 vssd1 vccd1 vccd1 _15085__1471/HI net1471 sky130_fd_sc_hd__conb_1
XANTENNA__11208__S net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_140_3247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09710__B2 net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07662_ net616 _03600_ _03603_ vssd1 vssd1 vccd1 vccd1 _03604_ sky130_fd_sc_hd__a21oi_2
XTAP_TAPCELL_ROW_140_3258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11435__C net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08865__X _04807_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09401_ _05341_ _05342_ vssd1 vssd1 vccd1 vccd1 _05343_ sky130_fd_sc_hd__or2_1
X_07593_ net1203 team_03_WB.instance_to_wrap.core.register_file.registers_state\[89\]
+ net785 team_03_WB.instance_to_wrap.core.register_file.registers_state\[121\] net736
+ vssd1 vssd1 vccd1 vccd1 _03535_ sky130_fd_sc_hd__o221a_1
XFILLER_0_133_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11154__D net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09332_ _05222_ _05236_ _05273_ vssd1 vssd1 vccd1 vccd1 _05274_ sky130_fd_sc_hd__or3b_1
XFILLER_0_62_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08277__A1 net1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08517__S net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_218 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_1118 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09202__A net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09263_ _03727_ _05147_ net608 vssd1 vssd1 vccd1 vccd1 _05205_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_173_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08214_ net1232 team_03_WB.instance_to_wrap.core.register_file.registers_state\[209\]
+ net962 team_03_WB.instance_to_wrap.core.register_file.registers_state\[241\] net936
+ vssd1 vssd1 vccd1 vccd1 _04156_ sky130_fd_sc_hd__o221a_1
XANTENNA__09696__X _05638_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08029__A1 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09226__B1 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09194_ net552 _04712_ _05135_ vssd1 vssd1 vccd1 vccd1 _05136_ sky130_fd_sc_hd__o21ai_1
XANTENNA__11170__C net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_402 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10067__B net1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08145_ _02800_ _02802_ _02811_ _02813_ net1212 vssd1 vssd1 vccd1 vccd1 _04087_ sky130_fd_sc_hd__o221a_1
XFILLER_0_31_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout400_A _06718_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_2751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_116_2762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07788__B1 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_1909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10793__A_N _05799_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08076_ net1186 team_03_WB.instance_to_wrap.core.register_file.registers_state\[854\]
+ vssd1 vssd1 vccd1 vccd1 _04018_ sky130_fd_sc_hd__or2_1
Xclkload150 clknet_leaf_116_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload150/Y sky130_fd_sc_hd__bufinv_16
Xclkload161 clknet_leaf_105_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload161/X sky130_fd_sc_hd__clkbuf_8
Xclkload172 clknet_leaf_88_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload172/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_144_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07027_ net1099 team_03_WB.instance_to_wrap.core.register_file.registers_state\[707\]
+ vssd1 vssd1 vccd1 vccd1 _02969_ sky130_fd_sc_hd__and2_1
XANTENNA__11179__A net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11336__A1 net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1407_A net1408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1028_X net1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_8_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1059 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_164_3737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout390_X net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_164_3748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout488_X net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout867_A net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold12 team_03_WB.instance_to_wrap.core.register_file.registers_state\[991\] vssd1
+ vssd1 vccd1 vccd1 net1505 sky130_fd_sc_hd__dlygate4sd3_1
Xhold23 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1001\] vssd1
+ vssd1 vccd1 vccd1 net1516 sky130_fd_sc_hd__dlygate4sd3_1
Xhold34 _02615_ vssd1 vssd1 vccd1 vccd1 net1527 sky130_fd_sc_hd__dlygate4sd3_1
X_08978_ _04916_ _04917_ _04919_ _04918_ net945 net865 vssd1 vssd1 vccd1 vccd1 _04920_
+ sky130_fd_sc_hd__mux4_1
Xhold45 team_03_WB.instance_to_wrap.core.register_file.registers_state\[957\] vssd1
+ vssd1 vccd1 vccd1 net1538 sky130_fd_sc_hd__dlygate4sd3_1
Xhold56 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1013\] vssd1
+ vssd1 vccd1 vccd1 net1549 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07392__A net1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold67 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[6\] vssd1 vssd1 vccd1
+ vccd1 net1560 sky130_fd_sc_hd__dlygate4sd3_1
Xhold78 team_03_WB.instance_to_wrap.core.register_file.registers_state\[946\] vssd1
+ vssd1 vccd1 vccd1 net1571 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11639__A2 net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07929_ net743 _03867_ _03868_ _03869_ _03870_ vssd1 vssd1 vccd1 vccd1 _03871_ sky130_fd_sc_hd__o32a_1
Xhold89 team_03_WB.instance_to_wrap.core.register_file.registers_state\[997\] vssd1
+ vssd1 vccd1 vccd1 net1582 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout655_X net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09701__A1 _02954_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10847__A0 net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10940_ team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[6\] net307 net689 vssd1
+ vssd1 vccd1 vccd1 _06525_ sky130_fd_sc_hd__a21o_1
XANTENNA__11345__C net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07712__B1 net1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11064__D _06463_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10871_ net833 _06468_ vssd1 vssd1 vccd1 vccd1 _06469_ sky130_fd_sc_hd__and2_2
XANTENNA_fanout822_X net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_1106 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input100_A wbs_dat_i[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12610_ net1350 vssd1 vssd1 vccd1 vccd1 _00374_ sky130_fd_sc_hd__inv_2
XFILLER_0_66_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_842 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13590_ net1344 vssd1 vssd1 vccd1 vccd1 _01354_ sky130_fd_sc_hd__inv_2
XFILLER_0_149_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14726__Q team_03_WB.instance_to_wrap.core.decoder.inst\[23\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11361__B net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07476__C1 net1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12541_ net1383 vssd1 vssd1 vccd1 vccd1 _00305_ sky130_fd_sc_hd__inv_2
XANTENNA__11272__B1 net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11811__A2 net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09217__B1 _02937_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12472_ net1380 vssd1 vssd1 vccd1 vccd1 _00236_ sky130_fd_sc_hd__inv_2
XFILLER_0_35_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14211_ clknet_leaf_32_wb_clk_i _01975_ _00576_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[565\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11788__S net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11423_ net296 net2457 net399 vssd1 vssd1 vccd1 vccd1 _02059_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11354_ net502 net629 _06729_ net401 net2138 vssd1 vssd1 vccd1 vccd1 _02103_ sky130_fd_sc_hd__a32o_1
XFILLER_0_22_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14142_ clknet_leaf_120_wb_clk_i _01906_ _00507_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[496\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07567__A net1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08440__A1 net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10305_ team_03_WB.instance_to_wrap.core.pc.current_pc\[22\] _06146_ vssd1 vssd1
+ vccd1 vccd1 _06147_ sky130_fd_sc_hd__and2_1
XFILLER_0_131_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14073_ clknet_leaf_169_wb_clk_i _01837_ _00438_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[427\]
+ sky130_fd_sc_hd__dfrtp_1
X_11285_ net712 _06527_ net831 vssd1 vssd1 vccd1 vccd1 _06710_ sky130_fd_sc_hd__and3_1
XFILLER_0_67_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10236_ net588 _02773_ net674 vssd1 vssd1 vccd1 vccd1 _06078_ sky130_fd_sc_hd__mux2_1
X_13024_ net1403 vssd1 vssd1 vccd1 vccd1 _00788_ sky130_fd_sc_hd__inv_2
Xfanout1010 net1012 vssd1 vssd1 vccd1 vccd1 net1010 sky130_fd_sc_hd__buf_2
XANTENNA__11239__D net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1021 net1022 vssd1 vssd1 vccd1 vccd1 net1021 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout1032 net1033 vssd1 vssd1 vccd1 vccd1 net1032 sky130_fd_sc_hd__clkbuf_4
X_10167_ _06008_ vssd1 vssd1 vccd1 vccd1 _06009_ sky130_fd_sc_hd__inv_2
Xfanout1043 net1044 vssd1 vssd1 vccd1 vccd1 net1043 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_174_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1054 net1055 vssd1 vssd1 vccd1 vccd1 net1054 sky130_fd_sc_hd__clkbuf_2
Xfanout1065 net1066 vssd1 vssd1 vccd1 vccd1 net1065 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_156_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1076 net1080 vssd1 vssd1 vccd1 vccd1 net1076 sky130_fd_sc_hd__buf_4
X_14975_ clknet_leaf_85_wb_clk_i _02727_ _01340_ vssd1 vssd1 vccd1 vccd1 net227 sky130_fd_sc_hd__dfrtp_1
X_10098_ _02924_ _02935_ _02936_ _05917_ vssd1 vssd1 vccd1 vccd1 _05942_ sky130_fd_sc_hd__a211o_1
Xfanout1087 net1088 vssd1 vssd1 vccd1 vccd1 net1087 sky130_fd_sc_hd__buf_2
Xfanout1098 net1101 vssd1 vssd1 vccd1 vccd1 net1098 sky130_fd_sc_hd__buf_2
X_13926_ clknet_leaf_28_wb_clk_i _01690_ _00291_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[280\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11255__C net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_55 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07703__B1 net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08900__C1 net1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13857_ clknet_leaf_179_wb_clk_i _01621_ _00222_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[211\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11552__A net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12808_ net1293 vssd1 vssd1 vccd1 vccd1 _00572_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_48_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13788_ clknet_leaf_149_wb_clk_i _01552_ _00153_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[142\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07467__C1 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11271__B net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_32_wb_clk_i clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_32_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_12739_ net1374 vssd1 vssd1 vccd1 vccd1 _00503_ sky130_fd_sc_hd__inv_2
XFILLER_0_84_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_2009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_44_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_167_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_96_2345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07219__C1 net1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_2356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14409_ clknet_leaf_74_wb_clk_i _02173_ _00774_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[763\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_4_346 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11566__A1 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08967__C1 net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold504 team_03_WB.instance_to_wrap.CPU_DAT_I\[25\] vssd1 vssd1 vccd1 vccd1 net1997
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold515 team_03_WB.instance_to_wrap.core.register_file.registers_state\[364\] vssd1
+ vssd1 vccd1 vccd1 net2008 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07865__S0 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold526 team_03_WB.instance_to_wrap.core.register_file.registers_state\[421\] vssd1
+ vssd1 vccd1 vccd1 net2019 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold537 team_03_WB.instance_to_wrap.core.register_file.registers_state\[227\] vssd1
+ vssd1 vccd1 vccd1 net2030 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold548 team_03_WB.instance_to_wrap.core.register_file.registers_state\[690\] vssd1
+ vssd1 vccd1 vccd1 net2041 sky130_fd_sc_hd__dlygate4sd3_1
Xhold559 team_03_WB.instance_to_wrap.core.register_file.registers_state\[163\] vssd1
+ vssd1 vccd1 vccd1 net2052 sky130_fd_sc_hd__dlygate4sd3_1
X_09950_ _05879_ net1707 net291 vssd1 vssd1 vccd1 vccd1 _02752_ sky130_fd_sc_hd__mux2_1
XANTENNA__09963__Y _05886_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08901_ net1239 team_03_WB.instance_to_wrap.core.register_file.registers_state\[460\]
+ net979 team_03_WB.instance_to_wrap.core.register_file.registers_state\[492\] net1215
+ vssd1 vssd1 vccd1 vccd1 _04843_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_70_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09881_ _05803_ _05811_ _05821_ _05646_ vssd1 vssd1 vccd1 vccd1 _05823_ sky130_fd_sc_hd__or4b_1
XTAP_TAPCELL_ROW_70_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08195__B1 net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08832_ net557 _04713_ _04773_ net572 vssd1 vssd1 vccd1 vccd1 _04774_ sky130_fd_sc_hd__o211a_1
Xhold1204 team_03_WB.instance_to_wrap.core.register_file.registers_state\[846\] vssd1
+ vssd1 vccd1 vccd1 net2697 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10541__A2 net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1215 team_03_WB.instance_to_wrap.core.register_file.registers_state\[136\] vssd1
+ vssd1 vccd1 vccd1 net2708 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07942__B1 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1226 team_03_WB.instance_to_wrap.core.register_file.registers_state\[219\] vssd1
+ vssd1 vccd1 vccd1 net2719 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1237 team_03_WB.instance_to_wrap.core.register_file.registers_state\[91\] vssd1
+ vssd1 vccd1 vccd1 net2730 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11446__B net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08763_ net1221 _04704_ vssd1 vssd1 vccd1 vccd1 _04705_ sky130_fd_sc_hd__or2_1
Xhold1248 team_03_WB.instance_to_wrap.core.register_file.registers_state\[710\] vssd1
+ vssd1 vccd1 vccd1 net2741 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1259 team_03_WB.instance_to_wrap.core.register_file.registers_state\[471\] vssd1
+ vssd1 vccd1 vccd1 net2752 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07714_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[397\] net800
+ _02869_ _03655_ vssd1 vssd1 vccd1 vccd1 _03656_ sky130_fd_sc_hd__o211a_1
XFILLER_0_79_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08694_ net1241 team_03_WB.instance_to_wrap.core.register_file.registers_state\[72\]
+ net957 team_03_WB.instance_to_wrap.core.register_file.registers_state\[104\] net918
+ vssd1 vssd1 vccd1 vccd1 _04636_ sky130_fd_sc_hd__o221a_1
XFILLER_0_79_135 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07645_ net1094 team_03_WB.instance_to_wrap.core.register_file.registers_state\[718\]
+ net798 team_03_WB.instance_to_wrap.core.register_file.registers_state\[750\] vssd1
+ vssd1 vccd1 vccd1 _03587_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_68_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1092_A net1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout448_A _06801_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07576_ net1092 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1016\]
+ net894 _03517_ net1153 vssd1 vssd1 vccd1 vccd1 _03518_ sky130_fd_sc_hd__o311a_1
XFILLER_0_165_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10057__A1 net30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09315_ _02938_ _05124_ vssd1 vssd1 vccd1 vccd1 _05257_ sky130_fd_sc_hd__nor2_1
XANTENNA__11181__B net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11254__B1 net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10078__A _02937_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_823 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout615_A net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_157_3596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_2802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1357_A net1358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_663 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09246_ _03391_ _05152_ net607 vssd1 vssd1 vccd1 vccd1 _05188_ sky130_fd_sc_hd__a21o_1
XFILLER_0_161_711 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09586__B _04382_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09177_ net546 net350 _05118_ vssd1 vssd1 vccd1 vccd1 _05119_ sky130_fd_sc_hd__o21ba_1
XANTENNA_fanout403_X net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11401__S net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_934 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08128_ team_03_WB.instance_to_wrap.core.decoder.inst\[26\] net1019 net684 vssd1
+ vssd1 vccd1 vccd1 _04070_ sky130_fd_sc_hd__a21oi_2
XANTENNA__08958__C1 net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08422__A1 net1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07818__C net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_160_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout984_A net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08059_ net1186 team_03_WB.instance_to_wrap.core.register_file.registers_state\[342\]
+ vssd1 vssd1 vccd1 vccd1 _04001_ sky130_fd_sc_hd__or2_1
X_11070_ net832 net279 vssd1 vssd1 vccd1 vccd1 _06613_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout772_X net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11059__D net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput102 wbs_we_i vssd1 vssd1 vccd1 vccd1 net102 sky130_fd_sc_hd__clkbuf_1
X_10021_ net77 net76 _05897_ _05898_ vssd1 vssd1 vccd1 vccd1 _05899_ sky130_fd_sc_hd__or4_1
XANTENNA__10532__A2 net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07933__B1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14760_ clknet_leaf_49_wb_clk_i net1682 _01125_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09686__B1 _03985_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11972_ net636 _06749_ net469 net365 net2261 vssd1 vssd1 vccd1 vccd1 _01571_ sky130_fd_sc_hd__a32o_1
XANTENNA__07850__A net1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13711_ clknet_leaf_136_wb_clk_i _01475_ _00076_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[65\]
+ sky130_fd_sc_hd__dfrtp_1
X_10923_ net313 net309 net316 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[9\]
+ vssd1 vssd1 vccd1 vccd1 _06511_ sky130_fd_sc_hd__o31a_1
XFILLER_0_168_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14691_ clknet_leaf_57_wb_clk_i _02455_ _01056_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.ADR_I\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10835__A3 net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_19_Right_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13642_ net1406 vssd1 vssd1 vccd1 vccd1 _01406_ sky130_fd_sc_hd__inv_2
X_10854_ _06450_ _06451_ _06452_ vssd1 vssd1 vccd1 vccd1 _06453_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_128_207 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10048__A1 net8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11091__B net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13573_ net1406 vssd1 vssd1 vccd1 vccd1 _01337_ sky130_fd_sc_hd__inv_2
XFILLER_0_94_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10785_ _06381_ _06382_ _06394_ vssd1 vssd1 vccd1 vccd1 _06395_ sky130_fd_sc_hd__or3b_4
XANTENNA__11522__D net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12524_ net1333 vssd1 vssd1 vccd1 vccd1 _00288_ sky130_fd_sc_hd__inv_2
XFILLER_0_82_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_435 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15084__1470 vssd1 vssd1 vccd1 vccd1 _15084__1470/HI net1470 sky130_fd_sc_hd__conb_1
XFILLER_0_48_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12455_ net1369 vssd1 vssd1 vccd1 vccd1 _00219_ sky130_fd_sc_hd__inv_2
XANTENNA__11311__S net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_934 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11548__B2 net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11406_ net276 net2621 net399 vssd1 vssd1 vccd1 vccd1 _02074_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_10_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12386_ net1360 vssd1 vssd1 vccd1 vccd1 _00150_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_28_Right_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10220__A1 _06057_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14125_ clknet_leaf_188_wb_clk_i _01889_ _00490_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[479\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_2242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11337_ net1250 net837 _06413_ net668 vssd1 vssd1 vccd1 vccd1 _06721_ sky130_fd_sc_hd__and4_1
XFILLER_0_120_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_150_wb_clk_i clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_150_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_91_2253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07584__X _03526_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14056_ clknet_leaf_18_wb_clk_i _01820_ _00421_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[410\]
+ sky130_fd_sc_hd__dfrtp_1
X_11268_ net501 net630 _06701_ net409 net1994 vssd1 vssd1 vccd1 vccd1 _02161_ sky130_fd_sc_hd__a32o_1
XANTENNA__11547__A net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13007_ net1336 vssd1 vssd1 vccd1 vccd1 _00771_ sky130_fd_sc_hd__inv_2
X_10219_ _06024_ _06060_ vssd1 vssd1 vccd1 vccd1 _06061_ sky130_fd_sc_hd__nor2_1
X_11199_ net281 net2434 net486 vssd1 vssd1 vccd1 vccd1 _02209_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_49 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10523__A2 net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11720__A1 net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09017__A net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11981__S net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_168_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14958_ clknet_leaf_94_wb_clk_i _02710_ _01323_ vssd1 vssd1 vccd1 vccd1 net210 sky130_fd_sc_hd__dfrtp_1
XANTENNA__09677__B1 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_37_Right_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07760__A net1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07688__C1 net1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13909_ clknet_leaf_126_wb_clk_i _01673_ _00274_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[263\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_159_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14889_ clknet_leaf_58_wb_clk_i _02652_ _01254_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.pc.current_pc\[18\]
+ sky130_fd_sc_hd__dfrtp_2
X_07430_ net1138 _03367_ _03369_ _03371_ net721 vssd1 vssd1 vccd1 vccd1 _03372_ sky130_fd_sc_hd__o41a_1
XTAP_TAPCELL_ROW_46_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12028__A2 net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10039__A1 net18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10039__B2 team_03_WB.instance_to_wrap.CPU_DAT_O\[24\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_730 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11236__B1 net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07361_ net821 _03290_ net717 vssd1 vssd1 vccd1 vccd1 _03303_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_31_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08101__B1 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09100_ net436 net428 _05041_ net550 vssd1 vssd1 vccd1 vccd1 _05042_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_21_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07292_ net1202 team_03_WB.instance_to_wrap.core.register_file.registers_state\[329\]
+ net783 team_03_WB.instance_to_wrap.core.register_file.registers_state\[361\] net1136
+ vssd1 vssd1 vccd1 vccd1 _03234_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_135_3146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_3157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10087__B_N _05697_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09031_ _04971_ _04972_ net865 vssd1 vssd1 vccd1 vccd1 _04973_ sky130_fd_sc_hd__o21a_1
XFILLER_0_150_87 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_46_Right_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11539__B2 net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_152_3493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08404__A1 net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_276 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold301 team_03_WB.instance_to_wrap.core.register_file.registers_state\[313\] vssd1
+ vssd1 vccd1 vccd1 net1794 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07838__S0 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_27_wb_clk_i_A clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold312 team_03_WB.instance_to_wrap.core.register_file.registers_state\[317\] vssd1
+ vssd1 vccd1 vccd1 net1805 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07000__A team_03_WB.instance_to_wrap.core.decoder.inst\[14\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold323 team_03_WB.instance_to_wrap.core.register_file.registers_state\[828\] vssd1
+ vssd1 vccd1 vccd1 net1816 sky130_fd_sc_hd__dlygate4sd3_1
Xhold334 team_03_WB.instance_to_wrap.core.register_file.registers_state\[692\] vssd1
+ vssd1 vccd1 vccd1 net1827 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07612__C1 net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold345 _02597_ vssd1 vssd1 vccd1 vccd1 net1838 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10913__X _06503_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12841__A net1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold356 team_03_WB.instance_to_wrap.CPU_DAT_O\[15\] vssd1 vssd1 vccd1 vccd1 net1849
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06966__A1 net1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_850 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_1132 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10064__C net1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold367 team_03_WB.instance_to_wrap.core.register_file.registers_state\[439\] vssd1
+ vssd1 vccd1 vccd1 net1860 sky130_fd_sc_hd__dlygate4sd3_1
Xhold378 team_03_WB.instance_to_wrap.core.register_file.registers_state\[434\] vssd1
+ vssd1 vccd1 vccd1 net1871 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09933_ _03821_ net662 vssd1 vssd1 vccd1 vccd1 _05871_ sky130_fd_sc_hd__nor2_1
Xhold389 team_03_WB.instance_to_wrap.core.register_file.registers_state\[293\] vssd1
+ vssd1 vccd1 vccd1 net1882 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout803 net804 vssd1 vssd1 vccd1 vccd1 net803 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_1_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout814 net816 vssd1 vssd1 vccd1 vccd1 net814 sky130_fd_sc_hd__clkbuf_4
Xfanout825 _02846_ vssd1 vssd1 vccd1 vccd1 net825 sky130_fd_sc_hd__buf_4
XFILLER_0_99_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10999__C net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout398_A _06752_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout836 net837 vssd1 vssd1 vccd1 vccd1 net836 sky130_fd_sc_hd__buf_2
Xfanout847 _06303_ vssd1 vssd1 vccd1 vccd1 net847 sky130_fd_sc_hd__buf_2
X_09864_ _03947_ net590 _05805_ _02945_ vssd1 vssd1 vccd1 vccd1 _05806_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__12052__S net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout858 _04084_ vssd1 vssd1 vccd1 vccd1 net858 sky130_fd_sc_hd__buf_8
XANTENNA__10514__A2 net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout869 net870 vssd1 vssd1 vccd1 vccd1 net869 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11711__A1 net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1105_A _02787_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07915__B1 net1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1001 team_03_WB.instance_to_wrap.core.register_file.registers_state\[400\] vssd1
+ vssd1 vccd1 vccd1 net2494 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1012 team_03_WB.instance_to_wrap.core.register_file.registers_state\[783\] vssd1
+ vssd1 vccd1 vccd1 net2505 sky130_fd_sc_hd__dlygate4sd3_1
X_08815_ net1052 team_03_WB.instance_to_wrap.core.register_file.registers_state\[961\]
+ net1004 team_03_WB.instance_to_wrap.core.register_file.registers_state\[993\] net1065
+ vssd1 vssd1 vccd1 vccd1 _04757_ sky130_fd_sc_hd__a221o_1
XFILLER_0_99_208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1023 team_03_WB.instance_to_wrap.core.register_file.registers_state\[134\] vssd1
+ vssd1 vccd1 vccd1 net2516 sky130_fd_sc_hd__dlygate4sd3_1
X_09795_ net578 _05736_ vssd1 vssd1 vccd1 vccd1 _05737_ sky130_fd_sc_hd__or2_1
Xhold1034 team_03_WB.instance_to_wrap.core.register_file.registers_state\[324\] vssd1
+ vssd1 vccd1 vccd1 net2527 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout565_A _03025_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07391__A1 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1045 team_03_WB.instance_to_wrap.core.register_file.registers_state\[577\] vssd1
+ vssd1 vccd1 vccd1 net2538 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_55_Right_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1056 team_03_WB.instance_to_wrap.core.register_file.registers_state\[833\] vssd1
+ vssd1 vccd1 vccd1 net2549 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1067 team_03_WB.instance_to_wrap.core.register_file.registers_state\[615\] vssd1
+ vssd1 vccd1 vccd1 net2560 sky130_fd_sc_hd__dlygate4sd3_1
X_08746_ net1052 team_03_WB.instance_to_wrap.core.register_file.registers_state\[323\]
+ net1005 team_03_WB.instance_to_wrap.core.register_file.registers_state\[355\] net1214
+ vssd1 vssd1 vccd1 vccd1 _04688_ sky130_fd_sc_hd__a221o_1
Xhold1078 team_03_WB.instance_to_wrap.core.register_file.registers_state\[229\] vssd1
+ vssd1 vccd1 vccd1 net2571 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_107_2569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1089 team_03_WB.instance_to_wrap.core.register_file.registers_state\[212\] vssd1
+ vssd1 vccd1 vccd1 net2582 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07670__A net1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12288__A net1402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout732_A net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07143__A1 net1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08677_ _04607_ _04618_ net853 vssd1 vssd1 vccd1 vccd1 _04619_ sky130_fd_sc_hd__mux2_4
XTAP_TAPCELL_ROW_159_3636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11192__A net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_159_3647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07628_ net1094 team_03_WB.instance_to_wrap.core.register_file.registers_state\[174\]
+ net896 vssd1 vssd1 vccd1 vccd1 _03570_ sky130_fd_sc_hd__or3_1
XFILLER_0_36_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07694__A2 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11227__A0 _06527_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout520_X net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07559_ net1188 team_03_WB.instance_to_wrap.core.register_file.registers_state\[344\]
+ net771 team_03_WB.instance_to_wrap.core.register_file.registers_state\[376\] vssd1
+ vssd1 vccd1 vccd1 _03501_ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout618_X net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_66_wb_clk_i_A clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_10570_ net1779 net531 net598 _05880_ vssd1 vssd1 vccd1 vccd1 _02553_ sky130_fd_sc_hd__a22o_1
XFILLER_0_9_983 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08643__A1 net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_64_Right_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10450__A1 team_03_WB.instance_to_wrap.core.pc.current_pc\[4\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09229_ _05170_ vssd1 vssd1 vccd1 vccd1 _05171_ sky130_fd_sc_hd__inv_2
XFILLER_0_133_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07851__C1 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_1043 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12240_ net1616 vssd1 vssd1 vccd1 vccd1 _01417_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__08006__A net1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout987_X net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12171_ net1636 vssd1 vssd1 vccd1 vccd1 _02382_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_2_Left_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11950__A1 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11122_ net281 net646 net703 net695 vssd1 vssd1 vccd1 vccd1 _06636_ sky130_fd_sc_hd__and4_1
Xhold890 team_03_WB.instance_to_wrap.core.register_file.registers_state\[495\] vssd1
+ vssd1 vccd1 vccd1 net2383 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11367__A net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11053_ net1043 net838 _06536_ net671 vssd1 vssd1 vccd1 vccd1 _06604_ sky130_fd_sc_hd__and4_1
XANTENNA__07057__S1 net1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07906__B1 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10004_ _05889_ net1733 net288 vssd1 vssd1 vccd1 vccd1 _02710_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_73_Right_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07283__C net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07382__A1 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09108__C1 net1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14812_ clknet_leaf_92_wb_clk_i net1645 _01177_ vssd1 vssd1 vccd1 vccd1 net163 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_118_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_1134 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07580__A net1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14743_ clknet_leaf_68_wb_clk_i _02507_ _01108_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_11955_ net618 _06732_ net451 net363 net2147 vssd1 vssd1 vccd1 vccd1 _01588_ sky130_fd_sc_hd__a32o_1
XFILLER_0_99_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_28_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06908__B net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_116 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11306__S net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10906_ net313 net309 net316 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[12\]
+ vssd1 vssd1 vccd1 vccd1 _06497_ sky130_fd_sc_hd__o31a_1
X_14674_ clknet_leaf_81_wb_clk_i _02438_ _01039_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.ADR_I\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_156_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11886_ net627 _06695_ net458 net372 net2021 vssd1 vssd1 vccd1 vccd1 _01655_ sky130_fd_sc_hd__a32o_1
XANTENNA__11218__A0 _06495_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_168_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13625_ net1430 vssd1 vssd1 vccd1 vccd1 _01389_ sky130_fd_sc_hd__inv_2
XFILLER_0_27_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10837_ net301 net2308 net519 vssd1 vssd1 vccd1 vccd1 _02329_ sky130_fd_sc_hd__mux2_1
XFILLER_0_144_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_82_Right_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_15_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_379 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13556_ net1416 vssd1 vssd1 vccd1 vccd1 _01320_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_41_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10768_ _05142_ net605 vssd1 vssd1 vccd1 vccd1 _06379_ sky130_fd_sc_hd__nand2_1
XANTENNA__09831__B1 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14914__Q team_03_WB.instance_to_wrap.CPU_DAT_O\[1\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_12507_ net1361 vssd1 vssd1 vccd1 vccd1 _00271_ sky130_fd_sc_hd__inv_2
XANTENNA__07842__C1 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13487_ net1343 vssd1 vssd1 vccd1 vccd1 _01251_ sky130_fd_sc_hd__inv_2
X_10699_ _05455_ _06310_ vssd1 vssd1 vccd1 vccd1 _06337_ sky130_fd_sc_hd__nor2_1
XANTENNA__09794__X _05736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12438_ net1280 vssd1 vssd1 vccd1 vccd1 _00202_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_130_3043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_3054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11976__S net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12369_ net1266 vssd1 vssd1 vccd1 vccd1 _00133_ sky130_fd_sc_hd__inv_2
X_14108_ clknet_leaf_147_wb_clk_i _01872_ _00473_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[462\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07070__B1 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15088_ net1474 vssd1 vssd1 vccd1 vccd1 la_data_out[24] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_39_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_91_Right_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11277__A net1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06930_ net1153 net1163 vssd1 vssd1 vccd1 vccd1 _02872_ sky130_fd_sc_hd__or2_4
X_14039_ clknet_leaf_116_wb_clk_i _01803_ _00404_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[393\]
+ sky130_fd_sc_hd__dfrtp_1
X_06861_ _02800_ _02802_ vssd1 vssd1 vccd1 vccd1 _02803_ sky130_fd_sc_hd__nor2_1
XANTENNA__08796__S1 net1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07373__A1 net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08600_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[549\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[517\]
+ net993 vssd1 vssd1 vccd1 vccd1 _04542_ sky130_fd_sc_hd__mux2_1
XANTENNA__07912__A3 net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09580_ _05396_ _05402_ net565 vssd1 vssd1 vccd1 vccd1 _05522_ sky130_fd_sc_hd__mux2_1
XFILLER_0_145_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08531_ net1218 _04471_ _04472_ vssd1 vssd1 vccd1 vccd1 _04473_ sky130_fd_sc_hd__o21ai_1
XANTENNA__11457__B1 net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_100_wb_clk_i_A clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08322__B1 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11216__S net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08462_ net933 _04402_ _04403_ vssd1 vssd1 vccd1 vccd1 _04404_ sky130_fd_sc_hd__o21a_1
XFILLER_0_161_31 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11209__A0 net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_102_2466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07413_ net1175 team_03_WB.instance_to_wrap.core.register_file.registers_state\[724\]
+ net763 team_03_WB.instance_to_wrap.core.register_file.registers_state\[756\] net741
+ vssd1 vssd1 vccd1 vccd1 _03355_ sky130_fd_sc_hd__o221a_1
X_08393_ net1245 team_03_WB.instance_to_wrap.core.register_file.registers_state\[345\]
+ net991 team_03_WB.instance_to_wrap.core.register_file.registers_state\[377\] net1078
+ vssd1 vssd1 vccd1 vccd1 _04335_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_102_2477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10908__X _06499_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_845 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_154_3533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07344_ net1170 team_03_WB.instance_to_wrap.core.register_file.registers_state\[92\]
+ net759 team_03_WB.instance_to_wrap.core.register_file.registers_state\[124\] net725
+ vssd1 vssd1 vccd1 vccd1 _03286_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_154_3544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_169_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09210__A net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07275_ net1140 _03216_ net724 vssd1 vssd1 vccd1 vccd1 _03217_ sky130_fd_sc_hd__o21a_1
XANTENNA__12047__S net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_171_3880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout313_A _05387_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_171_3891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_872 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1055_A net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09014_ _04923_ _04955_ vssd1 vssd1 vccd1 vccd1 _04956_ sky130_fd_sc_hd__nor2_1
XFILLER_0_5_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_170_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08389__B1 net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold120 _02611_ vssd1 vssd1 vccd1 vccd1 net1613 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold131 team_03_WB.instance_to_wrap.core.ru.state\[2\] vssd1 vssd1 vccd1 vccd1 net1624
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09050__A1 net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold142 team_03_WB.instance_to_wrap.core.register_file.registers_state\[974\] vssd1
+ vssd1 vccd1 vccd1 net1635 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1222_A net1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10735__A2 net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold153 team_03_WB.instance_to_wrap.core.register_file.registers_state\[951\] vssd1
+ vssd1 vccd1 vccd1 net1646 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07061__B1 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold164 _02590_ vssd1 vssd1 vccd1 vccd1 net1657 sky130_fd_sc_hd__dlygate4sd3_1
Xhold175 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[13\] vssd1 vssd1 vccd1
+ vccd1 net1668 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout682_A _05915_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold186 team_03_WB.instance_to_wrap.ADR_I\[3\] vssd1 vssd1 vccd1 vccd1 net1679 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout600 _06299_ vssd1 vssd1 vccd1 vccd1 net600 sky130_fd_sc_hd__clkbuf_2
Xhold197 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1006\] vssd1
+ vssd1 vccd1 vccd1 net1690 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout611 net612 vssd1 vssd1 vccd1 vccd1 net611 sky130_fd_sc_hd__buf_2
X_09916_ _02837_ _05142_ _05799_ _05857_ vssd1 vssd1 vccd1 vccd1 _05858_ sky130_fd_sc_hd__or4b_1
XFILLER_0_10_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout622 net625 vssd1 vssd1 vccd1 vccd1 net622 sky130_fd_sc_hd__clkbuf_4
Xfanout633 net634 vssd1 vssd1 vccd1 vccd1 net633 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout1010_X net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout644 net645 vssd1 vssd1 vccd1 vccd1 net644 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_109_2609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1108_X net1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout655 net659 vssd1 vssd1 vccd1 vccd1 net655 sky130_fd_sc_hd__buf_4
XANTENNA__09880__A _05821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout666 net667 vssd1 vssd1 vccd1 vccd1 net666 sky130_fd_sc_hd__clkbuf_2
Xfanout677 net678 vssd1 vssd1 vccd1 vccd1 net677 sky130_fd_sc_hd__buf_2
X_09847_ net570 net592 net667 _05788_ vssd1 vssd1 vccd1 vccd1 _05789_ sky130_fd_sc_hd__a22o_1
XANTENNA__11696__B1 net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout688 net690 vssd1 vssd1 vccd1 vccd1 net688 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout470_X net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout947_A net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07364__A1 net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout699 net700 vssd1 vssd1 vccd1 vccd1 net699 sky130_fd_sc_hd__buf_4
XANTENNA__11337__D net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09778_ _05270_ _05719_ vssd1 vssd1 vccd1 vccd1 _05720_ sky130_fd_sc_hd__xnor2_2
XTAP_TAPCELL_ROW_126_2967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08729_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[932\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[900\]
+ net977 vssd1 vssd1 vccd1 vccd1 _04671_ sky130_fd_sc_hd__mux2_1
XANTENNA__07116__A1 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout735_X net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_803 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09879__X _05821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11740_ net597 _06546_ net466 _06808_ net1870 vssd1 vssd1 vccd1 vccd1 _01796_ sky130_fd_sc_hd__a32o_1
XANTENNA__11353__C _06561_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08864__A1 net1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_189_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout902_X net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11671_ net2265 net264 net344 vssd1 vssd1 vccd1 vccd1 _01862_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_666 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13410_ net1415 vssd1 vssd1 vccd1 vccd1 _01174_ sky130_fd_sc_hd__inv_2
X_10622_ net2328 team_03_WB.instance_to_wrap.CPU_DAT_O\[7\] net842 vssd1 vssd1 vccd1
+ vccd1 _02506_ sky130_fd_sc_hd__mux2_1
XANTENNA__08077__C1 net1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08616__A1 net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14390_ clknet_leaf_152_wb_clk_i _02154_ _00755_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[744\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_12_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08435__S net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09813__B1 _05650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14734__Q team_03_WB.instance_to_wrap.core.decoder.inst\[31\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13341_ net1334 vssd1 vssd1 vccd1 vccd1 _01105_ sky130_fd_sc_hd__inv_2
XFILLER_0_84_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11620__B1 net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10553_ net1145 team_03_WB.instance_to_wrap.core.ru.state\[5\] vssd1 vssd1 vccd1
+ vccd1 _06296_ sky130_fd_sc_hd__nor2_1
XFILLER_0_148_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07824__C1 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10266__A _03528_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08092__A2 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_703 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1069 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10974__A2 _05845_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_347 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13272_ net1423 vssd1 vssd1 vccd1 vccd1 _01036_ sky130_fd_sc_hd__inv_2
XANTENNA_input76_A wbs_adr_i[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10484_ net1691 net1028 net905 net1676 vssd1 vssd1 vccd1 vccd1 _02625_ sky130_fd_sc_hd__a22o_1
XFILLER_0_121_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_161_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11796__S net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15011_ clknet_leaf_40_wb_clk_i net59 _01376_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[30\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__13577__A net1435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12223_ net1610 vssd1 vssd1 vccd1 vccd1 _01434_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__10187__A0 _04591_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09041__A1 net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12481__A net1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07575__A net1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12154_ net1675 vssd1 vssd1 vccd1 vccd1 _02399_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__08170__S net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11105_ _06628_ net2023 net419 vssd1 vssd1 vccd1 vccd1 _02251_ sky130_fd_sc_hd__mux2_1
XANTENNA__11097__A net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12085_ net624 _06651_ net455 net439 net1737 vssd1 vssd1 vccd1 vccd1 _01462_ sky130_fd_sc_hd__a32o_1
XFILLER_0_120_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11687__B1 net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11036_ net633 _06593_ vssd1 vssd1 vccd1 vccd1 _06594_ sky130_fd_sc_hd__nor2_1
XFILLER_0_21_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_34_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07355__A1 net1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11151__A2 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08552__B1 net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06919__A net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12987_ net1361 vssd1 vssd1 vccd1 vccd1 _00751_ sky130_fd_sc_hd__inv_2
XFILLER_0_115_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12100__A1 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08304__B1 net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14726_ clknet_leaf_53_wb_clk_i _02490_ _01091_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.decoder.inst\[23\]
+ sky130_fd_sc_hd__dfrtp_4
X_11938_ net263 net2528 net369 vssd1 vssd1 vccd1 vccd1 _01604_ sky130_fd_sc_hd__mux2_1
XANTENNA__11263__C _06477_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_157_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14657_ clknet_leaf_179_wb_clk_i _02421_ _01022_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1011\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_46_119 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09949__B net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11869_ net269 net2082 net378 vssd1 vssd1 vccd1 vccd1 _01671_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_60_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06961__S0 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13608_ net1320 vssd1 vssd1 vccd1 vccd1 _01372_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08068__C1 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14588_ clknet_leaf_151_wb_clk_i _02352_ _00953_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[942\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_54_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10414__B2 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13539_ net1326 vssd1 vssd1 vccd1 vccd1 _01303_ sky130_fd_sc_hd__inv_2
XANTENNA__11611__B1 net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_528 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07060_ net1097 team_03_WB.instance_to_wrap.core.register_file.registers_state\[578\]
+ net797 team_03_WB.instance_to_wrap.core.register_file.registers_state\[610\] net746
+ vssd1 vssd1 vccd1 vccd1 _03002_ sky130_fd_sc_hd__a221o_1
XFILLER_0_153_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09965__A _03756_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07291__B1 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_140_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput203 net203 vssd1 vssd1 vccd1 vccd1 gpio_oeb[7] sky130_fd_sc_hd__buf_2
XFILLER_0_2_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput214 net214 vssd1 vssd1 vccd1 vccd1 gpio_out[17] sky130_fd_sc_hd__buf_2
Xoutput225 net225 vssd1 vssd1 vccd1 vccd1 gpio_out[28] sky130_fd_sc_hd__buf_2
XFILLER_0_140_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput236 net236 vssd1 vssd1 vccd1 vccd1 gpio_out[8] sky130_fd_sc_hd__buf_2
XFILLER_0_2_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput247 net247 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[19] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_58_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput258 net258 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[3] sky130_fd_sc_hd__buf_2
XANTENNA__08240__C1 net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07594__A1 net1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11390__A2 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07962_ net613 _03900_ _03902_ vssd1 vssd1 vccd1 vccd1 _03904_ sky130_fd_sc_hd__a21oi_4
XANTENNA__08218__S0 net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11438__C net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09701_ _02954_ _04477_ _05126_ _05640_ _05642_ vssd1 vssd1 vccd1 vccd1 _05643_ sky130_fd_sc_hd__a311o_1
X_06913_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[164\] net782
+ net750 _02854_ vssd1 vssd1 vccd1 vccd1 _02855_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_147_3392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11678__B1 net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07893_ net1187 team_03_WB.instance_to_wrap.core.register_file.registers_state\[367\]
+ net877 _03834_ vssd1 vssd1 vccd1 vccd1 _03835_ sky130_fd_sc_hd__a31o_1
XANTENNA__11142__A2 net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08543__B1 net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09632_ team_03_WB.instance_to_wrap.core.decoder.inst\[28\] net1021 net535 _05571_
+ vssd1 vssd1 vccd1 vccd1 _05574_ sky130_fd_sc_hd__o2bb2a_1
XPHY_EDGE_ROW_74_Left_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06844_ net1196 vssd1 vssd1 vccd1 vccd1 _02787_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_104_2506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09205__A net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_2517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09563_ _05178_ _05180_ _05503_ vssd1 vssd1 vccd1 vccd1 _05505_ sky130_fd_sc_hd__or3_1
XANTENNA__09099__A1 net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15063__1449 vssd1 vssd1 vccd1 vccd1 _15063__1449/HI net1449 sky130_fd_sc_hd__conb_1
XFILLER_0_37_1150 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_172_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08514_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[959\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[927\]
+ net950 vssd1 vssd1 vccd1 vccd1 _04456_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_19_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_907 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09494_ net570 _05383_ vssd1 vssd1 vccd1 vccd1 _05436_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_121_2853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_121_2864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10653__A1 team_03_WB.instance_to_wrap.CPU_DAT_O\[8\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_93_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11850__A0 net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08445_ net1228 team_03_WB.instance_to_wrap.core.register_file.registers_state\[732\]
+ net953 team_03_WB.instance_to_wrap.core.register_file.registers_state\[764\] net933
+ vssd1 vssd1 vccd1 vccd1 _04387_ sky130_fd_sc_hd__o221a_1
XANTENNA__09859__B net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout430_A _04079_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_173_3920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1172_A net1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_173_3931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout528_A _06309_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08376_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[950\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[918\]
+ net970 vssd1 vssd1 vccd1 vccd1 _04318_ sky130_fd_sc_hd__mux2_1
XFILLER_0_162_124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07012__X _02954_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11602__A0 net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07327_ _03265_ _03268_ net822 vssd1 vssd1 vccd1 vccd1 _03269_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_45_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_83_Left_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout316_X net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1437_A net1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1058_X net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09810__A3 net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07258_ net1176 team_03_WB.instance_to_wrap.core.register_file.registers_state\[456\]
+ net774 team_03_WB.instance_to_wrap.core.register_file.registers_state\[488\] net1150
+ vssd1 vssd1 vccd1 vccd1 _03200_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_30_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07821__A2 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_143_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout897_A net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07189_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[1011\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[979\]
+ net762 vssd1 vssd1 vccd1 vccd1 _03131_ sky130_fd_sc_hd__mux2_1
XANTENNA__09023__A1 net1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1225_X net1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11905__A1 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1406 net1407 vssd1 vssd1 vccd1 vccd1 net1406 sky130_fd_sc_hd__buf_4
Xfanout1417 net1418 vssd1 vssd1 vccd1 vccd1 net1417 sky130_fd_sc_hd__buf_2
Xfanout430 _04079_ vssd1 vssd1 vccd1 vccd1 net430 sky130_fd_sc_hd__clkbuf_2
Xfanout1428 net1429 vssd1 vssd1 vccd1 vccd1 net1428 sky130_fd_sc_hd__buf_4
XANTENNA__08003__B _03943_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout441 _06819_ vssd1 vssd1 vccd1 vccd1 net441 sky130_fd_sc_hd__buf_6
Xfanout452 net453 vssd1 vssd1 vccd1 vccd1 net452 sky130_fd_sc_hd__clkbuf_4
Xfanout463 net481 vssd1 vssd1 vccd1 vccd1 net463 sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_92_Left_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout852_X net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07337__A1 team_03_WB.instance_to_wrap.core.decoder.inst\[29\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout474 net476 vssd1 vssd1 vccd1 vccd1 net474 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout485 _06779_ vssd1 vssd1 vccd1 vccd1 net485 sky130_fd_sc_hd__buf_4
XANTENNA__11133__A2 net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout496 net517 vssd1 vssd1 vccd1 vccd1 net496 sky130_fd_sc_hd__buf_2
X_12910_ net1310 vssd1 vssd1 vccd1 vccd1 _00674_ sky130_fd_sc_hd__inv_2
X_13890_ clknet_leaf_173_wb_clk_i _01654_ _00255_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[244\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_159_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14729__Q team_03_WB.instance_to_wrap.core.decoder.inst\[26\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12841_ net1253 vssd1 vssd1 vccd1 vccd1 _00605_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_17_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12094__B1 net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12772_ net1366 vssd1 vssd1 vccd1 vccd1 _00536_ sky130_fd_sc_hd__inv_2
XANTENNA__08298__C1 net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_167_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14511_ clknet_leaf_138_wb_clk_i _02275_ _00876_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[865\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10644__A1 team_03_WB.instance_to_wrap.CPU_DAT_O\[17\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_11723_ net596 _06469_ net457 _06808_ net1798 vssd1 vssd1 vccd1 vccd1 _01813_ sky130_fd_sc_hd__a32o_1
XANTENNA__08932__S1 net1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11841__B1 net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14442_ clknet_leaf_6_wb_clk_i _02206_ _00807_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[796\]
+ sky130_fd_sc_hd__dfrtp_1
X_11654_ net2486 _06620_ net342 vssd1 vssd1 vccd1 vccd1 _01879_ sky130_fd_sc_hd__mux2_1
XANTENNA__10708__B net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10605_ net1702 team_03_WB.instance_to_wrap.CPU_DAT_O\[24\] _06304_ vssd1 vssd1 vccd1
+ vccd1 _02523_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14373_ clknet_leaf_40_wb_clk_i _02137_ _00738_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[727\]
+ sky130_fd_sc_hd__dfrtp_1
X_11585_ net300 net2393 net448 vssd1 vssd1 vccd1 vccd1 _01944_ sky130_fd_sc_hd__mux2_1
XANTENNA__07499__S1 net1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_859 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10947__A2 _05757_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13324_ net1316 vssd1 vssd1 vccd1 vccd1 _01088_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_347 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10536_ net161 net1034 net1026 net1600 vssd1 vssd1 vccd1 vccd1 _02574_ sky130_fd_sc_hd__a22o_1
XFILLER_0_101_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_108_Right_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_1098 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13255_ net1399 vssd1 vssd1 vccd1 vccd1 _01019_ sky130_fd_sc_hd__inv_2
XANTENNA__10724__A _05833_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10467_ _02775_ _06279_ net286 vssd1 vssd1 vccd1 vccd1 _06280_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06921__B net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_199 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12206_ net1510 vssd1 vssd1 vccd1 vccd1 _02347_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08222__C1 net1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_57_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_57_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_20_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_36_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13186_ net1289 vssd1 vssd1 vccd1 vccd1 _00950_ sky130_fd_sc_hd__inv_2
X_10398_ team_03_WB.instance_to_wrap.core.pc.current_pc\[14\] _06141_ team_03_WB.instance_to_wrap.core.pc.current_pc\[15\]
+ vssd1 vssd1 vccd1 vccd1 _06224_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07576__A1 net1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11372__A2 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08773__B1 net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12137_ net1690 vssd1 vssd1 vccd1 vccd1 _02416_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__10580__B1 net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_1020 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12068_ net264 net2689 net358 vssd1 vssd1 vccd1 vccd1 _01478_ sky130_fd_sc_hd__mux2_1
X_11019_ net1249 net833 _06478_ net669 vssd1 vssd1 vccd1 vccd1 _06583_ sky130_fd_sc_hd__or4_1
XFILLER_0_159_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12085__B1 net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14709_ clknet_leaf_33_wb_clk_i _02473_ _01074_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.control_logic.instruction\[6\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__11832__B1 net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_119 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_288 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_20 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_828 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08230_ net1232 team_03_WB.instance_to_wrap.core.register_file.registers_state\[721\]
+ net962 team_03_WB.instance_to_wrap.core.register_file.registers_state\[753\] net936
+ vssd1 vssd1 vccd1 vccd1 _04172_ sky130_fd_sc_hd__o221a_1
XFILLER_0_157_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_144_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_145_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_166_1002 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_86 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_166_1024 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08161_ _04095_ _04102_ net871 vssd1 vssd1 vccd1 vccd1 _04103_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07112_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[1\] net800
+ net731 _03053_ vssd1 vssd1 vccd1 vccd1 _03054_ sky130_fd_sc_hd__o211a_1
X_08092_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[26\] net760
+ net739 _04033_ vssd1 vssd1 vccd1 vccd1 _04034_ sky130_fd_sc_hd__a211o_1
XFILLER_0_28_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11060__B2 net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08461__C1 net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_818 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_464 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_141_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07043_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[419\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[387\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[291\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[259\]
+ net780 net1133 vssd1 vssd1 vccd1 vccd1 _02985_ sky130_fd_sc_hd__mux4_1
Xclkload40 clknet_leaf_20_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload40/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_24_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload51 clknet_leaf_171_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload51/Y sky130_fd_sc_hd__bufinv_16
Xclkload62 clknet_leaf_42_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload62/Y sky130_fd_sc_hd__clkinv_2
XFILLER_0_3_764 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_1951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload73 clknet_leaf_53_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload73/Y sky130_fd_sc_hd__inv_6
XTAP_TAPCELL_ROW_77_1962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload84 clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload84/X sky130_fd_sc_hd__clkbuf_8
XANTENNA__07016__B1 net1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13010__A net1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload95 clknet_leaf_64_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload95/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_3_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08213__C1 net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_149_3432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11899__B1 net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_149_3443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08104__A net1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08994_ net1218 _04932_ _04933_ vssd1 vssd1 vccd1 vccd1 _04936_ sky130_fd_sc_hd__nand3_1
XANTENNA__10571__B1 net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_166_3790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07945_ net1088 team_03_WB.instance_to_wrap.core.register_file.registers_state\[695\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[663\] net793 net744
+ vssd1 vssd1 vccd1 vccd1 _03887_ sky130_fd_sc_hd__o221a_1
XANTENNA__09861__C _05676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout380_A net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout478_A net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12060__S net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07876_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[155\] net783
+ net737 _03817_ vssd1 vssd1 vccd1 vccd1 _03818_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_3_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_162_3698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09615_ _04778_ _05551_ _05555_ _05556_ vssd1 vssd1 vccd1 vccd1 _05557_ sky130_fd_sc_hd__o211ai_1
XANTENNA__11184__B net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06827_ team_03_WB.instance_to_wrap.core.pc.current_pc\[25\] vssd1 vssd1 vccd1 vccd1
+ _02770_ sky130_fd_sc_hd__inv_2
XANTENNA__10874__A1 team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[18\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout266_X net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout645_A _06458_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1387_A net1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09546_ net569 _05487_ net321 vssd1 vssd1 vccd1 vccd1 _05488_ sky130_fd_sc_hd__o21a_1
XANTENNA__12076__B1 net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08819__A1 net1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10626__A1 team_03_WB.instance_to_wrap.CPU_DAT_O\[3\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11823__B1 net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09477_ _05415_ _05418_ net563 vssd1 vssd1 vccd1 vccd1 _05419_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout812_A net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1175_X net1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11404__S net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08428_ net1228 team_03_WB.instance_to_wrap.core.register_file.registers_state\[730\]
+ net964 team_03_WB.instance_to_wrap.core.register_file.registers_state\[762\] net937
+ vssd1 vssd1 vccd1 vccd1 _04370_ sky130_fd_sc_hd__o221a_1
XFILLER_0_148_496 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_647 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkload1 clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload1/Y sky130_fd_sc_hd__inv_6
XFILLER_0_62_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08359_ net1236 team_03_WB.instance_to_wrap.core.register_file.registers_state\[214\]
+ net970 team_03_WB.instance_to_wrap.core.register_file.registers_state\[246\] net939
+ vssd1 vssd1 vccd1 vccd1 _04301_ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout1342_X net1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07255__B1 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11370_ net508 net637 _06737_ net402 net2002 vssd1 vssd1 vccd1 vccd1 _02095_ sky130_fd_sc_hd__a32o_1
XFILLER_0_6_591 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10321_ team_03_WB.instance_to_wrap.core.pc.current_pc\[28\] _06151_ team_03_WB.instance_to_wrap.core.pc.current_pc\[29\]
+ vssd1 vssd1 vccd1 vccd1 _06161_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_15_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_486 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07270__A3 net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13040_ net1412 vssd1 vssd1 vccd1 vccd1 _00804_ sky130_fd_sc_hd__inv_2
X_10252_ _06093_ vssd1 vssd1 vccd1 vccd1 _06094_ sky130_fd_sc_hd__inv_2
XANTENNA__11359__B _06473_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12000__B1 net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08014__A net1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07102__S0 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11354__A2 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10183_ _04619_ team_03_WB.instance_to_wrap.core.pc.current_pc\[7\] net675 vssd1
+ vssd1 vccd1 vccd1 _06025_ sky130_fd_sc_hd__mux2_1
Xfanout1203 net1204 vssd1 vssd1 vccd1 vccd1 net1203 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08949__A net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1214 net1216 vssd1 vssd1 vccd1 vccd1 net1214 sky130_fd_sc_hd__clkbuf_8
XANTENNA__09544__S net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1225 team_03_WB.instance_to_wrap.core.decoder.inst\[16\] vssd1 vssd1 vccd1
+ vccd1 net1225 sky130_fd_sc_hd__buf_4
Xfanout1236 net1238 vssd1 vssd1 vccd1 vccd1 net1236 sky130_fd_sc_hd__clkbuf_4
Xfanout1247 net1250 vssd1 vssd1 vccd1 vccd1 net1247 sky130_fd_sc_hd__buf_4
X_14991_ clknet_leaf_41_wb_clk_i net39 _01356_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input39_A gpio_in[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10550__Y _06293_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1258 net1259 vssd1 vssd1 vccd1 vccd1 net1258 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_31_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout271 _06491_ vssd1 vssd1 vccd1 vccd1 net271 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_31_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1269 net1270 vssd1 vssd1 vccd1 vccd1 net1269 sky130_fd_sc_hd__buf_4
Xfanout282 net283 vssd1 vssd1 vccd1 vccd1 net282 sky130_fd_sc_hd__buf_2
XANTENNA__11375__A net1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13942_ clknet_leaf_176_wb_clk_i _01706_ _00307_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[296\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout293 net294 vssd1 vssd1 vccd1 vccd1 net293 sky130_fd_sc_hd__buf_2
XANTENNA__09180__B1 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13873_ clknet_leaf_140_wb_clk_i _01637_ _00238_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[227\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_175_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_175_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__07621__A1_N net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1081 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12824_ net1379 vssd1 vssd1 vccd1 vccd1 _00588_ sky130_fd_sc_hd__inv_2
XFILLER_0_9_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_104_wb_clk_i clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_104_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_5_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11814__B1 net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12755_ net1256 vssd1 vssd1 vccd1 vccd1 _00519_ sky130_fd_sc_hd__inv_2
XFILLER_0_96_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_167_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10719__A _05596_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11314__S net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11706_ _06748_ net383 net340 net2161 vssd1 vssd1 vccd1 vccd1 _01828_ sky130_fd_sc_hd__a22o_1
XANTENNA__11290__A1 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_155_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12686_ net1274 vssd1 vssd1 vccd1 vccd1 _00450_ sky130_fd_sc_hd__inv_2
XANTENNA__10438__B _06136_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14425_ clknet_leaf_175_wb_clk_i _02189_ _00790_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[779\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_71_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_170_904 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11637_ _06711_ net385 net349 net2511 vssd1 vssd1 vccd1 vccd1 _01895_ sky130_fd_sc_hd__a22o_1
XFILLER_0_142_606 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08669__S0 net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12934__A net1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_122 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09786__A2 _05384_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11042__B2 net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14356_ clknet_leaf_132_wb_clk_i _02120_ _00721_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[710\]
+ sky130_fd_sc_hd__dfrtp_1
X_11568_ net2260 net484 _06797_ net507 vssd1 vssd1 vccd1 vccd1 _01957_ sky130_fd_sc_hd__a22o_1
XFILLER_0_107_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13307_ net1334 vssd1 vssd1 vccd1 vccd1 _01071_ sky130_fd_sc_hd__inv_2
XANTENNA__14922__Q team_03_WB.instance_to_wrap.CPU_DAT_O\[9\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold708 team_03_WB.instance_to_wrap.core.register_file.registers_state\[335\] vssd1
+ vssd1 vccd1 vccd1 net2201 sky130_fd_sc_hd__dlygate4sd3_1
X_10519_ net148 net1031 net1023 net1696 vssd1 vssd1 vccd1 vccd1 _02591_ sky130_fd_sc_hd__a22o_1
Xhold719 team_03_WB.instance_to_wrap.core.register_file.registers_state\[370\] vssd1
+ vssd1 vccd1 vccd1 net2212 sky130_fd_sc_hd__dlygate4sd3_1
X_14287_ clknet_leaf_135_wb_clk_i _02051_ _00652_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[641\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11499_ _06620_ net2481 net389 vssd1 vssd1 vccd1 vccd1 _02007_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15062__1448 vssd1 vssd1 vccd1 vccd1 _15062__1448/HI net1448 sky130_fd_sc_hd__conb_1
XPHY_EDGE_ROW_139_Left_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11269__B net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13238_ net1257 vssd1 vssd1 vccd1 vccd1 _01002_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_55_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11984__S net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13169_ net1270 vssd1 vssd1 vccd1 vccd1 _00933_ sky130_fd_sc_hd__inv_2
XANTENNA__11896__A3 net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_144_3340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_44 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11285__A net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07730_ _03670_ _03671_ net1165 vssd1 vssd1 vccd1 vccd1 _03672_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_137_77 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_140_3248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09710__A2 _05041_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07661_ net616 _03601_ vssd1 vssd1 vccd1 vccd1 _03603_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_140_3259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07182__C1 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11435__D net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_148_Left_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09400_ _03352_ _04475_ vssd1 vssd1 vccd1 vccd1 _05342_ sky130_fd_sc_hd__and2_1
XANTENNA__12058__A0 _06624_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07592_ _03531_ _03533_ net814 vssd1 vssd1 vccd1 vccd1 _03534_ sky130_fd_sc_hd__a21o_1
XFILLER_0_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09331_ _05230_ _05272_ vssd1 vssd1 vccd1 vccd1 _05273_ sky130_fd_sc_hd__and2_1
XFILLER_0_47_203 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09262_ _05198_ _05203_ vssd1 vssd1 vccd1 vccd1 _05204_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_118_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11820__A3 net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08213_ net1232 team_03_WB.instance_to_wrap.core.register_file.registers_state\[81\]
+ net962 team_03_WB.instance_to_wrap.core.register_file.registers_state\[113\] net919
+ vssd1 vssd1 vccd1 vccd1 _04155_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_138_3199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09226__A1 _03314_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09193_ net544 net434 net429 net592 vssd1 vssd1 vccd1 vccd1 _05135_ sky130_fd_sc_hd__or4_1
XFILLER_0_8_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_160_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10067__C net1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08144_ _02799_ _02801_ _02810_ _02812_ net1049 vssd1 vssd1 vccd1 vccd1 _04086_ sky130_fd_sc_hd__a221o_2
XANTENNA__07237__B1 net1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07938__A net1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08533__S net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06842__A net1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_116_2752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07788__A1 net1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_157_Left_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08985__B1 net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_2763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload140 clknet_leaf_74_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload140/Y sky130_fd_sc_hd__clkinv_4
XANTENNA__12055__S net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08075_ _04010_ _04011_ _04016_ net1163 vssd1 vssd1 vccd1 vccd1 _04017_ sky130_fd_sc_hd__o22a_1
Xclkload151 clknet_leaf_80_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload151/Y sky130_fd_sc_hd__inv_6
XFILLER_0_3_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1135_A net1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload162 clknet_leaf_106_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload162/Y sky130_fd_sc_hd__clkinv_2
XFILLER_0_101_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload173 clknet_leaf_89_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload173/Y sky130_fd_sc_hd__inv_6
XTAP_TAPCELL_ROW_168_3830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07026_ net1196 team_03_WB.instance_to_wrap.core.register_file.registers_state\[611\]
+ net883 _02967_ vssd1 vssd1 vccd1 vccd1 _02968_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_8_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11336__A2 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1302_A net1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_164_3738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11887__A3 net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_164_3749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold13 team_03_WB.instance_to_wrap.core.register_file.registers_state\[982\] vssd1
+ vssd1 vccd1 vccd1 net1506 sky130_fd_sc_hd__dlygate4sd3_1
X_08977_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[873\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[841\]
+ net986 vssd1 vssd1 vccd1 vccd1 _04919_ sky130_fd_sc_hd__mux2_1
Xhold24 team_03_WB.instance_to_wrap.core.register_file.registers_state\[942\] vssd1
+ vssd1 vccd1 vccd1 net1517 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout762_A net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold35 team_03_WB.instance_to_wrap.core.register_file.registers_state\[947\] vssd1
+ vssd1 vccd1 vccd1 net1528 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout383_X net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold46 team_03_WB.instance_to_wrap.core.register_file.registers_state\[980\] vssd1
+ vssd1 vccd1 vccd1 net1539 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_2_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_2_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xhold57 team_03_WB.instance_to_wrap.core.register_file.registers_state\[943\] vssd1
+ vssd1 vccd1 vccd1 net1550 sky130_fd_sc_hd__dlygate4sd3_1
X_07928_ net1181 team_03_WB.instance_to_wrap.core.register_file.registers_state\[183\]
+ net892 net1128 vssd1 vssd1 vccd1 vccd1 _03870_ sky130_fd_sc_hd__a211o_1
Xhold68 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1007\] vssd1
+ vssd1 vccd1 vccd1 net1561 sky130_fd_sc_hd__dlygate4sd3_1
Xhold79 team_03_WB.instance_to_wrap.core.register_file.registers_state\[964\] vssd1
+ vssd1 vccd1 vccd1 net1572 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_166_Left_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07859_ net1202 team_03_WB.instance_to_wrap.core.register_file.registers_state\[571\]
+ net886 vssd1 vssd1 vccd1 vccd1 _03801_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout648_X net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10870_ _06465_ _06466_ _06467_ net585 vssd1 vssd1 vccd1 vccd1 _06468_ sky130_fd_sc_hd__o211a_4
XFILLER_0_97_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09529_ _05469_ _05470_ net563 vssd1 vssd1 vccd1 vccd1 _05471_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout815_X net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07476__B1 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11272__A1 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12540_ net1409 vssd1 vssd1 vccd1 vccd1 _00304_ sky130_fd_sc_hd__inv_2
XANTENNA__11361__C _06477_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08673__C1 net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08009__A net1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_978 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12471_ net1392 vssd1 vssd1 vccd1 vccd1 _00235_ sky130_fd_sc_hd__inv_2
XFILLER_0_81_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10826__X _06430_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12754__A net1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14210_ clknet_leaf_174_wb_clk_i _01974_ _00575_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[564\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_62_740 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11422_ net270 net2506 net396 vssd1 vssd1 vccd1 vccd1 _02060_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07779__A1 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14141_ clknet_leaf_25_wb_clk_i _01905_ _00506_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[495\]
+ sky130_fd_sc_hd__dfrtp_1
X_11353_ _06446_ net711 _06561_ vssd1 vssd1 vccd1 vccd1 _06729_ sky130_fd_sc_hd__and3_1
XANTENNA__10783__B1 _06293_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07059__S net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10304_ team_03_WB.instance_to_wrap.core.pc.current_pc\[21\] team_03_WB.instance_to_wrap.core.pc.current_pc\[20\]
+ _06145_ vssd1 vssd1 vccd1 vccd1 _06146_ sky130_fd_sc_hd__and3_1
XFILLER_0_21_147 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14072_ clknet_leaf_19_wb_clk_i _01836_ _00437_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[426\]
+ sky130_fd_sc_hd__dfrtp_1
X_11284_ net516 net645 _06709_ net411 net2174 vssd1 vssd1 vccd1 vccd1 _02153_ sky130_fd_sc_hd__a32o_1
XFILLER_0_120_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13023_ net1287 vssd1 vssd1 vccd1 vccd1 _00787_ sky130_fd_sc_hd__inv_2
X_10235_ _06073_ _06074_ vssd1 vssd1 vccd1 vccd1 _06077_ sky130_fd_sc_hd__or2_1
XANTENNA__10535__B1 net1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1000 _04085_ vssd1 vssd1 vccd1 vccd1 net1000 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11878__A3 net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1011 net1012 vssd1 vssd1 vccd1 vccd1 net1011 sky130_fd_sc_hd__clkbuf_4
Xfanout1022 _02803_ vssd1 vssd1 vccd1 vccd1 net1022 sky130_fd_sc_hd__clkbuf_2
Xfanout1033 net1035 vssd1 vssd1 vccd1 vccd1 net1033 sky130_fd_sc_hd__clkbuf_2
X_10166_ _06006_ _06007_ vssd1 vssd1 vccd1 vccd1 _06008_ sky130_fd_sc_hd__or2_1
Xfanout1044 _02793_ vssd1 vssd1 vccd1 vccd1 net1044 sky130_fd_sc_hd__buf_4
XANTENNA__07951__A1 net1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1055 net1060 vssd1 vssd1 vccd1 vccd1 net1055 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11309__S net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1066 net1069 vssd1 vssd1 vccd1 vccd1 net1066 sky130_fd_sc_hd__clkbuf_8
Xfanout1077 net1080 vssd1 vssd1 vccd1 vccd1 net1077 sky130_fd_sc_hd__clkbuf_2
X_14974_ clknet_leaf_92_wb_clk_i _02726_ _01339_ vssd1 vssd1 vccd1 vccd1 net226 sky130_fd_sc_hd__dfrtp_1
X_10097_ _02832_ _02926_ _05940_ vssd1 vssd1 vccd1 vccd1 _05941_ sky130_fd_sc_hd__or3b_1
Xfanout1088 net1089 vssd1 vssd1 vccd1 vccd1 net1088 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_107_25 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1099 net1101 vssd1 vssd1 vccd1 vccd1 net1099 sky130_fd_sc_hd__buf_2
XANTENNA__10838__A1 net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13925_ clknet_leaf_37_wb_clk_i _01689_ _00290_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[279\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07703__A1 net1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08900__B1 net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload4_A clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13856_ clknet_leaf_191_wb_clk_i _01620_ _00221_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[210\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06927__A net1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09303__A _04591_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14917__Q team_03_WB.instance_to_wrap.CPU_DAT_O\[4\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_12807_ net1368 vssd1 vssd1 vccd1 vccd1 _00571_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_48_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09456__A1 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13787_ clknet_leaf_158_wb_clk_i _01551_ _00152_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[141\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_48_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10999_ net1044 net836 net278 net670 vssd1 vssd1 vccd1 vccd1 _06572_ sky130_fd_sc_hd__and4_1
XFILLER_0_84_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07467__B1 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12738_ net1351 vssd1 vssd1 vccd1 vccd1 _00502_ sky130_fd_sc_hd__inv_2
XFILLER_0_45_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11271__C net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10168__B net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11979__S net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_44_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12669_ net1383 vssd1 vssd1 vccd1 vccd1 _00433_ sky130_fd_sc_hd__inv_2
XFILLER_0_167_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14408_ clknet_leaf_9_wb_clk_i _02172_ _00773_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[762\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09759__A2 net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07758__A net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_2346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_160_Right_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_72_wb_clk_i clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_72_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_13_604 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_2357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08206__X _04148_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11566__A2 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_17_wb_clk_i_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__08967__B1 net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14339_ clknet_leaf_31_wb_clk_i _02103_ _00704_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[693\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold505 _02596_ vssd1 vssd1 vccd1 vccd1 net1998 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10184__A _03430_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold516 team_03_WB.instance_to_wrap.core.register_file.registers_state\[868\] vssd1
+ vssd1 vccd1 vccd1 net2009 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06978__C1 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07865__S1 net1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold527 team_03_WB.instance_to_wrap.core.register_file.registers_state\[739\] vssd1
+ vssd1 vccd1 vccd1 net2020 sky130_fd_sc_hd__dlygate4sd3_1
Xhold538 team_03_WB.instance_to_wrap.core.register_file.registers_state\[238\] vssd1
+ vssd1 vccd1 vccd1 net2031 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold549 team_03_WB.instance_to_wrap.core.register_file.registers_state\[366\] vssd1
+ vssd1 vccd1 vccd1 net2042 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09067__S0 net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08900_ net1239 team_03_WB.instance_to_wrap.core.register_file.registers_state\[332\]
+ net981 team_03_WB.instance_to_wrap.core.register_file.registers_state\[364\] net1076
+ vssd1 vssd1 vccd1 vccd1 _04842_ sky130_fd_sc_hd__o221a_1
X_09880_ _05821_ vssd1 vssd1 vccd1 vccd1 _05822_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_111_2660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_70_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10912__A net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10526__B1 net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08831_ net561 _04740_ _04772_ vssd1 vssd1 vccd1 vccd1 _04773_ sky130_fd_sc_hd__or3_1
Xhold1205 team_03_WB.instance_to_wrap.core.register_file.registers_state\[82\] vssd1
+ vssd1 vccd1 vccd1 net2698 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_57_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1216 team_03_WB.instance_to_wrap.core.register_file.registers_state\[93\] vssd1
+ vssd1 vccd1 vccd1 net2709 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11219__S net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08762_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[931\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[899\]
+ net980 vssd1 vssd1 vccd1 vccd1 _04704_ sky130_fd_sc_hd__mux2_1
Xhold1227 team_03_WB.instance_to_wrap.core.register_file.registers_state\[109\] vssd1
+ vssd1 vccd1 vccd1 net2720 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08876__X _04818_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1238 team_03_WB.instance_to_wrap.core.register_file.registers_state\[735\] vssd1
+ vssd1 vccd1 vccd1 net2731 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11446__C net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1249 team_03_WB.instance_to_wrap.core.register_file.registers_state\[111\] vssd1
+ vssd1 vccd1 vccd1 net2742 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10829__A1 net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07713_ net1104 team_03_WB.instance_to_wrap.core.register_file.registers_state\[429\]
+ net899 vssd1 vssd1 vccd1 vccd1 _03655_ sky130_fd_sc_hd__or3_1
XFILLER_0_135_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08693_ net940 _04633_ _04634_ vssd1 vssd1 vccd1 vccd1 _04635_ sky130_fd_sc_hd__o21a_1
XFILLER_0_79_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_147 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11743__A net1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07644_ net818 _03577_ net723 vssd1 vssd1 vccd1 vccd1 _03586_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_68_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07575_ net1189 team_03_WB.instance_to_wrap.core.register_file.registers_state\[984\]
+ vssd1 vssd1 vccd1 vccd1 _03517_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout343_A _06805_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1085_A net1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09314_ _04711_ _05255_ vssd1 vssd1 vccd1 vccd1 _05256_ sky130_fd_sc_hd__nor2_1
XANTENNA_clkbuf_leaf_56_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__10057__A2 net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07458__B1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11254__A1 net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08655__C1 net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_157_3597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_2803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09245_ _05185_ _05186_ vssd1 vssd1 vccd1 vccd1 _05187_ sky130_fd_sc_hd__nand2_1
XFILLER_0_63_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout510_A net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout608_A net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06843__Y _02786_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_291 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09176_ net436 net428 _05041_ net546 vssd1 vssd1 vccd1 vccd1 _05118_ sky130_fd_sc_hd__o31a_1
XFILLER_0_133_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08958__B1 net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08127_ net722 _04041_ _04047_ _04068_ vssd1 vssd1 vccd1 vccd1 _04069_ sky130_fd_sc_hd__o31a_4
XANTENNA__10094__A _05833_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09080__C1 net1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1138_X net1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_892 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08058_ net1090 team_03_WB.instance_to_wrap.core.register_file.registers_state\[374\]
+ net895 vssd1 vssd1 vccd1 vccd1 _04000_ sky130_fd_sc_hd__or3_1
XFILLER_0_3_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout598_X net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout977_A net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07009_ net1020 _02943_ _02947_ vssd1 vssd1 vccd1 vccd1 _02951_ sky130_fd_sc_hd__or3b_1
XANTENNA__10517__B1 net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08186__A1 net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1305_X net1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08499__A net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09094__S net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10020_ net75 net74 vssd1 vssd1 vccd1 vccd1 _05898_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout765_X net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07933__A1 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_95_wb_clk_i_A clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout932_X net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11971_ net634 _06748_ net466 net365 net2522 vssd1 vssd1 vccd1 vccd1 _01572_ sky130_fd_sc_hd__a32o_1
XANTENNA__09686__B2 net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13710_ clknet_leaf_131_wb_clk_i _01474_ _00075_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[64\]
+ sky130_fd_sc_hd__dfrtp_1
X_10922_ net690 _05706_ _06401_ vssd1 vssd1 vccd1 vccd1 _06510_ sky130_fd_sc_hd__a21oi_1
XANTENNA__15125__A net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14690_ clknet_leaf_56_wb_clk_i _02454_ _01055_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.ADR_I\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_15061__1447 vssd1 vssd1 vccd1 vccd1 _15061__1447/HI net1447 sky130_fd_sc_hd__conb_1
X_13641_ net1424 vssd1 vssd1 vccd1 vccd1 _01405_ sky130_fd_sc_hd__inv_2
X_10853_ net691 _05623_ net585 vssd1 vssd1 vccd1 vccd1 _06452_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_39_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07449__A0 _03389_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10048__A2 net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13572_ net1404 vssd1 vssd1 vccd1 vccd1 _01336_ sky130_fd_sc_hd__inv_2
XANTENNA__08646__C1 net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10784_ _06393_ _06391_ _06392_ vssd1 vssd1 vccd1 vccd1 _06394_ sky130_fd_sc_hd__and3b_4
XFILLER_0_27_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08110__A1 net1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11799__S net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12523_ net1297 vssd1 vssd1 vccd1 vccd1 _00287_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_23_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10556__X _06299_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12484__A net1376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_403 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_559 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07578__A net1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12454_ net1299 vssd1 vssd1 vccd1 vccd1 _00218_ sky130_fd_sc_hd__inv_2
XFILLER_0_124_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10716__B net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11548__A2 net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11405_ _06430_ net2616 net399 vssd1 vssd1 vccd1 vccd1 _02075_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08413__A2 net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12385_ net1290 vssd1 vssd1 vccd1 vccd1 _00149_ sky130_fd_sc_hd__inv_2
XFILLER_0_78_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10756__B1 net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14124_ clknet_leaf_21_wb_clk_i _01888_ _00489_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[478\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_50_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11336_ net498 net628 _06720_ net400 net2202 vssd1 vssd1 vccd1 vccd1 _02112_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_91_2243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_91_2254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14055_ clknet_leaf_108_wb_clk_i _01819_ _00420_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[409\]
+ sky130_fd_sc_hd__dfrtp_1
X_11267_ net1248 net839 net299 net671 vssd1 vssd1 vccd1 vccd1 _06701_ sky130_fd_sc_hd__and4_1
XANTENNA__10508__B1 net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15099__1482 vssd1 vssd1 vccd1 vccd1 _15099__1482/HI net1482 sky130_fd_sc_hd__conb_1
XFILLER_0_123_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08177__A1 net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07517__S net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13006_ net1269 vssd1 vssd1 vccd1 vccd1 _00770_ sky130_fd_sc_hd__inv_2
X_10218_ _06057_ _06059_ vssd1 vssd1 vccd1 vccd1 _06060_ sky130_fd_sc_hd__and2_1
X_11198_ team_03_WB.instance_to_wrap.core.decoder.inst\[11\] _06394_ _06455_ vssd1
+ vssd1 vccd1 vccd1 _06680_ sky130_fd_sc_hd__nand3_4
XANTENNA__07924__A1 net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_190_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_190_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_10149_ _03138_ _05990_ vssd1 vssd1 vccd1 vccd1 _05991_ sky130_fd_sc_hd__and2_1
XANTENNA__09677__A1 _03391_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14957_ clknet_leaf_100_wb_clk_i _02709_ _01322_ vssd1 vssd1 vccd1 vccd1 net209 sky130_fd_sc_hd__dfrtp_1
XANTENNA__07137__C1 net1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06928__Y _02870_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11563__A net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13908_ clknet_leaf_134_wb_clk_i _01672_ _00273_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[262\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07688__B1 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14888_ clknet_leaf_65_wb_clk_i _02651_ _01253_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.pc.current_pc\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_159_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13839_ clknet_leaf_137_wb_clk_i _01603_ _00204_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[193\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11236__A1 net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07360_ net1172 team_03_WB.instance_to_wrap.core.register_file.registers_state\[988\]
+ net760 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1020\] net1151
+ vssd1 vssd1 vccd1 vccd1 _03302_ sky130_fd_sc_hd__o221a_1
XFILLER_0_70_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_742 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08101__A1 net1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_764 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07291_ _03229_ _03232_ net825 vssd1 vssd1 vccd1 vccd1 _03233_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_143_712 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_3147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10907__A team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[12\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08591__B net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11502__S net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10995__B1 net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09030_ net1244 team_03_WB.instance_to_wrap.core.register_file.registers_state\[720\]
+ net989 team_03_WB.instance_to_wrap.core.register_file.registers_state\[752\] net946
+ vssd1 vssd1 vccd1 vccd1 _04972_ sky130_fd_sc_hd__o221a_1
XFILLER_0_155_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07488__A team_03_WB.instance_to_wrap.core.decoder.inst\[27\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07860__B1 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_99 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11539__A2 net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_564 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_152_3494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_2700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09062__C1 net1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold302 net195 vssd1 vssd1 vccd1 vccd1 net1795 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07838__S1 net1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_20 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold313 team_03_WB.instance_to_wrap.CPU_DAT_O\[22\] vssd1 vssd1 vccd1 vccd1 net1806
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold324 team_03_WB.instance_to_wrap.core.register_file.registers_state\[51\] vssd1
+ vssd1 vccd1 vccd1 net1817 sky130_fd_sc_hd__dlygate4sd3_1
Xhold335 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[20\] vssd1 vssd1 vccd1
+ vccd1 net1828 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold346 team_03_WB.instance_to_wrap.core.register_file.registers_state\[59\] vssd1
+ vssd1 vccd1 vccd1 net1839 sky130_fd_sc_hd__dlygate4sd3_1
Xhold357 team_03_WB.instance_to_wrap.core.register_file.registers_state\[546\] vssd1
+ vssd1 vccd1 vccd1 net1850 sky130_fd_sc_hd__dlygate4sd3_1
X_09932_ _05870_ net1732 net294 vssd1 vssd1 vccd1 vccd1 _02761_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_862 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold368 team_03_WB.instance_to_wrap.core.register_file.registers_state\[417\] vssd1
+ vssd1 vccd1 vccd1 net1861 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_1144 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold379 team_03_WB.instance_to_wrap.core.register_file.registers_state\[298\] vssd1
+ vssd1 vccd1 vccd1 net1872 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08168__A1 net1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout804 net805 vssd1 vssd1 vccd1 vccd1 net804 sky130_fd_sc_hd__buf_4
Xfanout815 net816 vssd1 vssd1 vccd1 vccd1 net815 sky130_fd_sc_hd__buf_4
Xfanout826 _02819_ vssd1 vssd1 vccd1 vccd1 net826 sky130_fd_sc_hd__buf_4
X_09863_ _03947_ net590 net538 vssd1 vssd1 vccd1 vccd1 _05805_ sky130_fd_sc_hd__o21a_1
XANTENNA__10999__D net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout837 _06386_ vssd1 vssd1 vccd1 vccd1 net837 sky130_fd_sc_hd__buf_4
Xfanout848 net849 vssd1 vssd1 vccd1 vccd1 net848 sky130_fd_sc_hd__buf_6
XANTENNA__08112__A net1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout293_A net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07376__C1 net1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout859 net860 vssd1 vssd1 vccd1 vccd1 net859 sky130_fd_sc_hd__buf_4
X_08814_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[801\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[769\]
+ net980 vssd1 vssd1 vccd1 vccd1 _04756_ sky130_fd_sc_hd__mux2_1
Xhold1002 team_03_WB.instance_to_wrap.core.register_file.registers_state\[341\] vssd1
+ vssd1 vccd1 vccd1 net2495 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1013 team_03_WB.instance_to_wrap.core.register_file.registers_state\[650\] vssd1
+ vssd1 vccd1 vccd1 net2506 sky130_fd_sc_hd__dlygate4sd3_1
X_09794_ _05084_ _05091_ _05117_ _05086_ net562 net571 vssd1 vssd1 vccd1 vccd1 _05736_
+ sky130_fd_sc_hd__mux4_2
XANTENNA_fanout1000_A _04085_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1024 team_03_WB.instance_to_wrap.core.register_file.registers_state\[146\] vssd1
+ vssd1 vccd1 vccd1 net2517 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1035 team_03_WB.instance_to_wrap.core.register_file.registers_state\[194\] vssd1
+ vssd1 vccd1 vccd1 net2528 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_139_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1046 team_03_WB.instance_to_wrap.core.register_file.registers_state\[183\] vssd1
+ vssd1 vccd1 vccd1 net2539 sky130_fd_sc_hd__dlygate4sd3_1
X_08745_ net862 _04685_ _04686_ _04684_ vssd1 vssd1 vccd1 vccd1 _04687_ sky130_fd_sc_hd__a31o_1
Xhold1057 team_03_WB.instance_to_wrap.core.register_file.registers_state\[432\] vssd1
+ vssd1 vccd1 vccd1 net2550 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_84_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09668__A1 net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10788__S net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout460_A net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1068 team_03_WB.instance_to_wrap.core.register_file.registers_state\[727\] vssd1
+ vssd1 vccd1 vccd1 net2561 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07128__C1 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1079 team_03_WB.instance_to_wrap.core.register_file.registers_state\[576\] vssd1
+ vssd1 vccd1 vccd1 net2572 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout558_A _03064_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09668__B2 net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11473__A net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07679__B1 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08676_ _04610_ _04611_ _04617_ _04614_ net1068 _02788_ vssd1 vssd1 vccd1 vccd1 _04618_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__08340__A1 net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_159_3637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08340__B2 net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_159_3648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07627_ net1192 net881 team_03_WB.instance_to_wrap.core.register_file.registers_state\[14\]
+ vssd1 vssd1 vccd1 vccd1 _03569_ sky130_fd_sc_hd__a21o_1
XANTENNA__11192__B net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_179_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_67_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout725_A net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12019__A3 net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout346_X net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1088_X net1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_731 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07558_ _03496_ _03499_ net821 vssd1 vssd1 vccd1 vccd1 _03500_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08782__A net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout513_X net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_194 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07489_ net1110 team_03_WB.instance_to_wrap.core.register_file.registers_state\[839\]
+ net803 team_03_WB.instance_to_wrap.core.register_file.registers_state\[871\] net1158
+ vssd1 vssd1 vccd1 vccd1 _03431_ sky130_fd_sc_hd__a221o_1
XFILLER_0_8_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_723 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11412__S net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09228_ _04532_ _05169_ vssd1 vssd1 vccd1 vccd1 _05170_ sky130_fd_sc_hd__or2_2
XFILLER_0_106_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07851__B1 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_907 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09159_ net431 net424 _04503_ net549 vssd1 vssd1 vccd1 vccd1 _05101_ sky130_fd_sc_hd__o31a_1
XFILLER_0_90_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1422_X net1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_161_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12170_ net1609 vssd1 vssd1 vccd1 vccd1 _02383_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__08721__S net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout882_X net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11121_ _06449_ net629 _06634_ vssd1 vssd1 vccd1 vccd1 _06635_ sky130_fd_sc_hd__or3_4
XFILLER_0_7_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold880 team_03_WB.instance_to_wrap.core.register_file.registers_state\[635\] vssd1
+ vssd1 vccd1 vccd1 net2373 sky130_fd_sc_hd__dlygate4sd3_1
Xhold891 team_03_WB.instance_to_wrap.core.register_file.registers_state\[718\] vssd1
+ vssd1 vccd1 vccd1 net2384 sky130_fd_sc_hd__dlygate4sd3_1
X_11052_ net515 net657 _06603_ net423 net2001 vssd1 vssd1 vccd1 vccd1 _02279_ sky130_fd_sc_hd__a32o_1
XANTENNA__11367__B net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08022__A net1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11163__B1 net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07367__C1 net1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10003_ _05888_ net1748 net290 vssd1 vssd1 vccd1 vccd1 _02711_ sky130_fd_sc_hd__mux2_1
XANTENNA__11702__A2 net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10910__B1 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09108__B1 net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input21_A DAT_I[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09552__S net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14811_ clknet_leaf_95_wb_clk_i net1714 _01176_ vssd1 vssd1 vccd1 vccd1 net162 sky130_fd_sc_hd__dfrtp_1
XANTENNA__11383__A net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14742_ clknet_leaf_69_wb_clk_i _02506_ _01107_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_11954_ net622 _06731_ net454 net363 net2046 vssd1 vssd1 vccd1 vccd1 _01589_ sky130_fd_sc_hd__a32o_1
XFILLER_0_98_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10905_ net693 _05697_ net586 vssd1 vssd1 vccd1 vccd1 _06496_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_28_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_128 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14673_ clknet_leaf_87_wb_clk_i _02437_ _01038_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.ADR_I\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_1107 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11885_ net629 _06694_ net461 net372 net2229 vssd1 vssd1 vccd1 vccd1 _01656_ sky130_fd_sc_hd__a32o_1
XPHY_EDGE_ROW_103_Left_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13624_ net1407 vssd1 vssd1 vccd1 vccd1 _01388_ sky130_fd_sc_hd__inv_2
XFILLER_0_156_325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10836_ _06436_ _06437_ _06435_ vssd1 vssd1 vccd1 vccd1 _06438_ sky130_fd_sc_hd__o21a_2
XFILLER_0_67_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09140__X _05082_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11769__A2 net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13555_ net1435 vssd1 vssd1 vccd1 vccd1 _01319_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_15_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08095__B1 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10767_ team_03_WB.instance_to_wrap.core.pc.current_pc\[0\] net604 vssd1 vssd1 vccd1
+ vccd1 _06378_ sky130_fd_sc_hd__or2_1
XFILLER_0_137_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09292__C1 _04953_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11175__C_N net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_857 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_41_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11322__S net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13103__A net1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12506_ net1375 vssd1 vssd1 vccd1 vccd1 _00270_ sky130_fd_sc_hd__inv_2
XFILLER_0_81_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07842__B1 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13486_ net1345 vssd1 vssd1 vccd1 vccd1 _01250_ sky130_fd_sc_hd__inv_2
XFILLER_0_82_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10698_ net1640 net527 net522 _06336_ vssd1 vssd1 vccd1 vccd1 _02462_ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12437_ net1272 vssd1 vssd1 vccd1 vccd1 _00201_ sky130_fd_sc_hd__inv_2
XFILLER_0_106_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10729__B1 net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_152_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_130_3044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_1019 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_3055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12368_ net1409 vssd1 vssd1 vccd1 vccd1 _00132_ sky130_fd_sc_hd__inv_2
XFILLER_0_22_275 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14930__Q team_03_WB.instance_to_wrap.CPU_DAT_O\[17\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_112_Left_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14107_ clknet_leaf_123_wb_clk_i _01871_ _00472_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[461\]
+ sky130_fd_sc_hd__dfrtp_1
X_11319_ _06626_ net2322 net406 vssd1 vssd1 vccd1 vccd1 _02126_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07070__A1 net1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15087_ net1473 vssd1 vssd1 vccd1 vccd1 la_data_out[23] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_39_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12299_ net1282 vssd1 vssd1 vccd1 vccd1 _00063_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_39_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14038_ clknet_leaf_154_wb_clk_i _01802_ _00403_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[392\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11277__B net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07358__C1 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11992__S net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06860_ team_03_WB.instance_to_wrap.core.control_logic.instruction\[6\] team_03_WB.instance_to_wrap.core.control_logic.instruction\[5\]
+ team_03_WB.instance_to_wrap.core.control_logic.instruction\[4\] vssd1 vssd1 vccd1
+ vccd1 _02802_ sky130_fd_sc_hd__nand3b_2
XFILLER_0_98_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08867__A _02937_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09462__S net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07373__A2 net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08570__A1 net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_31 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11293__A net1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08530_ net1062 _04469_ _04470_ vssd1 vssd1 vccd1 vccd1 _04472_ sky130_fd_sc_hd__or3_1
XANTENNA__11457__A1 net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08858__C1 net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_121_Left_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_65_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08461_ net1226 team_03_WB.instance_to_wrap.core.register_file.registers_state\[188\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[156\] net953 net917
+ vssd1 vssd1 vccd1 vccd1 _04403_ sky130_fd_sc_hd__a221o_1
X_07412_ net1175 team_03_WB.instance_to_wrap.core.register_file.registers_state\[596\]
+ vssd1 vssd1 vccd1 vccd1 _03354_ sky130_fd_sc_hd__or2_1
XFILLER_0_9_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_102_2467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_43 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08392_ net865 _04330_ _04333_ vssd1 vssd1 vccd1 vccd1 _04334_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_46_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_2478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_154_3534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07343_ net739 _03281_ _03282_ _03283_ _03284_ vssd1 vssd1 vccd1 vccd1 _03285_ sky130_fd_sc_hd__o32a_1
XFILLER_0_45_323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_174_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_154_3545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09822__A1 _04777_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11232__S net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13013__A net1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09210__B _05146_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07274_ _02872_ _03214_ _03215_ _02870_ _03213_ vssd1 vssd1 vccd1 vccd1 _03216_ sky130_fd_sc_hd__o221a_1
XFILLER_0_45_378 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08107__A net1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_171_3881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09013_ net436 net428 _04953_ net546 vssd1 vssd1 vccd1 vccd1 _04955_ sky130_fd_sc_hd__o31a_1
XANTENNA__07011__A net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_171_3892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_171_884 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15001__Q team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[20\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08389__A1 net1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1048_A net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold110 team_03_WB.instance_to_wrap.core.register_file.registers_state\[965\] vssd1
+ vssd1 vccd1 vccd1 net1603 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07946__A net1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold121 team_03_WB.instance_to_wrap.CPU_DAT_I\[1\] vssd1 vssd1 vccd1 vccd1 net1614
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold132 team_03_WB.instance_to_wrap.core.register_file.registers_state\[13\] vssd1
+ vssd1 vccd1 vccd1 net1625 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06850__A net1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold143 team_03_WB.instance_to_wrap.core.register_file.registers_state\[972\] vssd1
+ vssd1 vccd1 vccd1 net1636 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14840__Q net114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold154 net185 vssd1 vssd1 vccd1 vccd1 net1647 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07061__A1 net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11468__A net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15060__1446 vssd1 vssd1 vccd1 vccd1 _15060__1446/HI net1446 sky130_fd_sc_hd__conb_1
Xhold165 team_03_WB.instance_to_wrap.ADR_I\[14\] vssd1 vssd1 vccd1 vccd1 net1658 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12063__S net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold176 _02512_ vssd1 vssd1 vccd1 vccd1 net1669 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1215_A net1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07600__A3 net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold187 team_03_WB.instance_to_wrap.ADR_I\[6\] vssd1 vssd1 vccd1 vccd1 net1680 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout601 _06299_ vssd1 vssd1 vccd1 vccd1 net601 sky130_fd_sc_hd__clkbuf_4
Xhold198 net117 vssd1 vssd1 vccd1 vccd1 net1691 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout612 _02843_ vssd1 vssd1 vccd1 vccd1 net612 sky130_fd_sc_hd__buf_4
XFILLER_0_10_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09915_ _05646_ _05676_ _05856_ vssd1 vssd1 vccd1 vccd1 _05857_ sky130_fd_sc_hd__and3_1
Xfanout623 net625 vssd1 vssd1 vccd1 vccd1 net623 sky130_fd_sc_hd__clkbuf_2
XANTENNA__10091__B _05596_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09889__A1 net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07349__C1 net1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout634 net638 vssd1 vssd1 vccd1 vccd1 net634 sky130_fd_sc_hd__buf_4
XANTENNA_fanout675_A _05948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09889__B2 _05436_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout296_X net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout645 _06458_ vssd1 vssd1 vccd1 vccd1 net645 sky130_fd_sc_hd__buf_2
Xfanout656 net658 vssd1 vssd1 vccd1 vccd1 net656 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10499__A2 net1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout667 _04818_ vssd1 vssd1 vccd1 vccd1 net667 sky130_fd_sc_hd__buf_4
X_09846_ net540 _05787_ vssd1 vssd1 vccd1 vccd1 _05788_ sky130_fd_sc_hd__nand2_1
XANTENNA__08010__B1 net1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout678 net679 vssd1 vssd1 vccd1 vccd1 net678 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_fanout1003_X net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout689 net690 vssd1 vssd1 vccd1 vccd1 net689 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08561__A1 net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09777_ _05240_ _05241_ vssd1 vssd1 vccd1 vccd1 _05719_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout842_A net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06989_ _02929_ _02930_ vssd1 vssd1 vccd1 vccd1 _02931_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_126_2957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout463_X net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12299__A net1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_126_2968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11407__S net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08728_ net1222 _04668_ _04669_ _04665_ _04667_ vssd1 vssd1 vccd1 vccd1 _04670_ sky130_fd_sc_hd__a32o_1
XANTENNA__09510__B1 net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_25_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout630_X net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08659_ net865 _04599_ _04600_ _04598_ vssd1 vssd1 vccd1 vccd1 _04601_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_1_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout728_X net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11670_ net2545 _06630_ net345 vssd1 vssd1 vccd1 vccd1 _01863_ sky130_fd_sc_hd__mux2_1
XFILLER_0_113_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10621_ net2270 team_03_WB.instance_to_wrap.CPU_DAT_O\[8\] net842 vssd1 vssd1 vccd1
+ vccd1 _02507_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_12_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09813__B2 _05073_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13340_ net1326 vssd1 vssd1 vccd1 vccd1 _01104_ sky130_fd_sc_hd__inv_2
XFILLER_0_106_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10552_ net1144 _06293_ _06292_ vssd1 vssd1 vccd1 vccd1 _06295_ sky130_fd_sc_hd__a21o_2
XANTENNA__07824__B1 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13271_ net1404 vssd1 vssd1 vccd1 vccd1 _01035_ sky130_fd_sc_hd__inv_2
XANTENNA__10974__A3 net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_715 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10483_ net118 net1028 net906 net1628 vssd1 vssd1 vccd1 vccd1 _02626_ sky130_fd_sc_hd__a22o_1
XFILLER_0_84_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_129_wb_clk_i clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_129_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_106_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15010_ clknet_leaf_63_wb_clk_i net58 _01375_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_121_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12222_ net1660 vssd1 vssd1 vccd1 vccd1 _01435_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_122_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input69_A wbs_adr_i[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11384__B1 net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12153_ net1535 vssd1 vssd1 vccd1 vccd1 _02400_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__10282__A _03313_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11104_ net834 net296 vssd1 vssd1 vccd1 vccd1 _06628_ sky130_fd_sc_hd__and2_2
XANTENNA__11097__B net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12084_ net628 _06650_ net459 net440 net1843 vssd1 vssd1 vccd1 vccd1 _01463_ sky130_fd_sc_hd__a32o_1
XFILLER_0_21_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11035_ net710 _06503_ net701 vssd1 vssd1 vccd1 vccd1 _06593_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_34_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08552__A1 net1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11317__S net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11439__B2 net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09727__S1 net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12986_ net1377 vssd1 vssd1 vccd1 vccd1 _00750_ sky130_fd_sc_hd__inv_2
XFILLER_0_99_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08304__A1 net1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14725_ clknet_leaf_53_wb_clk_i _02489_ _01090_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.decoder.inst\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_169_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11937_ _06631_ net2740 net369 vssd1 vssd1 vccd1 vccd1 _01605_ sky130_fd_sc_hd__mux2_1
XANTENNA__11263__D net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14656_ clknet_leaf_192_wb_clk_i _02420_ _01021_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1010\]
+ sky130_fd_sc_hd__dfstp_1
X_11868_ _06527_ net2176 net377 vssd1 vssd1 vccd1 vccd1 _01672_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09311__A _04679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06961__S1 net1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10819_ net311 net310 net317 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[26\]
+ vssd1 vssd1 vccd1 vccd1 _06424_ sky130_fd_sc_hd__a31o_1
X_13607_ net1265 vssd1 vssd1 vccd1 vccd1 _01371_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_60_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08068__B1 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10457__A team_03_WB.instance_to_wrap.core.pc.current_pc\[4\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09804__A1 _02954_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14587_ clknet_leaf_121_wb_clk_i _02351_ _00952_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[941\]
+ sky130_fd_sc_hd__dfstp_1
X_11799_ net2340 _06628_ net329 vssd1 vssd1 vccd1 vccd1 _01739_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_892 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07815__B1 team_03_WB.instance_to_wrap.core.decoder.inst\[31\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13538_ net1317 vssd1 vssd1 vccd1 vccd1 _01302_ sky130_fd_sc_hd__inv_2
XFILLER_0_137_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10176__B net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11987__S net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13469_ net1328 vssd1 vssd1 vccd1 vccd1 _01233_ sky130_fd_sc_hd__inv_2
XANTENNA__09965__B net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12672__A net1402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07830__A3 net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07766__A net1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput204 net204 vssd1 vssd1 vccd1 vccd1 gpio_oeb[8] sky130_fd_sc_hd__buf_2
XFILLER_0_2_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput215 net215 vssd1 vssd1 vccd1 vccd1 gpio_out[18] sky130_fd_sc_hd__buf_2
Xoutput226 net226 vssd1 vssd1 vccd1 vccd1 gpio_out[29] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_58_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput237 net237 vssd1 vssd1 vccd1 vccd1 gpio_out[9] sky130_fd_sc_hd__clkbuf_4
Xoutput248 net248 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[1] sky130_fd_sc_hd__buf_2
XANTENNA__10192__A _04565_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput259 net259 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[5] sky130_fd_sc_hd__buf_2
XANTENNA__08791__A1 net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09981__A _05852_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07961_ net613 _03900_ _03902_ vssd1 vssd1 vccd1 vccd1 _03903_ sky130_fd_sc_hd__a21o_1
XANTENNA__08791__B2 net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08218__S1 net1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11438__D net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09700_ _03866_ net589 _05641_ vssd1 vssd1 vccd1 vccd1 _05642_ sky130_fd_sc_hd__a21oi_1
X_06912_ net1200 team_03_WB.instance_to_wrap.core.register_file.registers_state\[132\]
+ vssd1 vssd1 vccd1 vccd1 _02854_ sky130_fd_sc_hd__or2_1
X_07892_ net1091 team_03_WB.instance_to_wrap.core.register_file.registers_state\[335\]
+ net1150 vssd1 vssd1 vccd1 vccd1 _03834_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_147_3393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08543__A1 net1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09631_ _03314_ _04415_ net665 _05572_ vssd1 vssd1 vccd1 vccd1 _05573_ sky130_fd_sc_hd__a22o_1
XFILLER_0_4_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06843_ net1164 vssd1 vssd1 vccd1 vccd1 _02786_ sky130_fd_sc_hd__inv_2
XANTENNA__11227__S net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07897__A3 net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09562_ _05180_ _05503_ _05178_ vssd1 vssd1 vccd1 vccd1 _05504_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_104_2507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_2518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08513_ net871 _04451_ _04454_ vssd1 vssd1 vccd1 vccd1 _04455_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_19_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09493_ net581 _05433_ _05434_ vssd1 vssd1 vccd1 vccd1 _05435_ sky130_fd_sc_hd__and3_1
XFILLER_0_136_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_19_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11173__D net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_2854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_121_2865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08444_ net541 _04384_ _04355_ vssd1 vssd1 vccd1 vccd1 _04386_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_172_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06845__A net1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_738 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_173_3921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_173_3932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12058__S net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08375_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[822\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[790\]
+ net970 vssd1 vssd1 vccd1 vccd1 _04317_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout423_A _06560_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1165_A net1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07326_ net807 _03266_ _03267_ vssd1 vssd1 vccd1 vccd1 _03268_ sky130_fd_sc_hd__or3_1
XFILLER_0_18_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_162_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07806__B1 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07379__C net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10086__B _05730_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold1273_A team_03_WB.instance_to_wrap.CPU_DAT_O\[0\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_143_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07257_ net1191 team_03_WB.instance_to_wrap.core.register_file.registers_state\[328\]
+ vssd1 vssd1 vccd1 vccd1 _03199_ sky130_fd_sc_hd__or2_1
XANTENNA__09008__C1 net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout309_X net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1332_A net1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07676__A net1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07188_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[947\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[915\]
+ net762 vssd1 vssd1 vccd1 vccd1 _03130_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout792_A net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11366__B1 net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1120_X net1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1218_X net1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1407 net1408 vssd1 vssd1 vccd1 vccd1 net1407 sky130_fd_sc_hd__buf_4
XANTENNA_fanout580_X net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout420 _06560_ vssd1 vssd1 vccd1 vccd1 net420 sky130_fd_sc_hd__buf_8
Xfanout1418 net1436 vssd1 vssd1 vccd1 vccd1 net1418 sky130_fd_sc_hd__buf_2
Xfanout431 net438 vssd1 vssd1 vccd1 vccd1 net431 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_100_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1429 net1430 vssd1 vssd1 vccd1 vccd1 net1429 sky130_fd_sc_hd__buf_2
Xfanout442 _06819_ vssd1 vssd1 vccd1 vccd1 net442 sky130_fd_sc_hd__buf_4
XANTENNA__11669__A1 net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout453 net481 vssd1 vssd1 vccd1 vccd1 net453 sky130_fd_sc_hd__clkbuf_4
Xfanout464 net472 vssd1 vssd1 vccd1 vccd1 net464 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07337__A2 net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout475 net476 vssd1 vssd1 vccd1 vccd1 net475 sky130_fd_sc_hd__clkbuf_4
Xfanout486 _06680_ vssd1 vssd1 vccd1 vccd1 net486 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_6_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09829_ _05263_ _05264_ vssd1 vssd1 vccd1 vccd1 _05771_ sky130_fd_sc_hd__xnor2_1
Xfanout497 net500 vssd1 vssd1 vccd1 vccd1 net497 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout845_X net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07888__A3 net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12840_ net1291 vssd1 vssd1 vccd1 vccd1 _00604_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_17_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12771_ net1354 vssd1 vssd1 vccd1 vccd1 _00535_ sky130_fd_sc_hd__inv_2
XANTENNA__12757__A net1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11722_ _06454_ net596 net456 _06808_ net1889 vssd1 vssd1 vccd1 vccd1 _01814_ sky130_fd_sc_hd__a32o_1
X_14510_ clknet_leaf_129_wb_clk_i _02274_ _00875_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[864\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_139_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_81_2050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09131__A net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14441_ clknet_leaf_78_wb_clk_i _02205_ _00806_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[795\]
+ sky130_fd_sc_hd__dfrtp_1
X_11653_ net2233 _06619_ net343 vssd1 vssd1 vccd1 vccd1 _01880_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_805 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10604_ net1681 team_03_WB.instance_to_wrap.CPU_DAT_O\[25\] net841 vssd1 vssd1 vccd1
+ vccd1 _02524_ sky130_fd_sc_hd__mux2_1
X_14372_ clknet_leaf_23_wb_clk_i _02136_ _00737_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[726\]
+ sky130_fd_sc_hd__dfrtp_1
X_11584_ net301 net2306 net447 vssd1 vssd1 vccd1 vccd1 _01945_ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13323_ net1315 vssd1 vssd1 vccd1 vccd1 _01087_ sky130_fd_sc_hd__inv_2
XFILLER_0_49_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_16 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13588__A net1346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10535_ net162 net1032 net1024 net1713 vssd1 vssd1 vccd1 vccd1 _02575_ sky130_fd_sc_hd__a22o_1
XFILLER_0_36_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11600__S net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13254_ net1301 vssd1 vssd1 vccd1 vccd1 _01018_ sky130_fd_sc_hd__inv_2
X_10466_ _06047_ _06049_ vssd1 vssd1 vccd1 vccd1 _06279_ sky130_fd_sc_hd__xnor2_1
X_12205_ net1520 vssd1 vssd1 vccd1 vccd1 _02348_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_122_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13185_ net1261 vssd1 vssd1 vccd1 vccd1 _00949_ sky130_fd_sc_hd__inv_2
XANTENNA__08222__B1 net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10397_ _06222_ _06223_ team_03_WB.instance_to_wrap.core.pc.current_pc\[16\] net680
+ vssd1 vssd1 vccd1 vccd1 _02650_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_0_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_36_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_3_6_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_6_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_36_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12136_ net1561 vssd1 vssd1 vccd1 vccd1 _02417_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__11109__A0 net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_1032 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12067_ _06630_ net2693 net358 vssd1 vssd1 vccd1 vccd1 _01479_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_53_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_97_wb_clk_i clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_97_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_53_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09306__A net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11018_ net490 net646 _06582_ net420 net1927 vssd1 vssd1 vccd1 vccd1 _02292_ sky130_fd_sc_hd__a32o_1
XANTENNA__08210__A net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_26_wb_clk_i clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_26_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_126_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_142_3290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11842__Y _06812_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12085__A1 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12969_ net1253 vssd1 vssd1 vccd1 vccd1 _00733_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14708_ clknet_leaf_68_wb_clk_i _02472_ _01073_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.control_logic.instruction\[5\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_157_431 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_32 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14639_ clknet_leaf_135_wb_clk_i _02403_ _01004_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[993\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_16_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08160_ net1217 _04100_ _04101_ vssd1 vssd1 vccd1 vccd1 _04102_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_27_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_98 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07111_ net1104 team_03_WB.instance_to_wrap.core.register_file.registers_state\[33\]
+ net899 vssd1 vssd1 vccd1 vccd1 _03053_ sky130_fd_sc_hd__or3_1
XFILLER_0_70_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_884 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11060__A2 net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08091_ net1172 team_03_WB.instance_to_wrap.core.register_file.registers_state\[58\]
+ net880 vssd1 vssd1 vccd1 vccd1 _04033_ sky130_fd_sc_hd__and3_1
XFILLER_0_71_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_359 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10915__A net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11510__S net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkload30 clknet_leaf_176_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload30/X sky130_fd_sc_hd__clkbuf_8
X_07042_ net1100 team_03_WB.instance_to_wrap.core.register_file.registers_state\[451\]
+ net801 team_03_WB.instance_to_wrap.core.register_file.registers_state\[483\] vssd1
+ vssd1 vccd1 vccd1 _02984_ sky130_fd_sc_hd__a22o_1
XFILLER_0_30_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload41 clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload41/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_141_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload52 clknet_leaf_172_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload52/X sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_77_1952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload63 clknet_leaf_43_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload63/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__11348__B1 net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_707 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload74 clknet_leaf_54_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload74/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_2_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_77_1963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload85 clknet_leaf_33_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload85/Y sky130_fd_sc_hd__clkinv_2
XANTENNA__07016__A1 net1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload96 clknet_leaf_65_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload96/Y sky130_fd_sc_hd__bufinv_16
XANTENNA__08213__B1 net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_149_3433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_149_3444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08993_ net1062 _04934_ vssd1 vssd1 vccd1 vccd1 _04935_ sky130_fd_sc_hd__nand2_1
XFILLER_0_167_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_166_3780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07944_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[567\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[535\]
+ net767 vssd1 vssd1 vccd1 vccd1 _03886_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_166_3791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09861__D _05659_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07875_ net1189 team_03_WB.instance_to_wrap.core.register_file.registers_state\[187\]
+ vssd1 vssd1 vccd1 vccd1 _03817_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_3_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout373_A _06813_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_162_3699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06826_ team_03_WB.instance_to_wrap.core.pc.current_pc\[26\] vssd1 vssd1 vccd1 vccd1
+ _02769_ sky130_fd_sc_hd__inv_2
X_09614_ team_03_WB.instance_to_wrap.core.decoder.inst\[29\] net1021 net535 _05553_
+ vssd1 vssd1 vccd1 vccd1 _05556_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__10874__A2 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11184__C _06527_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_167_206 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09545_ _05413_ _05417_ net560 vssd1 vssd1 vccd1 vccd1 _05487_ sky130_fd_sc_hd__mux2_1
XANTENNA__10796__S net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06846__Y _02789_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1282_A net1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11481__A net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout638_A _06458_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_174_Right_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09476_ _05416_ _05417_ net554 vssd1 vssd1 vccd1 vccd1 _05418_ sky130_fd_sc_hd__mux2_1
XANTENNA__11823__A1 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07170__S net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08427_ net1228 team_03_WB.instance_to_wrap.core.register_file.registers_state\[602\]
+ net964 team_03_WB.instance_to_wrap.core.register_file.registers_state\[634\] net920
+ vssd1 vssd1 vccd1 vccd1 _04369_ sky130_fd_sc_hd__o221a_1
XFILLER_0_163_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1070_X net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout426_X net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout805_A _02850_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1168_X net1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_659 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_771 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07958__X _03900_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08358_ net1236 team_03_WB.instance_to_wrap.core.register_file.registers_state\[86\]
+ net972 team_03_WB.instance_to_wrap.core.register_file.registers_state\[118\] net921
+ vssd1 vssd1 vccd1 vccd1 _04300_ sky130_fd_sc_hd__o221a_1
XFILLER_0_163_456 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload2 clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload2/Y sky130_fd_sc_hd__clkinv_8
XANTENNA__11587__A0 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07309_ net1116 _03249_ _03250_ net1129 vssd1 vssd1 vccd1 vccd1 _03251_ sky130_fd_sc_hd__a211o_1
XFILLER_0_145_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08289_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[951\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[919\]
+ net963 vssd1 vssd1 vccd1 vccd1 _04231_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout1335_X net1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10320_ team_03_WB.instance_to_wrap.core.pc.current_pc\[30\] net678 _06157_ _06160_
+ vssd1 vssd1 vccd1 vccd1 _02664_ sky130_fd_sc_hd__o22a_1
XFILLER_0_81_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout795_X net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10251_ _06091_ _06092_ vssd1 vssd1 vccd1 vccd1 _06093_ sky130_fd_sc_hd__and2_1
XANTENNA__12000__A1 net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11359__C net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10011__A0 _03023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08755__A1 net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07102__S1 net1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10182_ team_03_WB.instance_to_wrap.core.decoder.inst\[28\] net826 _06023_ vssd1
+ vssd1 vccd1 vccd1 _06024_ sky130_fd_sc_hd__and3_1
XANTENNA__10831__Y _06434_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout962_X net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10562__B2 _05872_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1204 net1205 vssd1 vssd1 vccd1 vccd1 net1204 sky130_fd_sc_hd__buf_2
Xfanout1215 net1216 vssd1 vssd1 vccd1 vccd1 net1215 sky130_fd_sc_hd__buf_2
Xfanout1226 net1227 vssd1 vssd1 vccd1 vccd1 net1226 sky130_fd_sc_hd__clkbuf_4
Xfanout1237 net1238 vssd1 vssd1 vccd1 vccd1 net1237 sky130_fd_sc_hd__buf_2
X_14990_ clknet_leaf_64_wb_clk_i net38 _01355_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[9\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1248 net1250 vssd1 vssd1 vccd1 vccd1 net1248 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_79_1048 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1259 net1263 vssd1 vssd1 vccd1 vccd1 net1259 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_31_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11375__B net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout272 _06483_ vssd1 vssd1 vccd1 vccd1 net272 sky130_fd_sc_hd__buf_2
Xfanout283 net284 vssd1 vssd1 vccd1 vccd1 net283 sky130_fd_sc_hd__clkbuf_4
X_13941_ clknet_leaf_126_wb_clk_i _01705_ _00306_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[295\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout294 _05859_ vssd1 vssd1 vccd1 vccd1 net294 sky130_fd_sc_hd__buf_4
XANTENNA__11511__A0 _06628_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09180__A1 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13872_ clknet_leaf_158_wb_clk_i _01636_ _00237_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[226\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12823_ net1390 vssd1 vssd1 vccd1 vccd1 _00587_ sky130_fd_sc_hd__inv_2
XANTENNA__09468__C1 net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12487__A net1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11391__A net1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_141_Right_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12754_ net1396 vssd1 vssd1 vccd1 vccd1 _00518_ sky130_fd_sc_hd__inv_2
XANTENNA__09483__A2 _04503_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11705_ _06747_ net384 net340 net1916 vssd1 vssd1 vccd1 vccd1 _01829_ sky130_fd_sc_hd__a22o_1
XANTENNA__11290__A2 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12685_ net1311 vssd1 vssd1 vccd1 vccd1 _00449_ sky130_fd_sc_hd__inv_2
XFILLER_0_139_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_144_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_144_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_input91_X net91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14424_ clknet_leaf_3_wb_clk_i _02188_ _00789_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[778\]
+ sky130_fd_sc_hd__dfrtp_1
X_11636_ _06710_ net384 net348 net2463 vssd1 vssd1 vccd1 vccd1 _01896_ sky130_fd_sc_hd__a22o_1
XFILLER_0_65_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_170_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11578__A0 _06413_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08038__A3 net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08669__S1 net1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_730 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_170_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10294__X _06136_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11042__A2 net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14355_ clknet_leaf_102_wb_clk_i _02119_ _00720_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[709\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11567_ net638 net705 net268 net697 vssd1 vssd1 vccd1 vccd1 _06797_ sky130_fd_sc_hd__and4_1
XANTENNA__11330__S net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10518_ net149 net1032 net1024 net1670 vssd1 vssd1 vccd1 vccd1 _02592_ sky130_fd_sc_hd__a22o_1
X_13306_ net1314 vssd1 vssd1 vccd1 vccd1 _01070_ sky130_fd_sc_hd__inv_2
Xhold709 team_03_WB.instance_to_wrap.core.register_file.registers_state\[702\] vssd1
+ vssd1 vccd1 vccd1 net2202 sky130_fd_sc_hd__dlygate4sd3_1
X_14286_ clknet_leaf_127_wb_clk_i _02050_ _00651_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[640\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07747__C net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11498_ _06619_ net2275 net389 vssd1 vssd1 vccd1 vccd1 _02008_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13237_ net1276 vssd1 vssd1 vccd1 vccd1 _01001_ sky130_fd_sc_hd__inv_2
X_10449_ team_03_WB.instance_to_wrap.core.pc.current_pc\[6\] _06265_ net683 vssd1
+ vssd1 vccd1 vccd1 _02640_ sky130_fd_sc_hd__mux2_1
XANTENNA__12950__A net1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11269__C net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08746__A1 net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13168_ net1412 vssd1 vssd1 vccd1 vccd1 _00932_ sky130_fd_sc_hd__inv_2
XFILLER_0_23_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11750__B1 net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12119_ net238 net99 net101 vssd1 vssd1 vccd1 vccd1 _00010_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_72_1860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13099_ net1288 vssd1 vssd1 vccd1 vccd1 _00863_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_144_3330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_3341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11285__B _06527_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07660_ _03601_ vssd1 vssd1 vccd1 vccd1 _03602_ sky130_fd_sc_hd__inv_2
XFILLER_0_79_318 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_140_3249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06947__X _02889_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_172_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07591_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[153\] net787
+ net736 _03532_ vssd1 vssd1 vccd1 vccd1 _03533_ sky130_fd_sc_hd__a211o_1
XFILLER_0_149_228 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09330_ _04646_ _05229_ vssd1 vssd1 vccd1 vccd1 _05272_ sky130_fd_sc_hd__or2_1
XANTENNA__11505__S net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_46_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_87_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09261_ _05201_ _05202_ vssd1 vssd1 vccd1 vccd1 _05203_ sky130_fd_sc_hd__and2_1
XFILLER_0_8_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09202__C net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08212_ _04152_ _04153_ net860 vssd1 vssd1 vccd1 vccd1 _04154_ sky130_fd_sc_hd__a21o_1
XFILLER_0_172_220 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_968 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09192_ _05130_ _05133_ net556 vssd1 vssd1 vccd1 vccd1 _05134_ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08814__S net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11569__B1 net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_106 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10067__D net1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08143_ _02800_ _02802_ _02811_ _02813_ net1237 vssd1 vssd1 vccd1 vccd1 _04085_ sky130_fd_sc_hd__o221a_4
XANTENNA__07237__A1 net1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_116_2753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_2764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload130 clknet_leaf_144_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload130/X sky130_fd_sc_hd__clkbuf_8
X_08074_ net743 _04012_ _04013_ _04014_ _04015_ vssd1 vssd1 vccd1 vccd1 _04016_ sky130_fd_sc_hd__o32a_1
Xclkload141 clknet_leaf_75_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload141/X sky130_fd_sc_hd__clkbuf_4
Xclkload152 clknet_leaf_82_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload152/Y sky130_fd_sc_hd__clkinv_2
XFILLER_0_31_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload163 clknet_leaf_107_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload163/Y sky130_fd_sc_hd__clkinv_2
XTAP_TAPCELL_ROW_168_3820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07025_ net1099 team_03_WB.instance_to_wrap.core.register_file.registers_state\[579\]
+ vssd1 vssd1 vccd1 vccd1 _02967_ sky130_fd_sc_hd__and2_1
XFILLER_0_12_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload174 clknet_leaf_90_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload174/Y sky130_fd_sc_hd__inv_6
XTAP_TAPCELL_ROW_168_3831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1030_A net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08198__C1 net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08737__A1 net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1128_A net1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_8_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout490_A net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07945__C1 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_164_3739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12071__S net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold14 team_03_WB.instance_to_wrap.core.register_file.registers_state\[976\] vssd1
+ vssd1 vccd1 vccd1 net1507 sky130_fd_sc_hd__dlygate4sd3_1
X_08976_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[1001\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[969\]
+ net991 vssd1 vssd1 vccd1 vccd1 _04918_ sky130_fd_sc_hd__mux2_1
Xhold25 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1016\] vssd1
+ vssd1 vccd1 vccd1 net1518 sky130_fd_sc_hd__dlygate4sd3_1
Xhold36 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1019\] vssd1
+ vssd1 vccd1 vccd1 net1529 sky130_fd_sc_hd__dlygate4sd3_1
Xhold47 team_03_WB.instance_to_wrap.core.register_file.registers_state\[17\] vssd1
+ vssd1 vccd1 vccd1 net1540 sky130_fd_sc_hd__dlygate4sd3_1
Xhold58 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[14\] vssd1 vssd1 vccd1
+ vccd1 net1551 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07392__C net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07927_ net1087 net892 team_03_WB.instance_to_wrap.core.register_file.registers_state\[151\]
+ vssd1 vssd1 vccd1 vccd1 _03869_ sky130_fd_sc_hd__o21a_1
XANTENNA_clkbuf_leaf_85_wb_clk_i_A clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold69 team_03_WB.instance_to_wrap.ADR_I\[7\] vssd1 vssd1 vccd1 vccd1 net1562 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout376_X net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07858_ net1158 _03798_ _03799_ net823 vssd1 vssd1 vccd1 vccd1 _03800_ sky130_fd_sc_hd__o31a_1
XANTENNA__09701__A3 _05126_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout543_X net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07789_ _03729_ _03730_ vssd1 vssd1 vccd1 vccd1 _03731_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout922_A net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06920__B1 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08348__S0 net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11415__S net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09528_ _05348_ _05352_ net560 vssd1 vssd1 vccd1 vccd1 _05470_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_749 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09459_ net544 _04712_ _05132_ vssd1 vssd1 vccd1 vccd1 _05401_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_136_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07476__A1 net1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout710_X net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_148_272 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11272__A2 net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08673__B1 net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11361__D net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout808_X net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10480__B1 net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12470_ net1258 vssd1 vssd1 vccd1 vccd1 _00234_ sky130_fd_sc_hd__inv_2
XFILLER_0_164_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08724__S net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_938 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07228__A1 _03169_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11421_ net2397 net396 _06754_ net505 vssd1 vssd1 vccd1 vccd1 _02061_ sky130_fd_sc_hd__a22o_1
XFILLER_0_62_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10232__B1 _03864_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14140_ clknet_leaf_146_wb_clk_i _01904_ _00505_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[494\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_50_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11352_ net498 net626 _06728_ net401 net1955 vssd1 vssd1 vccd1 vccd1 _02104_ sky130_fd_sc_hd__a32o_1
XFILLER_0_132_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_342 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07567__C net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10783__A1 net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11980__A0 _06426_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10303_ team_03_WB.instance_to_wrap.core.pc.current_pc\[19\] team_03_WB.instance_to_wrap.core.pc.current_pc\[18\]
+ _06144_ vssd1 vssd1 vccd1 vccd1 _06145_ sky130_fd_sc_hd__and3_1
XFILLER_0_120_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14071_ clknet_leaf_112_wb_clk_i _01835_ _00436_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[425\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_132_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11283_ net715 _06523_ net831 vssd1 vssd1 vccd1 vccd1 _06709_ sky130_fd_sc_hd__and3_1
XFILLER_0_21_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12770__A net1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08728__A1 net1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13022_ net1410 vssd1 vssd1 vccd1 vccd1 _00786_ sky130_fd_sc_hd__inv_2
XANTENNA_input51_A gpio_in[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10234_ _06073_ _06074_ vssd1 vssd1 vccd1 vccd1 _06076_ sky130_fd_sc_hd__nor2_1
XFILLER_0_30_671 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1001 net1003 vssd1 vssd1 vccd1 vccd1 net1001 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07936__C1 net1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1012 net1013 vssd1 vssd1 vccd1 vccd1 net1012 sky130_fd_sc_hd__clkbuf_2
X_10165_ _03724_ _06005_ vssd1 vssd1 vccd1 vccd1 _06007_ sky130_fd_sc_hd__nor2_1
Xfanout1023 net1024 vssd1 vssd1 vccd1 vccd1 net1023 sky130_fd_sc_hd__clkbuf_4
Xfanout1034 net1035 vssd1 vssd1 vccd1 vccd1 net1034 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_50_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1045 net1046 vssd1 vssd1 vccd1 vccd1 net1045 sky130_fd_sc_hd__clkbuf_4
Xfanout1056 net1058 vssd1 vssd1 vccd1 vccd1 net1056 sky130_fd_sc_hd__buf_2
X_14973_ clknet_leaf_92_wb_clk_i _02725_ _01338_ vssd1 vssd1 vccd1 vccd1 net225 sky130_fd_sc_hd__dfrtp_1
X_10096_ net312 _05429_ _05936_ _05939_ vssd1 vssd1 vccd1 vccd1 _05940_ sky130_fd_sc_hd__or4_1
Xfanout1067 net1069 vssd1 vssd1 vccd1 vccd1 net1067 sky130_fd_sc_hd__buf_4
Xfanout1078 net1079 vssd1 vssd1 vccd1 vccd1 net1078 sky130_fd_sc_hd__buf_4
Xfanout1089 net1093 vssd1 vssd1 vccd1 vccd1 net1089 sky130_fd_sc_hd__buf_2
XANTENNA_output138_A net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_1046 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10838__A2 net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13924_ clknet_leaf_36_wb_clk_i _01688_ _00289_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[278\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08900__A1 net1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13855_ clknet_leaf_20_wb_clk_i _01619_ _00220_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[209\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_159_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06927__B net1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11325__S net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13106__A net1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_204 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12806_ net1300 vssd1 vssd1 vccd1 vccd1 _00570_ sky130_fd_sc_hd__inv_2
XANTENNA__09456__A2 _04080_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10998_ net2263 net423 _06571_ net512 vssd1 vssd1 vccd1 vccd1 _02301_ sky130_fd_sc_hd__a22o_1
X_13786_ clknet_leaf_142_wb_clk_i _01550_ _00151_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[140\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_48_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08113__C1 net1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07467__A1 net1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12737_ net1282 vssd1 vssd1 vccd1 vccd1 _00501_ sky130_fd_sc_hd__inv_2
XFILLER_0_139_283 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12668_ net1414 vssd1 vssd1 vccd1 vccd1 _00432_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09957__C net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07219__A1 net1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14407_ clknet_leaf_108_wb_clk_i _02171_ _00772_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[761\]
+ sky130_fd_sc_hd__dfrtp_1
X_11619_ _06693_ net381 net347 net2180 vssd1 vssd1 vccd1 vccd1 _01913_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_96_2347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09759__A3 _04922_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12599_ net1392 vssd1 vssd1 vccd1 vccd1 _00363_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_96_2358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08967__A1 net1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11566__A3 _06675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14338_ clknet_leaf_173_wb_clk_i _02102_ _00703_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[692\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_638 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold506 team_03_WB.instance_to_wrap.core.register_file.registers_state\[422\] vssd1
+ vssd1 vccd1 vccd1 net1999 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_133_3097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold517 team_03_WB.instance_to_wrap.core.register_file.registers_state\[276\] vssd1
+ vssd1 vccd1 vccd1 net2010 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11971__B1 net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_74_1900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold528 team_03_WB.instance_to_wrap.core.register_file.registers_state\[245\] vssd1
+ vssd1 vccd1 vccd1 net2021 sky130_fd_sc_hd__dlygate4sd3_1
Xhold539 team_03_WB.instance_to_wrap.core.register_file.registers_state\[312\] vssd1
+ vssd1 vccd1 vccd1 net2032 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12680__A net1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14269_ clknet_leaf_25_wb_clk_i _02033_ _00634_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[623\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09067__S1 net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09465__S net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_111_2650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_41_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_41_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__10912__B net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_2661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_70_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11723__B1 _06808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08830_ net434 net429 _04770_ net551 vssd1 vssd1 vccd1 vccd1 _04772_ sky130_fd_sc_hd__o31a_1
Xhold1206 team_03_WB.instance_to_wrap.core.register_file.registers_state\[65\] vssd1
+ vssd1 vccd1 vccd1 net2699 sky130_fd_sc_hd__dlygate4sd3_1
X_08761_ net1052 team_03_WB.instance_to_wrap.core.register_file.registers_state\[963\]
+ net1004 team_03_WB.instance_to_wrap.core.register_file.registers_state\[995\] net1065
+ vssd1 vssd1 vccd1 vccd1 _04703_ sky130_fd_sc_hd__a221o_1
Xhold1217 team_03_WB.instance_to_wrap.core.register_file.registers_state\[603\] vssd1
+ vssd1 vccd1 vccd1 net2710 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1228 team_03_WB.instance_to_wrap.core.register_file.registers_state\[595\] vssd1
+ vssd1 vccd1 vccd1 net2721 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_174_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1239 team_03_WB.instance_to_wrap.core.register_file.registers_state\[211\] vssd1
+ vssd1 vccd1 vccd1 net2732 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_174_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09144__A1 net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11446__D net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07712_ _03652_ _03653_ net1165 vssd1 vssd1 vccd1 vccd1 _03654_ sky130_fd_sc_hd__o21a_1
XFILLER_0_100_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10829__A2 net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08692_ net1241 team_03_WB.instance_to_wrap.core.register_file.registers_state\[168\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[136\] net976 net924
+ vssd1 vssd1 vccd1 vccd1 _04634_ sky130_fd_sc_hd__a221o_1
XANTENNA__07155__B1 _02870_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_2_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_07643_ net824 _03584_ vssd1 vssd1 vccd1 vccd1 _03585_ sky130_fd_sc_hd__nand2_1
XANTENNA__11743__B net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07052__A1_N net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15049__1490 vssd1 vssd1 vccd1 vccd1 net1490 _15049__1490/LO sky130_fd_sc_hd__conb_1
XFILLER_0_79_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_169_wb_clk_i_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_95_619 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07574_ net1189 team_03_WB.instance_to_wrap.core.register_file.registers_state\[856\]
+ vssd1 vssd1 vccd1 vccd1 _03516_ sky130_fd_sc_hd__or2_1
XFILLER_0_48_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09313_ net578 _05254_ vssd1 vssd1 vccd1 vccd1 _05255_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07458__A1 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08655__B1 net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11254__A2 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout336_A net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09244_ _04119_ _05184_ vssd1 vssd1 vccd1 vccd1 _05186_ sky130_fd_sc_hd__nand2_1
XFILLER_0_111_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1078_A net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_157_3598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_2804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09175_ _05115_ _05116_ vssd1 vssd1 vccd1 vccd1 _05117_ sky130_fd_sc_hd__nor2_1
XANTENNA__12066__S net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout503_A net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1245_A net1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08126_ net1146 _04057_ _04067_ vssd1 vssd1 vccd1 vccd1 _04068_ sky130_fd_sc_hd__o21ai_1
XANTENNA__08958__A1 net1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09080__B1 net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10765__A1 _05082_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11962__B1 net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_1_Right_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07630__A1 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08057_ _03995_ _03998_ net822 vssd1 vssd1 vccd1 vccd1 _03999_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout1412_A net1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07008_ _02949_ _02947_ vssd1 vssd1 vccd1 vccd1 _02950_ sky130_fd_sc_hd__and2b_1
XANTENNA_fanout493_X net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout872_A net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1200_X net1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout660_X net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08959_ net856 _04899_ _04900_ vssd1 vssd1 vccd1 vccd1 _04901_ sky130_fd_sc_hd__or3_1
XANTENNA_fanout758_X net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11970_ net638 _06747_ net468 net365 net2052 vssd1 vssd1 vccd1 vccd1 _01573_ sky130_fd_sc_hd__a32o_1
XANTENNA__09686__A2 _04178_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08343__C1 net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_16_Left_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_168_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10921_ net270 net2240 net518 vssd1 vssd1 vccd1 vccd1 _02316_ sky130_fd_sc_hd__mux2_1
XANTENNA__07850__C net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout925_X net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_811 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13640_ net1404 vssd1 vssd1 vccd1 vccd1 _01404_ sky130_fd_sc_hd__inv_2
XFILLER_0_169_879 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10852_ team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[20\] net307 net685 vssd1
+ vssd1 vccd1 vccd1 _06451_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_67_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07449__A1 _03390_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13571_ net1428 vssd1 vssd1 vccd1 vccd1 _01335_ sky130_fd_sc_hd__inv_2
X_10783_ net613 _05918_ _06385_ _06293_ vssd1 vssd1 vccd1 vccd1 _06393_ sky130_fd_sc_hd__a31o_1
XANTENNA__08646__B1 net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08110__A2 net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07859__A net1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12522_ net1288 vssd1 vssd1 vccd1 vccd1 _00286_ sky130_fd_sc_hd__inv_2
XFILLER_0_164_551 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_23_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_23_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input99_A wbs_cyc_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_151_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12453_ net1353 vssd1 vssd1 vccd1 vccd1 _00217_ sky130_fd_sc_hd__inv_2
XFILLER_0_152_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11404_ net278 net2667 net397 vssd1 vssd1 vccd1 vccd1 _02076_ sky130_fd_sc_hd__mux2_1
X_12384_ net1400 vssd1 vssd1 vccd1 vccd1 _00148_ sky130_fd_sc_hd__inv_2
XANTENNA__08413__A3 _04354_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11953__B1 net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11335_ net280 net709 net695 vssd1 vssd1 vccd1 vccd1 _06720_ sky130_fd_sc_hd__and3_1
X_14123_ clknet_leaf_40_wb_clk_i _01887_ _00488_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[477\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_162_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_91_2244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_2255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11266_ net514 net642 _06700_ net411 net2204 vssd1 vssd1 vccd1 vccd1 _02162_ sky130_fd_sc_hd__a32o_1
X_14054_ clknet_leaf_28_wb_clk_i _01818_ _00419_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[408\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08042__X _03984_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11705__B1 net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10217_ _06024_ _06058_ vssd1 vssd1 vccd1 vccd1 _06059_ sky130_fd_sc_hd__nor2_1
X_13005_ net1332 vssd1 vssd1 vccd1 vccd1 _00769_ sky130_fd_sc_hd__inv_2
X_11197_ net2244 net414 _06679_ net514 vssd1 vssd1 vccd1 vccd1 _02210_ sky130_fd_sc_hd__a22o_1
XFILLER_0_94_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07385__B1 net1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08582__C1 net1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07924__A2 _03864_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10148_ _04207_ net672 _05989_ vssd1 vssd1 vccd1 vccd1 _05990_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_94_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09126__A1 net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14956_ clknet_leaf_92_wb_clk_i _02708_ _01321_ vssd1 vssd1 vccd1 vccd1 net208 sky130_fd_sc_hd__dfrtp_1
X_10079_ _05921_ _05922_ net314 _05920_ vssd1 vssd1 vccd1 vccd1 _05923_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_89_2195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07137__B1 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09677__A2 _04119_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09314__A _04711_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11563__B net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07688__A1 net1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13907_ clknet_leaf_106_wb_clk_i _01671_ _00272_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[261\]
+ sky130_fd_sc_hd__dfrtp_1
X_14887_ clknet_leaf_65_wb_clk_i _02650_ _01252_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.pc.current_pc\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13838_ clknet_leaf_131_wb_clk_i _01602_ _00203_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[192\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_134_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_378 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11236__A2 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10894__S net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13769_ clknet_leaf_116_wb_clk_i _01533_ _00134_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[123\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10444__B1 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_21_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07290_ net808 _03230_ _03231_ vssd1 vssd1 vccd1 vccd1 _03232_ sky130_fd_sc_hd__or3_1
XFILLER_0_128_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10995__A1 net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08591__C _04532_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07121__X _03063_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_3148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10907__B net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_142_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07488__B _02819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_908 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_152_3495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_2701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_576 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10747__A1 _05718_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_295 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11944__B1 net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold303 team_03_WB.instance_to_wrap.core.register_file.registers_state\[11\] vssd1
+ vssd1 vccd1 vccd1 net1796 sky130_fd_sc_hd__dlygate4sd3_1
Xhold314 team_03_WB.instance_to_wrap.core.register_file.registers_state\[392\] vssd1
+ vssd1 vccd1 vccd1 net1807 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold325 team_03_WB.instance_to_wrap.CPU_DAT_I\[0\] vssd1 vssd1 vccd1 vccd1 net1818
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_159_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09600__A_N _05541_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold336 _02519_ vssd1 vssd1 vccd1 vccd1 net1829 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold347 team_03_WB.instance_to_wrap.core.register_file.registers_state\[66\] vssd1
+ vssd1 vccd1 vccd1 net1840 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold358 team_03_WB.instance_to_wrap.core.register_file.registers_state\[290\] vssd1
+ vssd1 vccd1 vccd1 net1851 sky130_fd_sc_hd__dlygate4sd3_1
Xhold369 net230 vssd1 vssd1 vccd1 vccd1 net1862 sky130_fd_sc_hd__dlygate4sd3_1
X_09931_ _03312_ net663 vssd1 vssd1 vccd1 vccd1 _05870_ sky130_fd_sc_hd__nor2_1
XFILLER_0_1_874 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout805 _02850_ vssd1 vssd1 vccd1 vccd1 net805 sky130_fd_sc_hd__buf_4
Xfanout816 _02848_ vssd1 vssd1 vccd1 vccd1 net816 sky130_fd_sc_hd__buf_4
X_09862_ _05278_ _05281_ _05300_ vssd1 vssd1 vccd1 vccd1 _05804_ sky130_fd_sc_hd__nand3_1
Xfanout827 net828 vssd1 vssd1 vccd1 vccd1 net827 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_110_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout838 net839 vssd1 vssd1 vccd1 vccd1 net838 sky130_fd_sc_hd__buf_4
Xfanout849 _04097_ vssd1 vssd1 vccd1 vccd1 net849 sky130_fd_sc_hd__buf_8
XANTENNA__07376__B1 net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11172__B2 net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07009__A net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08813_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[929\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[897\]
+ net980 vssd1 vssd1 vccd1 vccd1 _04755_ sky130_fd_sc_hd__mux2_1
Xhold1003 team_03_WB.instance_to_wrap.core.register_file.registers_state\[518\] vssd1
+ vssd1 vccd1 vccd1 net2496 sky130_fd_sc_hd__dlygate4sd3_1
X_09793_ _05421_ _05734_ net573 vssd1 vssd1 vccd1 vccd1 _05735_ sky130_fd_sc_hd__mux2_2
Xhold1014 team_03_WB.instance_to_wrap.core.register_file.registers_state\[617\] vssd1
+ vssd1 vccd1 vccd1 net2507 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1025 team_03_WB.instance_to_wrap.core.register_file.registers_state\[491\] vssd1
+ vssd1 vccd1 vccd1 net2518 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1036 team_03_WB.instance_to_wrap.core.register_file.registers_state\[924\] vssd1
+ vssd1 vccd1 vccd1 net2529 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1047 team_03_WB.instance_to_wrap.core.register_file.registers_state\[780\] vssd1
+ vssd1 vccd1 vccd1 net2540 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1058 team_03_WB.instance_to_wrap.core.register_file.registers_state\[723\] vssd1
+ vssd1 vccd1 vccd1 net2551 sky130_fd_sc_hd__dlygate4sd3_1
X_08744_ net1052 team_03_WB.instance_to_wrap.core.register_file.registers_state\[195\]
+ net1004 team_03_WB.instance_to_wrap.core.register_file.registers_state\[227\] net926
+ vssd1 vssd1 vccd1 vccd1 _04686_ sky130_fd_sc_hd__a221o_1
XFILLER_0_139_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07128__B1 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06848__A net1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1069 team_03_WB.instance_to_wrap.core.register_file.registers_state\[480\] vssd1
+ vssd1 vccd1 vccd1 net2562 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07679__A1 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08675_ _04615_ _04616_ vssd1 vssd1 vccd1 vccd1 _04617_ sky130_fd_sc_hd__and2_1
XFILLER_0_36_1024 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout453_A net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1195_A net1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10683__B1 net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_159_3638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07626_ net1094 team_03_WB.instance_to_wrap.core.register_file.registers_state\[46\]
+ net896 vssd1 vssd1 vccd1 vccd1 _03568_ sky130_fd_sc_hd__or3_1
XANTENNA__11192__C _06545_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_159_3649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09511__X _05453_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08628__B1 net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07557_ net806 _03497_ _03498_ vssd1 vssd1 vccd1 vccd1 _03499_ sky130_fd_sc_hd__or3_1
XANTENNA_fanout620_A net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12585__A net1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1362_A net1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout339_X net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout718_A net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_376 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07488_ team_03_WB.instance_to_wrap.core.decoder.inst\[27\] _02819_ vssd1 vssd1 vccd1
+ vccd1 _03430_ sky130_fd_sc_hd__and2_2
XFILLER_0_118_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08127__X _04069_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09227_ _03280_ _05168_ vssd1 vssd1 vccd1 vccd1 _05169_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_146_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1150_X net1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07851__A1 net1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout506_X net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1248_X net1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09158_ net569 _05099_ vssd1 vssd1 vccd1 vccd1 _05100_ sky130_fd_sc_hd__and2_1
XANTENNA__10738__A1 _05697_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11488__X _06778_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08109_ net728 _04048_ _04049_ net1114 vssd1 vssd1 vccd1 vccd1 _04051_ sky130_fd_sc_hd__a31o_1
XANTENNA__07603__A1 net1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08800__B1 net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09089_ net1055 team_03_WB.instance_to_wrap.core.register_file.registers_state\[653\]
+ net1003 team_03_WB.instance_to_wrap.core.register_file.registers_state\[685\] net925
+ vssd1 vssd1 vccd1 vccd1 _05031_ sky130_fd_sc_hd__a221o_1
X_11120_ net1042 net696 vssd1 vssd1 vccd1 vccd1 _06634_ sky130_fd_sc_hd__nand2_1
XFILLER_0_130_963 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11950__A3 net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold870 team_03_WB.instance_to_wrap.core.register_file.registers_state\[766\] vssd1
+ vssd1 vccd1 vccd1 net2363 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout875_X net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold881 team_03_WB.instance_to_wrap.core.register_file.registers_state\[848\] vssd1
+ vssd1 vccd1 vccd1 net2374 sky130_fd_sc_hd__dlygate4sd3_1
X_11051_ net707 net269 net830 vssd1 vssd1 vccd1 vccd1 _06603_ sky130_fd_sc_hd__and3_1
Xhold892 team_03_WB.instance_to_wrap.core.register_file.registers_state\[455\] vssd1
+ vssd1 vccd1 vccd1 net2385 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11367__C net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11163__A1 net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10002_ _05887_ net2497 net288 vssd1 vssd1 vccd1 vccd1 _02712_ sky130_fd_sc_hd__mux2_1
XANTENNA__07906__A2 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07462__S0 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10979__S net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09108__A1 net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_700 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14810_ clknet_leaf_104_wb_clk_i net1601 _01175_ vssd1 vssd1 vccd1 vccd1 net161 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_157_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08316__C1 net1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09134__A net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14741_ clknet_leaf_62_wb_clk_i _02505_ _01106_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11383__B _06527_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input14_A DAT_I[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07580__C net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11953_ net624 _06730_ net455 net363 net1878 vssd1 vssd1 vccd1 vccd1 _01590_ sky130_fd_sc_hd__a32o_1
XFILLER_0_87_939 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10904_ net298 net2715 net520 vssd1 vssd1 vccd1 vccd1 _02319_ sky130_fd_sc_hd__mux2_1
X_14672_ clknet_leaf_86_wb_clk_i _02436_ _01037_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.ADR_I\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11884_ net626 _06693_ net460 net372 net1976 vssd1 vssd1 vccd1 vccd1 _01657_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_84_2092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13623_ net1434 vssd1 vssd1 vccd1 vccd1 _01387_ sky130_fd_sc_hd__inv_2
XFILLER_0_67_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10835_ team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[23\] _05865_ net318 _06403_
+ net687 vssd1 vssd1 vccd1 vccd1 _06437_ sky130_fd_sc_hd__a41o_1
XFILLER_0_168_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11603__S net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13554_ net1427 vssd1 vssd1 vccd1 vccd1 _01318_ sky130_fd_sc_hd__inv_2
XFILLER_0_39_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_871 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10766_ net1552 net530 net525 _06377_ vssd1 vssd1 vccd1 vccd1 _02435_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_41_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09831__A2 _04711_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12505_ net1365 vssd1 vssd1 vccd1 vccd1 _00269_ sky130_fd_sc_hd__inv_2
XANTENNA__07842__A1 net1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10697_ _06317_ _06333_ _06335_ net606 vssd1 vssd1 vccd1 vccd1 _06336_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_164_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13485_ net1345 vssd1 vssd1 vccd1 vccd1 _01249_ sky130_fd_sc_hd__inv_2
X_12436_ net1310 vssd1 vssd1 vccd1 vccd1 _00200_ sky130_fd_sc_hd__inv_2
XANTENNA__11926__A0 _06624_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11398__X _06752_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_3045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07055__C1 net1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12367_ net1336 vssd1 vssd1 vccd1 vccd1 _00131_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14106_ clknet_leaf_144_wb_clk_i _01870_ _00471_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[460\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07528__S net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09309__A net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11318_ _06625_ net2706 net406 vssd1 vssd1 vccd1 vccd1 _02127_ sky130_fd_sc_hd__mux2_1
X_15086_ net1472 vssd1 vssd1 vccd1 vccd1 la_data_out[22] sky130_fd_sc_hd__buf_2
X_12298_ net1279 vssd1 vssd1 vccd1 vccd1 _00062_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_39_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14037_ clknet_leaf_126_wb_clk_i _01801_ _00402_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[391\]
+ sky130_fd_sc_hd__dfrtp_1
X_11249_ net276 net716 net828 vssd1 vssd1 vccd1 vccd1 _06692_ sky130_fd_sc_hd__and3_1
XFILLER_0_38_44 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10889__S net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10901__A1 net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12103__B1 net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11293__B net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_43 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14939_ clknet_leaf_52_wb_clk_i _02694_ _01304_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_O\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11457__A2 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_2560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08460_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[60\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[28\]
+ net953 vssd1 vssd1 vccd1 vccd1 _04402_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_65_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07411_ net1084 team_03_WB.instance_to_wrap.core.register_file.registers_state\[628\]
+ net889 vssd1 vssd1 vccd1 vccd1 _03353_ sky130_fd_sc_hd__or3_1
XFILLER_0_86_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08391_ net856 _04331_ _04332_ vssd1 vssd1 vccd1 vccd1 _04333_ sky130_fd_sc_hd__or3_1
XANTENNA__09807__C1 net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_2468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_102_2479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11513__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07342_ net1172 team_03_WB.instance_to_wrap.core.register_file.registers_state\[188\]
+ net888 net1123 vssd1 vssd1 vccd1 vccd1 _03284_ sky130_fd_sc_hd__a211o_1
XFILLER_0_174_156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_173 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08086__A1 net1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_154_3535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_154_3546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10968__A1 team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[1\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11090__A0 _06479_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07273_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[937\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[905\]
+ net788 vssd1 vssd1 vccd1 vccd1 _03215_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09012_ _04953_ vssd1 vssd1 vccd1 vccd1 _04954_ sky130_fd_sc_hd__inv_2
XFILLER_0_116_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_171_3882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_171_3893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold100 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1012\] vssd1
+ vssd1 vccd1 vccd1 net1593 sky130_fd_sc_hd__dlygate4sd3_1
Xhold111 team_03_WB.instance_to_wrap.core.register_file.registers_state\[961\] vssd1
+ vssd1 vccd1 vccd1 net1604 sky130_fd_sc_hd__dlygate4sd3_1
Xhold122 _02572_ vssd1 vssd1 vccd1 vccd1 net1615 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_70 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold133 team_03_WB.instance_to_wrap.core.register_file.registers_state\[28\] vssd1
+ vssd1 vccd1 vccd1 net1626 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08794__C1 net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold144 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1015\] vssd1
+ vssd1 vccd1 vccd1 net1637 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09219__A net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold155 net120 vssd1 vssd1 vccd1 vccd1 net1648 sky130_fd_sc_hd__dlygate4sd3_1
Xhold166 _02617_ vssd1 vssd1 vccd1 vccd1 net1659 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08123__A net1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold177 team_03_WB.instance_to_wrap.CPU_DAT_I\[21\] vssd1 vssd1 vccd1 vccd1 net1670
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold188 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[25\] vssd1 vssd1 vccd1
+ vccd1 net1681 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout602 net603 vssd1 vssd1 vccd1 vccd1 net602 sky130_fd_sc_hd__buf_2
X_09914_ _05659_ _05822_ _05855_ vssd1 vssd1 vccd1 vccd1 _05856_ sky130_fd_sc_hd__and3_1
Xhold199 net201 vssd1 vssd1 vccd1 vccd1 net1692 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout613 net616 vssd1 vssd1 vccd1 vccd1 net613 sky130_fd_sc_hd__buf_4
XFILLER_0_10_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout624 net625 vssd1 vssd1 vccd1 vccd1 net624 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout1110_A net1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10091__C _05821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout635 net638 vssd1 vssd1 vccd1 vccd1 net635 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11145__B2 net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1208_A net1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08546__C1 net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout646 net647 vssd1 vssd1 vccd1 vccd1 net646 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08010__A1 net1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input6_A DAT_I[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09845_ net570 net592 vssd1 vssd1 vccd1 vccd1 _05787_ sky130_fd_sc_hd__or2_1
Xfanout657 net658 vssd1 vssd1 vccd1 vccd1 net657 sky130_fd_sc_hd__buf_4
XFILLER_0_77_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout570_A net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11696__A2 net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout668 _06564_ vssd1 vssd1 vccd1 vccd1 net668 sky130_fd_sc_hd__clkbuf_4
Xfanout679 net681 vssd1 vssd1 vccd1 vccd1 net679 sky130_fd_sc_hd__buf_2
XANTENNA_fanout289_X net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11484__A net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout668_A _06564_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07364__A3 net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09776_ _05709_ _05712_ _05717_ vssd1 vssd1 vccd1 vccd1 _05718_ sky130_fd_sc_hd__or3_4
XANTENNA__08269__S net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06988_ team_03_WB.instance_to_wrap.core.decoder.inst\[14\] _02827_ _02829_ vssd1
+ vssd1 vccd1 vccd1 _02930_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_126_2958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08727_ net1046 team_03_WB.instance_to_wrap.core.register_file.registers_state\[580\]
+ net998 team_03_WB.instance_to_wrap.core.register_file.registers_state\[612\] net943
+ vssd1 vssd1 vccd1 vccd1 _04669_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout835_A _06387_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09510__A1 net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1198_X net1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08658_ net1057 team_03_WB.instance_to_wrap.core.register_file.registers_state\[199\]
+ net1010 team_03_WB.instance_to_wrap.core.register_file.registers_state\[231\] net930
+ vssd1 vssd1 vccd1 vccd1 _04600_ sky130_fd_sc_hd__a221o_1
XFILLER_0_166_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_1_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07609_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[953\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[921\]
+ net789 vssd1 vssd1 vccd1 vccd1 _03551_ sky130_fd_sc_hd__mux2_1
X_08589_ net867 _04530_ _04525_ net851 vssd1 vssd1 vccd1 vccd1 _04531_ sky130_fd_sc_hd__o211a_1
XANTENNA__11423__S net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10620_ net2760 team_03_WB.instance_to_wrap.CPU_DAT_O\[9\] net840 vssd1 vssd1 vccd1
+ vccd1 _02508_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08077__A1 net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10959__A1 _06538_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_1107 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_882 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09813__A2 _05545_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10551_ net1144 _06293_ _06292_ vssd1 vssd1 vccd1 vccd1 _06294_ sky130_fd_sc_hd__a21oi_4
XANTENNA__07824__A1 net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11620__A2 net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07696__X _03638_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10482_ net119 net1029 net906 net1765 vssd1 vssd1 vccd1 vccd1 _02627_ sky130_fd_sc_hd__a22o_1
X_13270_ net1257 vssd1 vssd1 vccd1 vccd1 _01034_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout992_X net992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_727 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07037__C1 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12221_ net2310 vssd1 vssd1 vccd1 vccd1 _01436_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__11384__A1 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08785__C1 net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12152_ net1505 vssd1 vssd1 vccd1 vccd1 _02401_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__08033__A net1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11103_ _06627_ net2644 net416 vssd1 vssd1 vccd1 vccd1 _02252_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_169_wb_clk_i clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_169_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_12083_ _06787_ net459 net440 net2217 vssd1 vssd1 vccd1 vccd1 _01464_ sky130_fd_sc_hd__a22o_1
XFILLER_0_60_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08537__C1 net1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11034_ net2216 net422 _06592_ net507 vssd1 vssd1 vccd1 vccd1 _02286_ sky130_fd_sc_hd__a22o_1
XANTENNA__08001__A1 net1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11687__A2 net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input17_X net17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11439__A2 net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12985_ net1352 vssd1 vssd1 vccd1 vccd1 _00749_ sky130_fd_sc_hd__inv_2
XANTENNA__10647__A0 team_03_WB.instance_to_wrap.core.decoder.inst\[14\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14724_ clknet_leaf_50_wb_clk_i _02488_ _01089_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.decoder.inst\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09799__A _03489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_596 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11936_ net264 net2631 net370 vssd1 vssd1 vccd1 vccd1 _01606_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14655_ clknet_leaf_168_wb_clk_i _02419_ _01020_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1009\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_129_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11867_ net295 net2195 net378 vssd1 vssd1 vccd1 vccd1 _01673_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13606_ net1317 vssd1 vssd1 vccd1 vccd1 _01370_ sky130_fd_sc_hd__inv_2
XANTENNA__13114__A net1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08068__A1 net1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10818_ net691 _05541_ vssd1 vssd1 vccd1 vccd1 _06423_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_60_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14586_ clknet_leaf_148_wb_clk_i _02350_ _00951_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[940\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_39_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_144_318 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09804__A2 _05735_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11798_ net2503 _06627_ net327 vssd1 vssd1 vccd1 vccd1 _01740_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07276__C1 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13537_ net1317 vssd1 vssd1 vccd1 vccd1 _01301_ sky130_fd_sc_hd__inv_2
XFILLER_0_171_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10749_ team_03_WB.instance_to_wrap.core.pc.current_pc\[7\] net604 vssd1 vssd1 vccd1
+ vccd1 _06367_ sky130_fd_sc_hd__or2_1
XFILLER_0_153_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11611__A2 net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13468_ net1327 vssd1 vssd1 vccd1 vccd1 _01232_ sky130_fd_sc_hd__inv_2
XANTENNA__06951__A team_03_WB.instance_to_wrap.core.decoder.inst\[25\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08642__S net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09568__B2 _02945_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12419_ net1374 vssd1 vssd1 vccd1 vccd1 _00183_ sky130_fd_sc_hd__inv_2
X_13399_ net1431 vssd1 vssd1 vccd1 vccd1 _01163_ sky130_fd_sc_hd__inv_2
Xoutput205 net205 vssd1 vssd1 vccd1 vccd1 gpio_oeb[9] sky130_fd_sc_hd__buf_2
XANTENNA__07579__B1 net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput216 net216 vssd1 vssd1 vccd1 vccd1 gpio_out[19] sky130_fd_sc_hd__buf_2
XFILLER_0_2_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput227 net227 vssd1 vssd1 vccd1 vccd1 gpio_out[30] sky130_fd_sc_hd__clkbuf_4
XANTENNA__08776__C1 net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput238 net238 vssd1 vssd1 vccd1 vccd1 wbs_ack_o sky130_fd_sc_hd__buf_2
XANTENNA__08240__A1 net1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput249 net249 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[21] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_58_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15069_ net1455 vssd1 vssd1 vccd1 vccd1 la_data_out[5] sky130_fd_sc_hd__buf_2
X_07960_ net613 _03901_ vssd1 vssd1 vccd1 vccd1 _03902_ sky130_fd_sc_hd__nor2_1
XANTENNA__08528__C1 net1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11575__Y _06801_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06911_ net1154 net881 vssd1 vssd1 vccd1 vccd1 _02853_ sky130_fd_sc_hd__nand2_1
XFILLER_0_65_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11678__A2 net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07891_ net807 _03828_ _03831_ _03832_ vssd1 vssd1 vccd1 vccd1 _03833_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_147_3394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_155_Right_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11508__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09630_ net539 _05571_ vssd1 vssd1 vccd1 vccd1 _05572_ sky130_fd_sc_hd__nand2_1
XANTENNA__09740__A1 net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06842_ net1154 vssd1 vssd1 vccd1 vccd1 _02785_ sky130_fd_sc_hd__inv_2
X_09561_ _05308_ _05501_ _05182_ _05190_ vssd1 vssd1 vccd1 vccd1 _05503_ sky130_fd_sc_hd__a211oi_1
XTAP_TAPCELL_ROW_104_2508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_104_2519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10638__A0 net1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08512_ _04452_ _04453_ net859 vssd1 vssd1 vccd1 vccd1 _04454_ sky130_fd_sc_hd__o21a_1
X_09492_ _05313_ _05432_ _05320_ vssd1 vssd1 vccd1 vccd1 _05434_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_19_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07503__B1 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_2855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08443_ net541 _04384_ vssd1 vssd1 vccd1 vccd1 _04385_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_121_2866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_173_3922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_173_3933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08374_ net1207 _04312_ _04315_ net851 vssd1 vssd1 vccd1 vccd1 _04316_ sky130_fd_sc_hd__o31a_1
XFILLER_0_135_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08118__A net1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07325_ net1182 team_03_WB.instance_to_wrap.core.register_file.registers_state\[221\]
+ net768 team_03_WB.instance_to_wrap.core.register_file.registers_state\[253\] net744
+ vssd1 vssd1 vccd1 vccd1 _03267_ sky130_fd_sc_hd__o221a_1
XANTENNA__15012__Q team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[31\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12863__A net1347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10086__C net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout416_A _06610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_554 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1158_A net1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10810__B1 net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07256_ net1096 team_03_WB.instance_to_wrap.core.register_file.registers_state\[360\]
+ net896 vssd1 vssd1 vccd1 vccd1 _03198_ sky130_fd_sc_hd__or3_1
XFILLER_0_6_774 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_30_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07187_ net1115 _03123_ _03124_ _03126_ _03128_ vssd1 vssd1 vccd1 vccd1 _03129_ sky130_fd_sc_hd__o32a_1
XFILLER_0_170_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1325_A net1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11366__A1 net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07168__S net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout785_A net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1113_X net1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout410 _06684_ vssd1 vssd1 vccd1 vccd1 net410 sky130_fd_sc_hd__clkbuf_8
Xfanout1408 net1437 vssd1 vssd1 vccd1 vccd1 net1408 sky130_fd_sc_hd__clkbuf_4
Xfanout1419 net1422 vssd1 vssd1 vccd1 vccd1 net1419 sky130_fd_sc_hd__buf_4
Xfanout421 _06560_ vssd1 vssd1 vccd1 vccd1 net421 sky130_fd_sc_hd__buf_4
Xfanout432 net437 vssd1 vssd1 vccd1 vccd1 net432 sky130_fd_sc_hd__buf_2
Xfanout443 net446 vssd1 vssd1 vccd1 vccd1 net443 sky130_fd_sc_hd__buf_6
Xfanout454 net457 vssd1 vssd1 vccd1 vccd1 net454 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout952_A net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout465 net472 vssd1 vssd1 vccd1 vccd1 net465 sky130_fd_sc_hd__clkbuf_2
XANTENNA__11418__S net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout476 net481 vssd1 vssd1 vccd1 vccd1 net476 sky130_fd_sc_hd__buf_2
X_09828_ _05442_ _05669_ net574 vssd1 vssd1 vccd1 vccd1 _05770_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_122_Right_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout487 _06680_ vssd1 vssd1 vccd1 vccd1 net487 sky130_fd_sc_hd__buf_4
Xfanout498 net500 vssd1 vssd1 vccd1 vccd1 net498 sky130_fd_sc_hd__clkbuf_2
X_09759_ _03243_ net537 _04922_ _05700_ vssd1 vssd1 vccd1 vccd1 _05701_ sky130_fd_sc_hd__o31a_1
XANTENNA_fanout740_X net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10892__A3 net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout838_X net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08917__S0 net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08298__A1 net1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12770_ net1296 vssd1 vssd1 vccd1 vccd1 _00534_ sky130_fd_sc_hd__inv_2
XANTENNA__08298__B2 net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11721_ net2107 net275 net335 vssd1 vssd1 vccd1 vccd1 _01815_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_81_2040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11841__A2 net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_739 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_154_605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14440_ clknet_leaf_12_wb_clk_i _02204_ _00805_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[794\]
+ sky130_fd_sc_hd__dfrtp_1
X_11652_ net2752 _06618_ net342 vssd1 vssd1 vccd1 vccd1 _01881_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08028__A net1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10603_ net1873 net2783 net840 vssd1 vssd1 vccd1 vccd1 _02525_ sky130_fd_sc_hd__mux2_1
XANTENNA__09798__A1 net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07258__C1 net1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11054__B1 net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14371_ clknet_leaf_34_wb_clk_i _02135_ _00736_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[725\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_817 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11583_ net276 net2532 net450 vssd1 vssd1 vccd1 vccd1 _01946_ sky130_fd_sc_hd__mux2_1
XANTENNA__10801__A0 _06409_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13322_ net1308 vssd1 vssd1 vccd1 vccd1 _01086_ sky130_fd_sc_hd__inv_2
XANTENNA_input81_A wbs_adr_i[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10534_ net163 net1031 net1023 net1644 vssd1 vssd1 vccd1 vccd1 _02576_ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_150_833 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11389__A net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10465_ team_03_WB.instance_to_wrap.core.pc.current_pc\[3\] net683 _06275_ _06278_
+ vssd1 vssd1 vccd1 vccd1 _02637_ sky130_fd_sc_hd__o22a_1
XFILLER_0_122_535 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13253_ net1348 vssd1 vssd1 vccd1 vccd1 _01017_ sky130_fd_sc_hd__inv_2
XFILLER_0_122_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_161_1137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12204_ net1534 vssd1 vssd1 vccd1 vccd1 _02349_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__08222__A1 net1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10396_ net284 _06143_ _06220_ net680 vssd1 vssd1 vccd1 vccd1 _06223_ sky130_fd_sc_hd__o31a_1
X_13184_ net1403 vssd1 vssd1 vccd1 vccd1 _00948_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_36_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11676__X _06806_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07576__A3 net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08773__A2 net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12135_ net1503 vssd1 vssd1 vccd1 vccd1 _02418_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__10580__A2 net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07981__B1 _02871_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12066_ _06528_ net2754 net357 vssd1 vssd1 vccd1 vccd1 _01480_ sky130_fd_sc_hd__mux2_1
XFILLER_0_159_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_8_Left_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_53_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11328__S net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11017_ net703 net273 net827 vssd1 vssd1 vccd1 vccd1 _06582_ sky130_fd_sc_hd__and3_2
XFILLER_0_95_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07733__B1 net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08930__C1 net1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_142_3291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12968_ net1295 vssd1 vssd1 vccd1 vccd1 _00732_ sky130_fd_sc_hd__inv_2
XANTENNA__08637__S net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_66_wb_clk_i clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_66_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_clkbuf_leaf_36_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09322__A _04711_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14707_ clknet_leaf_47_wb_clk_i _02471_ _01072_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.control_logic.instruction\[4\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_169_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11919_ _06620_ net2324 net368 vssd1 vssd1 vccd1 vccd1 _01623_ sky130_fd_sc_hd__mux2_1
XANTENNA__11832__A2 net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_966 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12899_ net1356 vssd1 vssd1 vccd1 vccd1 _00663_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_44 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_238 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14638_ clknet_leaf_130_wb_clk_i _02402_ _01003_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[992\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_56_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14569_ clknet_leaf_78_wb_clk_i _02333_ _00934_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[923\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12683__A net1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07110_ _03050_ _03051_ net815 vssd1 vssd1 vccd1 vccd1 _03052_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_15_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08090_ _04031_ vssd1 vssd1 vccd1 vccd1 _04032_ sky130_fd_sc_hd__inv_2
XANTENNA__08461__A1 net1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10474__Y _06285_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10915__B _06503_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload20 clknet_leaf_8_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload20/Y sky130_fd_sc_hd__clkinv_4
X_07041_ net1100 team_03_WB.instance_to_wrap.core.register_file.registers_state\[323\]
+ net801 team_03_WB.instance_to_wrap.core.register_file.registers_state\[355\] net1155
+ vssd1 vssd1 vccd1 vccd1 _02983_ sky130_fd_sc_hd__a221o_1
XFILLER_0_71_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload31 clknet_leaf_177_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload31/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_28_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload42 clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload42/Y sky130_fd_sc_hd__bufinv_16
Xclkload53 clknet_leaf_11_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload53/Y sky130_fd_sc_hd__clkinv_2
XANTENNA__11348__A1 net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload64 clknet_leaf_46_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload64/Y sky130_fd_sc_hd__clkinv_1
XTAP_TAPCELL_ROW_77_1953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_1964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload75 clknet_leaf_55_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload75/X sky130_fd_sc_hd__clkbuf_8
XANTENNA__08213__A1 net1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload86 clknet_leaf_35_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload86/X sky130_fd_sc_hd__clkbuf_8
Xclkload97 clknet_leaf_67_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload97/Y sky130_fd_sc_hd__inv_8
XTAP_TAPCELL_ROW_149_3434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10931__A _06517_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08992_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[426\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[394\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[298\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[266\]
+ net955 net1070 vssd1 vssd1 vccd1 vccd1 _04934_ sky130_fd_sc_hd__mux4_1
XFILLER_0_76_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10571__A2 net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_166_3781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07943_ net1181 team_03_WB.instance_to_wrap.core.register_file.registers_state\[727\]
+ net766 team_03_WB.instance_to_wrap.core.register_file.registers_state\[759\] net743
+ vssd1 vssd1 vccd1 vccd1 _03885_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_166_3792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_75_wb_clk_i_A clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09713__A1 _05551_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07874_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[59\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[27\]
+ net783 vssd1 vssd1 vccd1 vccd1 _03816_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_3_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_3_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09613_ _03280_ _04532_ net665 _05554_ vssd1 vssd1 vccd1 vccd1 _05555_ sky130_fd_sc_hd__a22o_1
X_06825_ team_03_WB.instance_to_wrap.core.pc.current_pc\[27\] vssd1 vssd1 vccd1 vccd1
+ _02768_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_123_2906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11184__D net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout366_A _06815_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09544_ _05405_ _05414_ net560 vssd1 vssd1 vccd1 vccd1 _05486_ sky130_fd_sc_hd__mux2_1
XANTENNA__12076__A2 net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09232__A _04415_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11481__B net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11284__B1 net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09475_ net543 _04179_ _05083_ vssd1 vssd1 vccd1 vccd1 _05417_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12069__S net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout533_A _06298_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08426_ _04362_ _04367_ net871 vssd1 vssd1 vccd1 vccd1 _04368_ sky130_fd_sc_hd__mux2_1
XFILLER_0_164_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_164_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_163_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout321_X net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout700_A _06561_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08357_ net939 _04297_ _04298_ vssd1 vssd1 vccd1 vccd1 _04299_ sky130_fd_sc_hd__o21a_1
XANTENNA__06862__Y _02804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_783 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout419_X net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload3 clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload3/X sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout1063_X net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_468 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07308_ net1185 team_03_WB.instance_to_wrap.core.register_file.registers_state\[989\]
+ net769 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1021\] net1162
+ vssd1 vssd1 vccd1 vccd1 _03250_ sky130_fd_sc_hd__o221a_1
XFILLER_0_33_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08282__S net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10384__Y _06213_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08288_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[887\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[855\]
+ net963 vssd1 vssd1 vccd1 vccd1 _04230_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_861 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07239_ net1191 team_03_WB.instance_to_wrap.core.register_file.registers_state\[840\]
+ net774 team_03_WB.instance_to_wrap.core.register_file.registers_state\[872\] net1131
+ vssd1 vssd1 vccd1 vccd1 _03181_ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout1230_X net1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1328_X net1328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10250_ _03426_ _06090_ vssd1 vssd1 vccd1 vccd1 _06092_ sky130_fd_sc_hd__or2_1
XANTENNA__12000__A2 _06756_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout788_X net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10181_ _04646_ team_03_WB.instance_to_wrap.core.pc.current_pc\[8\] net675 vssd1
+ vssd1 vccd1 vccd1 _06023_ sky130_fd_sc_hd__mux2_1
XANTENNA__10562__A2 net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1205 net1206 vssd1 vssd1 vccd1 vccd1 net1205 sky130_fd_sc_hd__buf_2
XFILLER_0_121_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1216 team_03_WB.instance_to_wrap.core.decoder.inst\[17\] vssd1 vssd1 vccd1
+ vccd1 net1216 sky130_fd_sc_hd__clkbuf_8
Xfanout1227 net1238 vssd1 vssd1 vccd1 vccd1 net1227 sky130_fd_sc_hd__clkbuf_4
Xfanout1238 team_03_WB.instance_to_wrap.core.decoder.inst\[15\] vssd1 vssd1 vccd1
+ vccd1 net1238 sky130_fd_sc_hd__buf_4
XANTENNA_fanout955_X net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1249 net1250 vssd1 vssd1 vccd1 vccd1 net1249 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09704__A1 net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout273 _06473_ vssd1 vssd1 vccd1 vccd1 net273 sky130_fd_sc_hd__buf_2
X_13940_ clknet_leaf_134_wb_clk_i _01704_ _00305_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[294\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_31_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout284 net286 vssd1 vssd1 vccd1 vccd1 net284 sky130_fd_sc_hd__clkbuf_4
Xfanout295 _06523_ vssd1 vssd1 vccd1 vccd1 net295 sky130_fd_sc_hd__buf_2
XANTENNA__09180__A2 _04807_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13871_ clknet_leaf_135_wb_clk_i _01635_ _00236_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[225\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07810__S0 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12768__A net1402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12822_ net1280 vssd1 vssd1 vccd1 vccd1 _00586_ sky130_fd_sc_hd__inv_2
XFILLER_0_9_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11391__B net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12753_ net1267 vssd1 vssd1 vccd1 vccd1 _00517_ sky130_fd_sc_hd__inv_2
XFILLER_0_96_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11814__A2 net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11704_ _06746_ net385 net340 net2259 vssd1 vssd1 vccd1 vccd1 _01830_ sky130_fd_sc_hd__a22o_1
XFILLER_0_16_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12684_ net1332 vssd1 vssd1 vccd1 vccd1 _00448_ sky130_fd_sc_hd__inv_2
XFILLER_0_167_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13599__A net1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14423_ clknet_leaf_110_wb_clk_i _02187_ _00788_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[777\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11635_ _06709_ net386 net349 net2329 vssd1 vssd1 vccd1 vccd1 _01897_ sky130_fd_sc_hd__a22o_1
XFILLER_0_25_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_102 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07597__A net1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08192__S net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14354_ clknet_leaf_166_wb_clk_i _02118_ _00719_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[708\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input84_X net84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11566_ net505 net633 _06675_ net484 net1875 vssd1 vssd1 vccd1 vccd1 _01958_ sky130_fd_sc_hd__a32o_1
XANTENNA__08045__X _03987_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_184_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_184_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_135_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13305_ net1333 vssd1 vssd1 vccd1 vccd1 _01069_ sky130_fd_sc_hd__inv_2
X_10517_ net150 net1032 net1023 net1735 vssd1 vssd1 vccd1 vccd1 _02593_ sky130_fd_sc_hd__a22o_1
XFILLER_0_122_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07651__C1 net1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14285_ clknet_leaf_188_wb_clk_i _02049_ _00650_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[639\]
+ sky130_fd_sc_hd__dfrtp_1
X_11497_ _06618_ net2711 net389 vssd1 vssd1 vccd1 vccd1 _02009_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_113_wb_clk_i clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_113_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_13236_ net1318 vssd1 vssd1 vccd1 vccd1 _01000_ sky130_fd_sc_hd__inv_2
XFILLER_0_122_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10448_ _06264_ _06263_ net285 vssd1 vssd1 vccd1 vccd1 _06265_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_55_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_2297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_55_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07403__C1 net1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13167_ net1338 vssd1 vssd1 vccd1 vccd1 _00931_ sky130_fd_sc_hd__inv_2
X_10379_ net282 _06207_ _06208_ vssd1 vssd1 vccd1 vccd1 _06209_ sky130_fd_sc_hd__nand3_1
XFILLER_0_0_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_1850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12118_ net1143 net914 vssd1 vssd1 vccd1 vccd1 net239 sky130_fd_sc_hd__or2_1
XANTENNA__09317__A net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_1861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13098_ net1284 vssd1 vssd1 vccd1 vccd1 _00862_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_144_3331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_3342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11285__C net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12049_ _06618_ net2751 net356 vssd1 vssd1 vccd1 vccd1 _01497_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07182__A1 net1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12678__A net1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_159_wb_clk_i_A clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_07590_ net1205 team_03_WB.instance_to_wrap.core.register_file.registers_state\[185\]
+ vssd1 vssd1 vccd1 vccd1 _03532_ sky130_fd_sc_hd__and2_1
XANTENNA__08367__S net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11266__B1 net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09260_ net589 _05200_ vssd1 vssd1 vccd1 vccd1 _05202_ sky130_fd_sc_hd__nand2_1
XANTENNA__08891__A net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11018__B1 net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08211_ net1232 team_03_WB.instance_to_wrap.core.register_file.registers_state\[177\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[145\] net960 net918
+ vssd1 vssd1 vccd1 vccd1 _04153_ sky130_fd_sc_hd__a221o_1
X_09191_ _05131_ _05132_ vssd1 vssd1 vccd1 vccd1 _05133_ sky130_fd_sc_hd__nor2_1
XFILLER_0_172_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11569__A1 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08142_ net1219 _02820_ vssd1 vssd1 vccd1 vccd1 _04084_ sky130_fd_sc_hd__nand2_1
XANTENNA_wire589_X net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07300__A team_03_WB.instance_to_wrap.core.decoder.inst\[29\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_160_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload120 clknet_leaf_164_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload120/Y sky130_fd_sc_hd__inv_6
X_08073_ net1088 team_03_WB.instance_to_wrap.core.register_file.registers_state\[662\]
+ net893 net1128 vssd1 vssd1 vccd1 vccd1 _04015_ sky130_fd_sc_hd__a211o_1
XFILLER_0_125_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_2754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload131 clknet_leaf_145_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload131/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_102_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_116_2765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_1132 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload142 clknet_leaf_76_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload142/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload153 clknet_leaf_83_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload153/Y sky130_fd_sc_hd__clkinv_2
X_07024_ net748 _02964_ _02965_ net1165 vssd1 vssd1 vccd1 vccd1 _02966_ sky130_fd_sc_hd__a31o_1
XANTENNA__09926__S net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload164 clknet_leaf_108_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload164/Y sky130_fd_sc_hd__clkinv_4
Xclkload175 clknet_leaf_91_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload175/Y sky130_fd_sc_hd__inv_8
XTAP_TAPCELL_ROW_168_3821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_168_3832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10932__Y _06519_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1023_A net1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11741__A1 net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09227__A _03280_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08975_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[937\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[905\]
+ net993 vssd1 vssd1 vccd1 vccd1 _04917_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout483_A _06779_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold15 team_03_WB.instance_to_wrap.core.register_file.registers_state\[931\] vssd1
+ vssd1 vccd1 vccd1 net1508 sky130_fd_sc_hd__dlygate4sd3_1
Xhold26 team_03_WB.instance_to_wrap.core.register_file.registers_state\[932\] vssd1
+ vssd1 vccd1 vccd1 net1519 sky130_fd_sc_hd__dlygate4sd3_1
Xhold37 team_03_WB.instance_to_wrap.core.register_file.registers_state\[949\] vssd1
+ vssd1 vccd1 vccd1 net1530 sky130_fd_sc_hd__dlygate4sd3_1
X_07926_ net1181 team_03_WB.instance_to_wrap.core.register_file.registers_state\[55\]
+ net876 vssd1 vssd1 vccd1 vccd1 _03868_ sky130_fd_sc_hd__and3_1
Xhold48 team_03_WB.instance_to_wrap.core.register_file.registers_state\[958\] vssd1
+ vssd1 vccd1 vccd1 net1541 sky130_fd_sc_hd__dlygate4sd3_1
Xhold59 team_03_WB.instance_to_wrap.ADR_I\[1\] vssd1 vssd1 vccd1 vccd1 net1552 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09698__B1 _04820_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07970__A net1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07857_ net1202 team_03_WB.instance_to_wrap.core.register_file.registers_state\[859\]
+ net783 team_03_WB.instance_to_wrap.core.register_file.registers_state\[891\] net1167
+ vssd1 vssd1 vccd1 vccd1 _03799_ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout650_A net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout271_X net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout748_A net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1392_A net1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08370__B1 net1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout369_X net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10600__S net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07788_ net1086 team_03_WB.instance_to_wrap.core.register_file.registers_state\[971\]
+ net795 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1003\] net1125
+ vssd1 vssd1 vccd1 vccd1 _03730_ sky130_fd_sc_hd__a221o_1
XFILLER_0_97_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09527_ _05349_ _05360_ net553 vssd1 vssd1 vccd1 vccd1 _05469_ sky130_fd_sc_hd__mux2_1
XANTENNA__08348__S1 net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_503 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout915_A net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1180_X net1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout536_X net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08122__B1 net1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1278_X net1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09458_ _05129_ _05131_ vssd1 vssd1 vccd1 vccd1 _05400_ sky130_fd_sc_hd__nor2_1
XFILLER_0_137_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_750 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_148_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08409_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[889\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[857\]
+ net991 vssd1 vssd1 vccd1 vccd1 _04351_ sky130_fd_sc_hd__mux2_1
XFILLER_0_163_232 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09389_ _05306_ _05307_ _05311_ _05330_ vssd1 vssd1 vccd1 vccd1 _05331_ sky130_fd_sc_hd__o31a_1
XANTENNA_fanout703_X net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11431__S net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_163_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11420_ _06503_ _06751_ vssd1 vssd1 vccd1 vccd1 _06754_ sky130_fd_sc_hd__nor2_1
XANTENNA__08425__A1 net1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07633__C1 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11351_ net300 net711 net696 vssd1 vssd1 vccd1 vccd1 _06728_ sky130_fd_sc_hd__and3_1
XFILLER_0_22_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10302_ team_03_WB.instance_to_wrap.core.pc.current_pc\[17\] team_03_WB.instance_to_wrap.core.pc.current_pc\[16\]
+ _06142_ vssd1 vssd1 vccd1 vccd1 _06144_ sky130_fd_sc_hd__and3_2
XFILLER_0_85_1097 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14070_ clknet_leaf_154_wb_clk_i _01834_ _00435_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[424\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_89_Left_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11282_ net503 net632 _06708_ net410 net1911 vssd1 vssd1 vccd1 vccd1 _02154_ sky130_fd_sc_hd__a32o_1
X_13021_ net1382 vssd1 vssd1 vccd1 vccd1 _00785_ sky130_fd_sc_hd__inv_2
X_10233_ _06074_ vssd1 vssd1 vccd1 vccd1 _06075_ sky130_fd_sc_hd__inv_2
XFILLER_0_30_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10535__A2 net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11732__A1 _06509_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07936__B1 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input44_A gpio_in[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10164_ _03724_ _06005_ vssd1 vssd1 vccd1 vccd1 _06006_ sky130_fd_sc_hd__and2_1
XANTENNA__09137__A net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1002 net1003 vssd1 vssd1 vccd1 vccd1 net1002 sky130_fd_sc_hd__clkbuf_4
Xfanout1013 _04085_ vssd1 vssd1 vccd1 vccd1 net1013 sky130_fd_sc_hd__clkbuf_4
Xfanout1024 net1025 vssd1 vssd1 vccd1 vccd1 net1024 sky130_fd_sc_hd__clkbuf_4
XANTENNA__13655__Q team_03_WB.instance_to_wrap.core.register_file.registers_state\[9\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1035 _06283_ vssd1 vssd1 vccd1 vccd1 net1035 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_50_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1046 net1060 vssd1 vssd1 vccd1 vccd1 net1046 sky130_fd_sc_hd__buf_4
X_14972_ clknet_leaf_84_wb_clk_i _02724_ _01337_ vssd1 vssd1 vccd1 vccd1 net224 sky130_fd_sc_hd__dfrtp_1
X_10095_ _05435_ _05453_ _05518_ _05938_ vssd1 vssd1 vccd1 vccd1 _05939_ sky130_fd_sc_hd__or4b_1
Xfanout1057 net1058 vssd1 vssd1 vccd1 vccd1 net1057 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_22_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1068 net1069 vssd1 vssd1 vccd1 vccd1 net1068 sky130_fd_sc_hd__buf_2
Xfanout1079 net1080 vssd1 vssd1 vccd1 vccd1 net1079 sky130_fd_sc_hd__buf_4
X_13923_ clknet_leaf_31_wb_clk_i _01687_ _00288_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[277\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_156_1058 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10838__A3 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11606__S net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13854_ clknet_leaf_121_wb_clk_i _01618_ _00219_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[208\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_98_Left_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12805_ net1351 vssd1 vssd1 vccd1 vccd1 _00569_ sky130_fd_sc_hd__inv_2
XFILLER_0_97_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11248__B1 net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13785_ clknet_leaf_162_wb_clk_i _01549_ _00150_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[139\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_48_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08113__B1 net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_160 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10997_ net640 _06570_ vssd1 vssd1 vccd1 vccd1 _06571_ sky130_fd_sc_hd__nor2_1
XANTENNA__09456__A3 _04770_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11799__A1 _06628_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12736_ net1401 vssd1 vssd1 vccd1 vccd1 _00500_ sky130_fd_sc_hd__inv_2
XFILLER_0_127_402 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08915__S net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08664__A1 net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_582 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_139_295 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12667_ net1362 vssd1 vssd1 vccd1 vccd1 _00431_ sky130_fd_sc_hd__inv_2
XANTENNA__07872__C1 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14406_ clknet_leaf_27_wb_clk_i _02170_ _00771_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[760\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_170_714 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_3190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08416__A1 net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11618_ _06692_ net382 net347 net2358 vssd1 vssd1 vccd1 vccd1 _01914_ sky130_fd_sc_hd__a22o_1
XFILLER_0_155_799 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12598_ net1257 vssd1 vssd1 vccd1 vccd1 _00362_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_96_2348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_915 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14337_ clknet_leaf_183_wb_clk_i _02101_ _00702_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[691\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_13_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11549_ net504 net632 _06659_ net484 net1698 vssd1 vssd1 vccd1 vccd1 _01968_ sky130_fd_sc_hd__a32o_1
XANTENNA__06978__A1 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold507 team_03_WB.instance_to_wrap.core.register_file.registers_state\[457\] vssd1
+ vssd1 vccd1 vccd1 net2000 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_116 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold518 net200 vssd1 vssd1 vccd1 vccd1 net2011 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_133_3098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11971__A1 net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold529 team_03_WB.instance_to_wrap.core.register_file.registers_state\[681\] vssd1
+ vssd1 vccd1 vccd1 net2022 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_1901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_994 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14268_ clknet_leaf_150_wb_clk_i _02032_ _00633_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[622\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13219_ net1358 vssd1 vssd1 vccd1 vccd1 _00983_ sky130_fd_sc_hd__inv_2
XFILLER_0_111_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14199_ clknet_leaf_111_wb_clk_i _01963_ _00564_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[553\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_111_2651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_2662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11723__A1 net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10526__A2 net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08134__A_N _03459_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1013 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1207 team_03_WB.instance_to_wrap.core.register_file.registers_state\[67\] vssd1
+ vssd1 vccd1 vccd1 net2700 sky130_fd_sc_hd__dlygate4sd3_1
X_08760_ net1208 _04701_ vssd1 vssd1 vccd1 vccd1 _04702_ sky130_fd_sc_hd__or2_1
Xhold1218 team_03_WB.instance_to_wrap.core.register_file.registers_state\[599\] vssd1
+ vssd1 vccd1 vccd1 net2711 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_81_wb_clk_i clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_81_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xhold1229 team_03_WB.instance_to_wrap.core.register_file.registers_state\[338\] vssd1
+ vssd1 vccd1 vccd1 net2722 sky130_fd_sc_hd__dlygate4sd3_1
X_07711_ net1197 team_03_WB.instance_to_wrap.core.register_file.registers_state\[461\]
+ net778 team_03_WB.instance_to_wrap.core.register_file.registers_state\[493\] net1155
+ vssd1 vssd1 vccd1 vccd1 _03653_ sky130_fd_sc_hd__o221a_1
XANTENNA__10829__A3 net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08691_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[40\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[8\]
+ net975 vssd1 vssd1 vccd1 vccd1 _04633_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_10_wb_clk_i clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_10_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__07155__A1 net1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11516__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07642_ net1119 _03582_ _03583_ vssd1 vssd1 vccd1 vccd1 _03584_ sky130_fd_sc_hd__a21o_1
XFILLER_0_73_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09213__C net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07573_ net1092 team_03_WB.instance_to_wrap.core.register_file.registers_state\[888\]
+ net895 vssd1 vssd1 vccd1 vccd1 _03515_ sky130_fd_sc_hd__or3_1
X_09312_ net609 _05125_ vssd1 vssd1 vccd1 vccd1 _05254_ sky130_fd_sc_hd__nor2_1
XFILLER_0_119_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08655__A1 net1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_146_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09243_ _04119_ _05184_ vssd1 vssd1 vccd1 vccd1 _05185_ sky130_fd_sc_hd__or2_1
XFILLER_0_75_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_146_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_2805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_446 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_157_3599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout329_A _06810_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_336 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11104__X _06628_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09174_ net436 net427 net588 net550 vssd1 vssd1 vccd1 vccd1 _05116_ sky130_fd_sc_hd__o31a_1
XFILLER_0_44_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_145_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11411__A0 _06468_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08125_ net1141 _04062_ _04064_ _04066_ net722 vssd1 vssd1 vccd1 vccd1 _04067_ sky130_fd_sc_hd__o41a_1
XANTENNA__09080__A1 net1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10943__X _06528_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1140_A net1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10094__C _05841_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1238_A team_03_WB.instance_to_wrap.core.decoder.inst\[15\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11962__A1 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08056_ net807 _03996_ _03997_ vssd1 vssd1 vccd1 vccd1 _03998_ sky130_fd_sc_hd__or3_1
XANTENNA_fanout698_A net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07007_ net1020 _02943_ vssd1 vssd1 vccd1 vccd1 _02949_ sky130_fd_sc_hd__or2_1
XFILLER_0_3_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1405_A net1408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10517__A2 net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1026_X net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11714__A1 net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07918__B1 _02872_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout865_A net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout486_X net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08958_ net1244 team_03_WB.instance_to_wrap.core.register_file.registers_state\[201\]
+ net986 team_03_WB.instance_to_wrap.core.register_file.registers_state\[233\] net945
+ vssd1 vssd1 vccd1 vccd1 _04900_ sky130_fd_sc_hd__o221a_1
X_07909_ net729 _03849_ _03850_ net1117 vssd1 vssd1 vccd1 vccd1 _03851_ sky130_fd_sc_hd__o31a_1
X_08889_ net584 _04830_ vssd1 vssd1 vccd1 vccd1 _04831_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout653_X net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07146__A1 net1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08343__B1 net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09686__A3 _04820_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11426__S net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10920_ _06507_ _06508_ _06506_ vssd1 vssd1 vccd1 vccd1 _06509_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_86_609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10851_ team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[20\] net305 vssd1
+ vssd1 vccd1 vccd1 _06450_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout820_X net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout918_X net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1090 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13570_ net1432 vssd1 vssd1 vccd1 vccd1 _01334_ sky130_fd_sc_hd__inv_2
XANTENNA__08646__A1 net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10782_ _06381_ _06382_ _06388_ net1144 vssd1 vssd1 vccd1 vccd1 _06392_ sky130_fd_sc_hd__o31a_1
XFILLER_0_52_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12521_ net1260 vssd1 vssd1 vccd1 vccd1 _00285_ sky130_fd_sc_hd__inv_2
XANTENNA__07854__C1 net1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12452_ net1376 vssd1 vssd1 vccd1 vccd1 _00216_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_43_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07578__C net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11402__A0 net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11403_ net302 net2407 net397 vssd1 vssd1 vccd1 vccd1 _02077_ sky130_fd_sc_hd__mux2_1
X_12383_ net1350 vssd1 vssd1 vccd1 vccd1 _00147_ sky130_fd_sc_hd__inv_2
XANTENNA__10756__A2 net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11953__A1 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07875__A net1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14122_ clknet_leaf_0_wb_clk_i _01886_ _00487_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[476\]
+ sky130_fd_sc_hd__dfrtp_1
X_11334_ net492 net621 _06719_ net400 net1954 vssd1 vssd1 vccd1 vccd1 _02113_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_10_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_2245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11397__A net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14053_ clknet_leaf_14_wb_clk_i _01817_ _00418_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[407\]
+ sky130_fd_sc_hd__dfrtp_1
X_11265_ net714 net272 net830 vssd1 vssd1 vccd1 vccd1 _06700_ sky130_fd_sc_hd__and3_1
XANTENNA__10508__A2 net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07909__B1 net1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13004_ net1312 vssd1 vssd1 vccd1 vccd1 _00768_ sky130_fd_sc_hd__inv_2
X_10216_ _06023_ _03206_ vssd1 vssd1 vccd1 vccd1 _06058_ sky130_fd_sc_hd__and2b_1
X_11196_ net657 net707 net266 net699 vssd1 vssd1 vccd1 vccd1 _06679_ sky130_fd_sc_hd__and4_1
XFILLER_0_118_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10147_ team_03_WB.instance_to_wrap.core.pc.current_pc\[18\] net672 vssd1 vssd1 vccd1
+ vccd1 _05989_ sky130_fd_sc_hd__nand2_1
XFILLER_0_27_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14955_ clknet_leaf_103_wb_clk_i _02707_ _01320_ vssd1 vssd1 vccd1 vccd1 net207 sky130_fd_sc_hd__dfrtp_1
X_10078_ _02937_ _05342_ vssd1 vssd1 vccd1 vccd1 _05922_ sky130_fd_sc_hd__nor2_1
XANTENNA__07137__A1 net1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_2196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13906_ clknet_leaf_117_wb_clk_i _01670_ _00271_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[260\]
+ sky130_fd_sc_hd__dfrtp_1
X_14886_ clknet_leaf_65_wb_clk_i _02649_ _01251_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.pc.current_pc\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11563__C _06527_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13837_ clknet_leaf_183_wb_clk_i _01601_ _00202_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[191\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_98_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_67_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_139_3230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13768_ clknet_leaf_8_wb_clk_i _01532_ _00133_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[122\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10444__A1 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09330__A _04646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11641__B1 net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_63_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12719_ net1337 vssd1 vssd1 vccd1 vccd1 _00483_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_63_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13699_ clknet_leaf_31_wb_clk_i _01463_ _00064_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[53\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_143_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_135_3138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11071__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_46 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10907__C net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10995__A2 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_3149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07860__A2 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09062__A1 net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_152_3496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_2702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11944__A1 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09476__S net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07073__B1 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold304 team_03_WB.instance_to_wrap.core.register_file.registers_state\[438\] vssd1
+ vssd1 vccd1 vccd1 net1797 sky130_fd_sc_hd__dlygate4sd3_1
Xhold315 team_03_WB.instance_to_wrap.CPU_DAT_O\[29\] vssd1 vssd1 vccd1 vccd1 net1808
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07612__A2 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold326 _02571_ vssd1 vssd1 vccd1 vccd1 net1819 sky130_fd_sc_hd__dlygate4sd3_1
Xhold337 net176 vssd1 vssd1 vccd1 vccd1 net1830 sky130_fd_sc_hd__dlygate4sd3_1
Xhold348 team_03_WB.instance_to_wrap.core.register_file.registers_state\[570\] vssd1
+ vssd1 vccd1 vccd1 net1841 sky130_fd_sc_hd__dlygate4sd3_1
X_09930_ _05869_ net1922 net293 vssd1 vssd1 vccd1 vccd1 _02762_ sky130_fd_sc_hd__mux2_1
Xhold359 team_03_WB.instance_to_wrap.ADR_I\[13\] vssd1 vssd1 vccd1 vccd1 net1852 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_992 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_15_Right_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout806 net810 vssd1 vssd1 vccd1 vccd1 net806 sky130_fd_sc_hd__buf_6
XFILLER_0_1_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09861_ _05802_ _05686_ _05676_ _05659_ vssd1 vssd1 vccd1 vccd1 _05803_ sky130_fd_sc_hd__nand4b_1
Xfanout817 net820 vssd1 vssd1 vccd1 vccd1 net817 sky130_fd_sc_hd__buf_6
Xfanout828 _06558_ vssd1 vssd1 vccd1 vccd1 net828 sky130_fd_sc_hd__clkbuf_8
XANTENNA__07376__A1 net1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout839 _06386_ vssd1 vssd1 vccd1 vccd1 net839 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11172__A2 net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08112__C net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08812_ net873 _04753_ net852 vssd1 vssd1 vccd1 vccd1 _04754_ sky130_fd_sc_hd__a21oi_1
X_09792_ _05526_ _05600_ net568 vssd1 vssd1 vccd1 vccd1 _05734_ sky130_fd_sc_hd__mux2_1
Xhold1004 net212 vssd1 vssd1 vccd1 vccd1 net2497 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1015 team_03_WB.instance_to_wrap.core.register_file.registers_state\[611\] vssd1
+ vssd1 vccd1 vccd1 net2508 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1026 team_03_WB.instance_to_wrap.core.register_file.registers_state\[508\] vssd1
+ vssd1 vccd1 vccd1 net2519 sky130_fd_sc_hd__dlygate4sd3_1
X_08743_ net1052 team_03_WB.instance_to_wrap.core.register_file.registers_state\[67\]
+ net1004 team_03_WB.instance_to_wrap.core.register_file.registers_state\[99\] net942
+ vssd1 vssd1 vccd1 vccd1 _04685_ sky130_fd_sc_hd__a221o_1
Xhold1037 team_03_WB.instance_to_wrap.core.register_file.registers_state\[865\] vssd1
+ vssd1 vccd1 vccd1 net2530 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1048 team_03_WB.instance_to_wrap.core.register_file.registers_state\[140\] vssd1
+ vssd1 vccd1 vccd1 net2541 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1059 team_03_WB.instance_to_wrap.core.register_file.registers_state\[877\] vssd1
+ vssd1 vccd1 vccd1 net2552 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07128__A1 net1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13027__A net1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout279_A _06418_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10132__A0 _04354_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08674_ net1056 team_03_WB.instance_to_wrap.core.register_file.registers_state\[711\]
+ net1009 team_03_WB.instance_to_wrap.core.register_file.registers_state\[743\] net930
+ vssd1 vssd1 vccd1 vccd1 _04616_ sky130_fd_sc_hd__a221o_1
XFILLER_0_68_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07025__A net1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07625_ _03529_ _03566_ vssd1 vssd1 vccd1 vccd1 _03567_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_159_3639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11880__B1 net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_24_Right_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11192__D net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1090_A net1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1188_A net1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07556_ net1187 team_03_WB.instance_to_wrap.core.register_file.registers_state\[216\]
+ net771 team_03_WB.instance_to_wrap.core.register_file.registers_state\[248\] net745
+ vssd1 vssd1 vccd1 vccd1 _03498_ sky130_fd_sc_hd__o221a_1
XFILLER_0_9_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09240__A _04323_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10435__B2 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07836__C1 net1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11632__B1 net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07487_ _03391_ _03428_ vssd1 vssd1 vccd1 vccd1 _03429_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout613_A net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09226_ _03314_ _05160_ net607 vssd1 vssd1 vccd1 vccd1 _05168_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_118_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_522 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09157_ _05095_ _05098_ net554 vssd1 vssd1 vccd1 vccd1 _05099_ sky130_fd_sc_hd__mux2_1
XANTENNA__10199__A0 _04711_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout401_X net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08487__S0 net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08108_ net1173 team_03_WB.instance_to_wrap.core.register_file.registers_state\[730\]
+ net766 team_03_WB.instance_to_wrap.core.register_file.registers_state\[762\] net743
+ vssd1 vssd1 vccd1 vccd1 _04050_ sky130_fd_sc_hd__o221a_1
XFILLER_0_71_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08290__S net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08143__X _04085_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09088_ _05028_ _05029_ net1224 vssd1 vssd1 vccd1 vccd1 _05030_ sky130_fd_sc_hd__o21a_1
XPHY_EDGE_ROW_169_Right_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_33_Right_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout982_A net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09534__B1_N _05475_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08039_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[273\] net792
+ _03980_ vssd1 vssd1 vccd1 vccd1 _03981_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_82_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold860 team_03_WB.instance_to_wrap.core.register_file.registers_state\[334\] vssd1
+ vssd1 vccd1 vccd1 net2353 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1408_X net1408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold871 team_03_WB.instance_to_wrap.core.register_file.registers_state\[912\] vssd1
+ vssd1 vccd1 vccd1 net2364 sky130_fd_sc_hd__dlygate4sd3_1
Xhold882 team_03_WB.instance_to_wrap.core.register_file.registers_state\[347\] vssd1
+ vssd1 vccd1 vccd1 net2375 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11699__B1 net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11050_ net2673 net422 _06602_ net509 vssd1 vssd1 vccd1 vccd1 _02280_ sky130_fd_sc_hd__a22o_1
XANTENNA__08013__C1 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold893 team_03_WB.instance_to_wrap.core.register_file.registers_state\[580\] vssd1
+ vssd1 vccd1 vccd1 net2386 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout770_X net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07367__A1 net1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11163__A2 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout868_X net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10001_ _05886_ net1767 net288 vssd1 vssd1 vccd1 vccd1 _02713_ sky130_fd_sc_hd__mux2_1
XANTENNA__08022__C net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07462__S1 net1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10910__A2 _05676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_200 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14740_ clknet_leaf_68_wb_clk_i _02504_ _01105_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_11952_ net629 _06729_ net461 net364 net2287 vssd1 vssd1 vccd1 vccd1 _01591_ sky130_fd_sc_hd__a32o_1
XANTENNA__11383__C net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_42_Right_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10903_ net686 _06493_ _06494_ _06492_ vssd1 vssd1 vccd1 vccd1 _06495_ sky130_fd_sc_hd__o31a_4
XANTENNA__11871__A0 net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14671_ clknet_leaf_86_wb_clk_i _02435_ _01036_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.ADR_I\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_28_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11883_ net629 _06692_ net461 net372 net2098 vssd1 vssd1 vccd1 vccd1 _01658_ sky130_fd_sc_hd__a32o_1
XANTENNA__12776__A net1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13622_ net1420 vssd1 vssd1 vccd1 vccd1 _01386_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_45_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_699 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10834_ net313 net309 net316 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[23\]
+ vssd1 vssd1 vccd1 vccd1 _06436_ sky130_fd_sc_hd__o31a_1
XFILLER_0_67_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09816__B1 _02954_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13553_ net1416 vssd1 vssd1 vccd1 vccd1 _01317_ sky130_fd_sc_hd__inv_2
XANTENNA__11623__B1 net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10765_ team_03_WB.instance_to_wrap.core.pc.current_pc\[1\] _05082_ net604 vssd1
+ vssd1 vccd1 vccd1 _06377_ sky130_fd_sc_hd__mux2_1
XANTENNA__09292__A1 _04893_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_41_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12504_ net1375 vssd1 vssd1 vccd1 vccd1 _00268_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_41_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13484_ net1404 vssd1 vssd1 vccd1 vccd1 _01248_ sky130_fd_sc_hd__inv_2
X_10696_ _06312_ _06334_ vssd1 vssd1 vccd1 vccd1 _06335_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_54_369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_1113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12435_ net1260 vssd1 vssd1 vccd1 vccd1 _00199_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_51_Right_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10729__A2 net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07055__B1 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_130_3035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_130_3046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08252__C1 net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12366_ net1269 vssd1 vssd1 vccd1 vccd1 _00130_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_136_Right_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14105_ clknet_leaf_154_wb_clk_i _01869_ _00470_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[459\]
+ sky130_fd_sc_hd__dfrtp_1
X_11317_ _06624_ net2384 net406 vssd1 vssd1 vccd1 vccd1 _02128_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15085_ net1471 vssd1 vssd1 vccd1 vccd1 la_data_out[21] sky130_fd_sc_hd__buf_2
XANTENNA__09309__B _05126_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12297_ net1253 vssd1 vssd1 vccd1 vccd1 _00061_ sky130_fd_sc_hd__inv_2
X_14036_ clknet_leaf_134_wb_clk_i _01800_ _00401_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[390\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_120_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11248_ net515 net644 _06691_ net411 net2234 vssd1 vssd1 vccd1 vccd1 _02171_ sky130_fd_sc_hd__a32o_1
XANTENNA__11277__D net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07358__A1 net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07358__B2 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11179_ net632 _06669_ vssd1 vssd1 vccd1 vccd1 _06670_ sky130_fd_sc_hd__nor2_1
XFILLER_0_101_1141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10901__A2 net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12103__A1 net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_60_Right_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14938_ clknet_leaf_49_wb_clk_i _02693_ _01303_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_O\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_145_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11293__C _06545_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08858__A1 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_106_2550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11862__A0 _06499_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14869_ clknet_leaf_57_wb_clk_i net1824 _01234_ vssd1 vssd1 vccd1 vccd1 net126 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_159_154 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07410_ _02782_ _03351_ net613 vssd1 vssd1 vccd1 vccd1 _03352_ sky130_fd_sc_hd__mux2_1
XANTENNA__08375__S net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08390_ net1244 team_03_WB.instance_to_wrap.core.register_file.registers_state\[217\]
+ net990 team_03_WB.instance_to_wrap.core.register_file.registers_state\[249\] net947
+ vssd1 vssd1 vccd1 vccd1 _04332_ sky130_fd_sc_hd__o221a_1
XFILLER_0_174_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_102_2469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10417__A1 net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11614__B1 net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07341_ net1083 net888 team_03_WB.instance_to_wrap.core.register_file.registers_state\[156\]
+ vssd1 vssd1 vccd1 vccd1 _03283_ sky130_fd_sc_hd__o21a_1
XFILLER_0_161_67 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_154_3536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_703 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_154_3547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07272_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[809\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[777\]
+ net788 vssd1 vssd1 vccd1 vccd1 _03214_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_14_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09011_ net849 _04931_ _04937_ _04952_ vssd1 vssd1 vccd1 vccd1 _04953_ sky130_fd_sc_hd__a31o_4
XTAP_TAPCELL_ROW_171_3883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_171_3894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07046__B1 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold101 net132 vssd1 vssd1 vccd1 vccd1 net1594 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_599 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08243__C1 net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold112 team_03_WB.instance_to_wrap.core.register_file.registers_state\[971\] vssd1
+ vssd1 vccd1 vccd1 net1605 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07946__C net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold123 team_03_WB.instance_to_wrap.core.register_file.registers_state\[7\] vssd1
+ vssd1 vccd1 vccd1 net1616 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08794__B1 net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold134 team_03_WB.instance_to_wrap.core.register_file.registers_state\[10\] vssd1
+ vssd1 vccd1 vccd1 net1627 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_103_Right_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold145 team_03_WB.instance_to_wrap.ADR_I\[4\] vssd1 vssd1 vccd1 vccd1 net1638 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_650 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold156 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1018\] vssd1
+ vssd1 vccd1 vccd1 net1649 sky130_fd_sc_hd__dlygate4sd3_1
Xhold167 team_03_WB.instance_to_wrap.core.register_file.registers_state\[25\] vssd1
+ vssd1 vccd1 vccd1 net1660 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_940 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09934__S net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09913_ _05854_ _05718_ _05697_ _05686_ vssd1 vssd1 vccd1 vccd1 _05855_ sky130_fd_sc_hd__and4b_1
Xhold178 _02592_ vssd1 vssd1 vccd1 vccd1 net1671 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout603 _06295_ vssd1 vssd1 vccd1 vccd1 net603 sky130_fd_sc_hd__clkbuf_4
Xhold189 _02524_ vssd1 vssd1 vccd1 vccd1 net1682 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout614 net615 vssd1 vssd1 vccd1 vccd1 net614 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07349__A1 net1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout625 net631 vssd1 vssd1 vccd1 vccd1 net625 sky130_fd_sc_hd__buf_2
XANTENNA_fanout396_A _06752_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11145__A2 net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout636 net637 vssd1 vssd1 vccd1 vccd1 net636 sky130_fd_sc_hd__clkbuf_4
X_09844_ net582 _05785_ vssd1 vssd1 vccd1 vccd1 _05786_ sky130_fd_sc_hd__nand2_1
Xfanout647 net659 vssd1 vssd1 vccd1 vccd1 net647 sky130_fd_sc_hd__buf_4
XFILLER_0_42_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout658 net659 vssd1 vssd1 vccd1 vccd1 net658 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08641__S0 net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1103_A net1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout669 _06564_ vssd1 vssd1 vccd1 vccd1 net669 sky130_fd_sc_hd__buf_2
XANTENNA__09235__A _04235_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11484__B net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09775_ net351 _05485_ _05714_ _05716_ vssd1 vssd1 vccd1 vccd1 _05717_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout563_A net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06987_ _02838_ _02928_ vssd1 vssd1 vccd1 vccd1 _02929_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_126_2959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08726_ net1047 team_03_WB.instance_to_wrap.core.register_file.registers_state\[708\]
+ net999 team_03_WB.instance_to_wrap.core.register_file.registers_state\[740\] net928
+ vssd1 vssd1 vccd1 vccd1 _04668_ sky130_fd_sc_hd__a221o_1
XFILLER_0_69_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10656__A1 team_03_WB.instance_to_wrap.CPU_DAT_O\[5\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11853__A0 net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08657_ net1057 team_03_WB.instance_to_wrap.core.register_file.registers_state\[71\]
+ net1010 team_03_WB.instance_to_wrap.core.register_file.registers_state\[103\] net946
+ vssd1 vssd1 vccd1 vccd1 _04599_ sky130_fd_sc_hd__a221o_1
XFILLER_0_96_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout351_X net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout730_A net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout828_A _06558_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1093_X net1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_139_828 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout449_X net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07608_ net1203 team_03_WB.instance_to_wrap.core.register_file.registers_state\[601\]
+ net787 team_03_WB.instance_to_wrap.core.register_file.registers_state\[633\] net736
+ vssd1 vssd1 vccd1 vccd1 _03550_ sky130_fd_sc_hd__o221a_1
XANTENNA__08285__S net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08138__X _04080_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08588_ _04526_ _04527_ _04529_ _04528_ net938 net861 vssd1 vssd1 vccd1 vccd1 _04530_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_138_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11605__A0 _06545_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07539_ net1102 team_03_WB.instance_to_wrap.core.register_file.registers_state\[326\]
+ net799 team_03_WB.instance_to_wrap.core.register_file.registers_state\[358\] net1156
+ vssd1 vssd1 vccd1 vccd1 _03481_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_119_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout616_X net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_12_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1358_X net1358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11005__A net1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10550_ team_03_WB.instance_to_wrap.core.d_hit net687 vssd1 vssd1 vccd1 vccd1 _06293_
+ sky130_fd_sc_hd__nor2_4
XFILLER_0_148_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_147_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09209_ _04073_ _05147_ net608 vssd1 vssd1 vccd1 vccd1 _05151_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_107_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10481_ net1648 net1029 net906 net1617 vssd1 vssd1 vccd1 vccd1 _02628_ sky130_fd_sc_hd__a22o_1
XFILLER_0_134_566 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12220_ net1500 vssd1 vssd1 vccd1 vccd1 _01437_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__07037__B1 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13220__A net1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12030__B1 net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout985_X net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11384__A2 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12151_ net1764 vssd1 vssd1 vccd1 vccd1 _02402_ sky130_fd_sc_hd__clkbuf_1
X_11102_ net832 net270 vssd1 vssd1 vccd1 vccd1 _06627_ sky130_fd_sc_hd__and2_2
XANTENNA_clkbuf_4_5__f_wb_clk_i_A clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12082_ _06786_ net460 net440 net1936 vssd1 vssd1 vccd1 vccd1 _01465_ sky130_fd_sc_hd__a22o_1
Xhold690 team_03_WB.instance_to_wrap.core.register_file.registers_state\[787\] vssd1
+ vssd1 vccd1 vccd1 net2183 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08537__B1 net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11033_ net635 _06591_ vssd1 vssd1 vccd1 vccd1 _06592_ sky130_fd_sc_hd__nor2_1
XFILLER_0_21_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_34_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_138_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_138_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_86_2133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12097__B1 net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12984_ net1380 vssd1 vssd1 vccd1 vccd1 _00748_ sky130_fd_sc_hd__inv_2
XANTENNA__10647__A1 team_03_WB.instance_to_wrap.CPU_DAT_O\[14\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11844__A0 _06409_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_26_wb_clk_i_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_14723_ clknet_leaf_52_wb_clk_i _02487_ _01088_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.decoder.inst\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_115_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11935_ _06630_ net2723 net370 vssd1 vssd1 vccd1 vccd1 _01607_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09799__B _04591_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14654_ clknet_leaf_115_wb_clk_i _02418_ _01019_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1008\]
+ sky130_fd_sc_hd__dfstp_1
X_11866_ _06683_ net457 net375 net2257 vssd1 vssd1 vccd1 vccd1 _01674_ sky130_fd_sc_hd__a22o_1
X_13605_ net1329 vssd1 vssd1 vccd1 vccd1 _01369_ sky130_fd_sc_hd__inv_2
X_10817_ net302 net2200 net521 vssd1 vssd1 vccd1 vccd1 _02333_ sky130_fd_sc_hd__mux2_1
X_14585_ clknet_leaf_175_wb_clk_i _02349_ _00950_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[939\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_60_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11797_ net2337 _06505_ net329 vssd1 vssd1 vccd1 vccd1 _01741_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_60_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13536_ net1317 vssd1 vssd1 vccd1 vccd1 _01300_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_219 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07276__B1 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10748_ net1612 net529 net524 _06366_ vssd1 vssd1 vccd1 vccd1 _02442_ sky130_fd_sc_hd__a22o_1
XFILLER_0_125_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13467_ net1340 vssd1 vssd1 vccd1 vccd1 _01231_ sky130_fd_sc_hd__inv_2
X_10679_ net606 _06320_ vssd1 vssd1 vccd1 vccd1 _06321_ sky130_fd_sc_hd__nand2_1
XFILLER_0_152_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06951__B net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09568__A2 _04235_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_216 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12021__B1 net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12418_ net1360 vssd1 vssd1 vccd1 vccd1 _00182_ sky130_fd_sc_hd__inv_2
XFILLER_0_51_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13398_ net1423 vssd1 vssd1 vccd1 vccd1 _01162_ sky130_fd_sc_hd__inv_2
XFILLER_0_23_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07766__C net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput206 net206 vssd1 vssd1 vccd1 vccd1 gpio_out[0] sky130_fd_sc_hd__buf_2
Xoutput217 net217 vssd1 vssd1 vccd1 vccd1 gpio_out[20] sky130_fd_sc_hd__buf_2
XFILLER_0_26_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08776__B1 net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput228 net228 vssd1 vssd1 vccd1 vccd1 gpio_out[31] sky130_fd_sc_hd__clkbuf_4
X_12349_ net1388 vssd1 vssd1 vccd1 vccd1 _00113_ sky130_fd_sc_hd__inv_2
Xoutput239 net239 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[0] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_58_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10583__B1 net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_34_Left_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15068_ net1454 vssd1 vssd1 vccd1 vccd1 la_data_out[4] sky130_fd_sc_hd__buf_2
XANTENNA__08528__B1 net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06910_ net1132 net896 vssd1 vssd1 vccd1 vccd1 _02852_ sky130_fd_sc_hd__nor2_1
X_14019_ clknet_leaf_37_wb_clk_i _01783_ _00384_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[373\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_65_wb_clk_i_A clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__10335__B1 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07890_ net745 _03830_ net812 vssd1 vssd1 vccd1 vccd1 _03832_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_147_3384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_147_3395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10886__A1 team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[16\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06841_ net1148 vssd1 vssd1 vccd1 vccd1 _02784_ sky130_fd_sc_hd__inv_2
X_09560_ _05308_ _05501_ _05190_ vssd1 vssd1 vccd1 vccd1 _05502_ sky130_fd_sc_hd__a21o_1
XANTENNA__12088__B1 net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08894__A net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_2509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09205__D _05144_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08511_ net1227 team_03_WB.instance_to_wrap.core.register_file.registers_state\[735\]
+ net956 team_03_WB.instance_to_wrap.core.register_file.registers_state\[767\] net934
+ vssd1 vssd1 vccd1 vccd1 _04453_ sky130_fd_sc_hd__o221a_1
X_09491_ _05313_ _05320_ _05432_ vssd1 vssd1 vccd1 vccd1 _05433_ sky130_fd_sc_hd__or3_1
XANTENNA__11835__B1 net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10929__A net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_43_Left_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08442_ net431 net426 _04382_ vssd1 vssd1 vccd1 vccd1 _04384_ sky130_fd_sc_hd__or3_2
XTAP_TAPCELL_ROW_121_2856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_121_2867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07303__A net1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_826 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_173_3923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08373_ net937 _04313_ _04314_ net1063 vssd1 vssd1 vccd1 vccd1 _04315_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_173_3934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07324_ net1185 team_03_WB.instance_to_wrap.core.register_file.registers_state\[93\]
+ net768 team_03_WB.instance_to_wrap.core.register_file.registers_state\[125\] net728
+ vssd1 vssd1 vccd1 vccd1 _03266_ sky130_fd_sc_hd__o221a_1
XFILLER_0_34_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08464__C1 net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10810__A1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07255_ _03193_ _03196_ net824 vssd1 vssd1 vccd1 vccd1 _03197_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09008__A1 net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout311_A _05388_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1053_A net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout409_A _06684_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08216__C1 net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12012__B1 net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07186_ net741 _03127_ net1161 vssd1 vssd1 vccd1 vccd1 _03128_ sky130_fd_sc_hd__a21o_1
XANTENNA__11366__A2 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_52_Left_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1220_A net1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10574__B1 net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07973__A net1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout680_A net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout400 _06718_ vssd1 vssd1 vccd1 vccd1 net400 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_111_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1409 net1413 vssd1 vssd1 vccd1 vccd1 net1409 sky130_fd_sc_hd__buf_4
Xfanout411 _06684_ vssd1 vssd1 vccd1 vccd1 net411 sky130_fd_sc_hd__buf_4
XANTENNA_fanout778_A net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout422 _06560_ vssd1 vssd1 vccd1 vccd1 net422 sky130_fd_sc_hd__buf_6
XANTENNA_fanout399_X net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout433 net437 vssd1 vssd1 vccd1 vccd1 net433 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_100_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout444 net445 vssd1 vssd1 vccd1 vccd1 net444 sky130_fd_sc_hd__clkbuf_8
Xfanout455 net457 vssd1 vssd1 vccd1 vccd1 net455 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout1106_X net1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout466 net472 vssd1 vssd1 vccd1 vccd1 net466 sky130_fd_sc_hd__clkbuf_4
X_09827_ _05768_ vssd1 vssd1 vccd1 vccd1 _05769_ sky130_fd_sc_hd__inv_2
Xfanout477 net480 vssd1 vssd1 vccd1 vccd1 net477 sky130_fd_sc_hd__clkbuf_4
Xfanout488 _06680_ vssd1 vssd1 vccd1 vccd1 net488 sky130_fd_sc_hd__buf_8
Xfanout499 net500 vssd1 vssd1 vccd1 vccd1 net499 sky130_fd_sc_hd__buf_4
XANTENNA_fanout945_A net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09758_ _03243_ _04922_ _05699_ _04818_ vssd1 vssd1 vccd1 vccd1 _05700_ sky130_fd_sc_hd__a22o_1
XANTENNA__12079__B1 net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10629__A1 team_03_WB.instance_to_wrap.CPU_DAT_O\[0\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_61_Left_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08709_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[36\] net985
+ vssd1 vssd1 vccd1 vccd1 _04651_ sky130_fd_sc_hd__or2_1
XANTENNA__08917__S1 net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11826__B1 net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09689_ _04537_ net353 _05630_ vssd1 vssd1 vccd1 vccd1 _05631_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout733_X net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11434__S net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13215__A net1347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11720_ net1921 net300 net337 vssd1 vssd1 vccd1 vccd1 _01816_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_81_2041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_166_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07213__A net1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout900_X net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11651_ net2356 _06617_ net343 vssd1 vssd1 vccd1 vccd1 _01882_ sky130_fd_sc_hd__mux2_1
XANTENNA__09131__C net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10602_ net2087 net1650 net843 vssd1 vssd1 vccd1 vccd1 _02526_ sky130_fd_sc_hd__mux2_1
XANTENNA__07258__B1 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11054__A1 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14370_ clknet_leaf_184_wb_clk_i _02134_ _00735_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[724\]
+ sky130_fd_sc_hd__dfrtp_1
X_11582_ _06430_ net2694 net450 vssd1 vssd1 vccd1 vccd1 _01947_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_146_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13321_ net1318 vssd1 vssd1 vccd1 vccd1 _01085_ sky130_fd_sc_hd__inv_2
X_10533_ net164 net1032 net1024 net1622 vssd1 vssd1 vccd1 vccd1 _02577_ sky130_fd_sc_hd__a22o_1
XFILLER_0_135_864 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_150_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12003__A0 net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_70_Left_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13252_ net1370 vssd1 vssd1 vccd1 vccd1 _01016_ sky130_fd_sc_hd__inv_2
X_10464_ net285 _06277_ net683 vssd1 vssd1 vccd1 vccd1 _06278_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_150_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11389__B net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input74_A wbs_adr_i[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10293__B team_03_WB.instance_to_wrap.core.pc.current_pc\[4\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08044__A net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_161_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_150_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12203_ net1509 vssd1 vssd1 vccd1 vccd1 _02350_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_150_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13183_ net1347 vssd1 vssd1 vccd1 vccd1 _00947_ sky130_fd_sc_hd__inv_2
X_10395_ net304 net303 _06084_ _06221_ vssd1 vssd1 vccd1 vccd1 _06222_ sky130_fd_sc_hd__a211o_1
XANTENNA__07430__B1 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12134_ net1554 vssd1 vssd1 vccd1 vccd1 _02419_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_36_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12065_ _06629_ net2769 net358 vssd1 vssd1 vccd1 vccd1 _01481_ sky130_fd_sc_hd__mux2_1
XANTENNA__10120__A_N _03640_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_53_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11016_ net494 net647 _06581_ net420 net1801 vssd1 vssd1 vccd1 vccd1 _02293_ sky130_fd_sc_hd__a32o_1
XANTENNA__08930__B1 net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_149_wb_clk_i_A clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_142_3281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_142_3292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11817__B1 net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12967_ net1369 vssd1 vssd1 vccd1 vccd1 _00731_ sky130_fd_sc_hd__inv_2
XANTENNA__12085__A3 net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14706_ clknet_leaf_32_wb_clk_i _02470_ _01071_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.control_logic.instruction\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_16_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11918_ _06619_ net2635 net368 vssd1 vssd1 vccd1 vccd1 _01624_ sky130_fd_sc_hd__mux2_1
XANTENNA__10101__X _05945_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08694__C1 net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08219__A net1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12898_ net1296 vssd1 vssd1 vccd1 vccd1 _00662_ sky130_fd_sc_hd__inv_2
XFILLER_0_75_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_158_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11849_ net277 net2024 net378 vssd1 vssd1 vccd1 vccd1 _01691_ sky130_fd_sc_hd__mux2_1
X_14637_ clknet_leaf_189_wb_clk_i _02401_ _01002_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[991\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_145_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11045__B2 net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08446__C1 net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14568_ clknet_leaf_12_wb_clk_i _02332_ _00933_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[922\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_144_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06962__A net1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_35_wb_clk_i clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_35_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_109_Left_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06991__D_N team_03_WB.instance_to_wrap.core.decoder.inst\[30\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13519_ net1307 vssd1 vssd1 vccd1 vccd1 _01283_ sky130_fd_sc_hd__inv_2
XFILLER_0_42_114 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14499_ clknet_leaf_34_wb_clk_i _02263_ _00864_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[853\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_71_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload10 clknet_leaf_4_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload10/Y sky130_fd_sc_hd__inv_6
X_07040_ _02978_ _02981_ net818 vssd1 vssd1 vccd1 vccd1 _02982_ sky130_fd_sc_hd__o21ai_1
Xclkload21 clknet_leaf_9_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload21/Y sky130_fd_sc_hd__inv_8
XFILLER_0_152_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkload32 clknet_leaf_178_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload32/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_140_322 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09097__S0 net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload43 clknet_leaf_23_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload43/Y sky130_fd_sc_hd__inv_4
XFILLER_0_2_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload54 clknet_leaf_14_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload54/Y sky130_fd_sc_hd__clkinv_2
XANTENNA__11348__A2 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload65 clknet_leaf_44_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload65/X sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_77_1954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload76 clknet_leaf_56_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload76/Y sky130_fd_sc_hd__inv_6
XTAP_TAPCELL_ROW_77_1965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09410__A1 net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload87 clknet_leaf_69_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload87/Y sky130_fd_sc_hd__inv_6
XANTENNA__08889__A net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_149_3435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload98 clknet_leaf_68_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload98/Y sky130_fd_sc_hd__clkinv_4
XANTENNA__11899__A3 net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_219 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_188_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_08991_ net1045 team_03_WB.instance_to_wrap.core.register_file.registers_state\[458\]
+ net995 team_03_WB.instance_to_wrap.core.register_file.registers_state\[490\] net1070
+ vssd1 vssd1 vccd1 vccd1 _04933_ sky130_fd_sc_hd__a221o_1
XFILLER_0_76_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07972__A1 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11519__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07942_ net1182 team_03_WB.instance_to_wrap.core.register_file.registers_state\[599\]
+ net766 team_03_WB.instance_to_wrap.core.register_file.registers_state\[631\] net729
+ vssd1 vssd1 vccd1 vccd1 _03884_ sky130_fd_sc_hd__o221a_1
XANTENNA__10423__S net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_166_3782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_166_3793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_118_Left_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10859__A1 team_03_WB.instance_to_wrap.core.decoder.inst\[10\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07873_ _03813_ _03814_ net813 vssd1 vssd1 vccd1 vccd1 _03815_ sky130_fd_sc_hd__o21a_1
XANTENNA_clkbuf_4_4__f_wb_clk_i_X clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09612_ net538 _05553_ vssd1 vssd1 vccd1 vccd1 _05554_ sky130_fd_sc_hd__nand2_1
X_06824_ team_03_WB.instance_to_wrap.core.pc.current_pc\[28\] vssd1 vssd1 vccd1 vccd1
+ _02767_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_3_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06932__C1 net1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09543_ net576 _05484_ _05481_ vssd1 vssd1 vccd1 vccd1 _05485_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout359_A _06817_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11284__A1 net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09474_ _05085_ _05115_ vssd1 vssd1 vccd1 vccd1 _05416_ sky130_fd_sc_hd__nor2_1
XANTENNA__11481__C _06541_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11823__A3 net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08425_ net1220 _04365_ _04366_ vssd1 vssd1 vccd1 vccd1 _04367_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_93_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_149_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1170_A net1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1268_A net1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_959 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08356_ net1236 team_03_WB.instance_to_wrap.core.register_file.registers_state\[182\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[150\] net972 net922
+ vssd1 vssd1 vccd1 vccd1 _04298_ sky130_fd_sc_hd__a221o_1
XFILLER_0_19_689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload4 clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload4/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_73_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07307_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[957\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[925\]
+ net769 vssd1 vssd1 vccd1 vccd1 _03249_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08287_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[823\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[791\]
+ net965 vssd1 vssd1 vccd1 vccd1 _04229_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout314_X net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10795__B1 net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_119 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1435_A net1436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07238_ net1148 _03175_ _03177_ _03178_ _03179_ vssd1 vssd1 vccd1 vccd1 _03180_ sky130_fd_sc_hd__o32a_1
XFILLER_0_33_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout895_A net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07169_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[179\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[147\]
+ net763 vssd1 vssd1 vccd1 vccd1 _03111_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout1223_X net1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12000__A3 net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10180_ _06018_ _06019_ _03242_ vssd1 vssd1 vccd1 vccd1 _06022_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_121_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07963__A1 net1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11429__S net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1206 team_03_WB.instance_to_wrap.core.decoder.inst\[20\] vssd1 vssd1 vccd1
+ vccd1 net1206 sky130_fd_sc_hd__clkbuf_8
Xfanout1217 net1218 vssd1 vssd1 vccd1 vccd1 net1217 sky130_fd_sc_hd__clkbuf_4
Xfanout1228 net1229 vssd1 vssd1 vccd1 vccd1 net1228 sky130_fd_sc_hd__clkbuf_4
Xfanout1239 net1246 vssd1 vssd1 vccd1 vccd1 net1239 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07208__A net1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout850_X net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout263 _06546_ vssd1 vssd1 vccd1 vccd1 net263 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_31_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout285 net286 vssd1 vssd1 vccd1 vccd1 net285 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout948_X net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07176__C1 net1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11375__D net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout296 _06513_ vssd1 vssd1 vccd1 vccd1 net296 sky130_fd_sc_hd__buf_2
XANTENNA__09180__A3 net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13870_ clknet_leaf_131_wb_clk_i _01634_ _00235_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[224\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07810__S1 net1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12821_ net1273 vssd1 vssd1 vccd1 vccd1 _00585_ sky130_fd_sc_hd__inv_2
XFILLER_0_97_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12752_ net1401 vssd1 vssd1 vccd1 vccd1 _00516_ sky130_fd_sc_hd__inv_2
XFILLER_0_167_731 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11391__C _06545_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11703_ _06745_ net386 net341 net2019 vssd1 vssd1 vccd1 vccd1 _01831_ sky130_fd_sc_hd__a22o_1
XFILLER_0_167_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12683_ net1282 vssd1 vssd1 vccd1 vccd1 _00447_ sky130_fd_sc_hd__inv_2
XFILLER_0_127_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14422_ clknet_leaf_176_wb_clk_i _02186_ _00787_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[776\]
+ sky130_fd_sc_hd__dfrtp_1
X_11634_ _06708_ net380 net346 net2387 vssd1 vssd1 vccd1 vccd1 _01898_ sky130_fd_sc_hd__a22o_1
XANTENNA__08428__C1 net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14353_ clknet_leaf_139_wb_clk_i _02117_ _00718_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[707\]
+ sky130_fd_sc_hd__dfrtp_1
X_11565_ net515 net643 _06674_ net485 net1832 vssd1 vssd1 vccd1 vccd1 _01959_ sky130_fd_sc_hd__a32o_1
XFILLER_0_24_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_141_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13304_ net1333 vssd1 vssd1 vccd1 vccd1 _01068_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_147 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10516_ net151 net1030 net1025 net1595 vssd1 vssd1 vccd1 vccd1 _02594_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_98_2390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_480 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14284_ clknet_leaf_19_wb_clk_i _02048_ _00649_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[638\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_165_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11496_ _06617_ net2665 net388 vssd1 vssd1 vccd1 vccd1 _02010_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_878 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13235_ net1265 vssd1 vssd1 vccd1 vccd1 _00999_ sky130_fd_sc_hd__inv_2
X_10447_ team_03_WB.instance_to_wrap.core.pc.current_pc\[6\] _06135_ vssd1 vssd1 vccd1
+ vccd1 _06264_ sky130_fd_sc_hd__xor2_1
XANTENNA__10538__B1 net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_55_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_94_2298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07817__S net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13166_ net1305 vssd1 vssd1 vccd1 vccd1 _00930_ sky130_fd_sc_hd__inv_2
X_10378_ _05986_ _05987_ _06087_ vssd1 vssd1 vccd1 vccd1 _06208_ sky130_fd_sc_hd__o21ai_1
X_12117_ team_03_WB.instance_to_wrap.WRITE_I _02777_ team_03_WB.instance_to_wrap.wb.curr_state\[0\]
+ _02797_ net2650 vssd1 vssd1 vccd1 vccd1 _00009_ sky130_fd_sc_hd__a32o_1
XANTENNA__11750__A2 net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_153_wb_clk_i clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_153_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_20_397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_1851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13097_ net1255 vssd1 vssd1 vccd1 vccd1 _00861_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_72_1862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_144_3332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12048_ _06617_ net2488 net356 vssd1 vssd1 vccd1 vccd1 _01498_ sky130_fd_sc_hd__mux2_1
XANTENNA__12959__A net1347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10710__B1 net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06957__A net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_161_3690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13999_ clknet_leaf_138_wb_clk_i _01763_ _00364_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[353\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_149_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11266__A1 net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08667__C1 net1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09620__X _05562_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_904 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_303 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11802__S net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08210_ net935 _04151_ vssd1 vssd1 vccd1 vccd1 _04152_ sky130_fd_sc_hd__or2_1
XANTENNA__11018__A1 net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09190_ net434 net429 _04679_ net552 vssd1 vssd1 vccd1 vccd1 _05132_ sky130_fd_sc_hd__o31a_1
XFILLER_0_90_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07890__B1 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_604 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08236__X _04178_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11569__A2 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08141_ net1064 net1015 vssd1 vssd1 vccd1 vccd1 _04083_ sky130_fd_sc_hd__nor2_1
XFILLER_0_56_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09631__A1 _03314_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07300__B net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload110 clknet_leaf_158_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload110/Y sky130_fd_sc_hd__bufinv_16
X_08072_ net1183 team_03_WB.instance_to_wrap.core.register_file.registers_state\[694\]
+ net876 vssd1 vssd1 vccd1 vccd1 _04014_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_116_2755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload121 clknet_leaf_165_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload121/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_125_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_116_2766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload132 clknet_leaf_120_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload132/Y sky130_fd_sc_hd__inv_8
Xclkload143 clknet_leaf_77_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload143/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_114_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload154 clknet_leaf_84_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload154/Y sky130_fd_sc_hd__bufinv_16
X_07023_ net1099 team_03_WB.instance_to_wrap.core.register_file.registers_state\[675\]
+ net897 vssd1 vssd1 vccd1 vccd1 _02965_ sky130_fd_sc_hd__or3_1
XFILLER_0_11_92 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_140_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_168_3822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload165 clknet_leaf_109_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload165/Y sky130_fd_sc_hd__bufinv_16
XANTENNA__10529__B1 net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload176 clknet_leaf_92_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload176/X sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_168_3833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08198__A1 net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_1008 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_126_Left_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07945__A1 net1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07945__B2 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08974_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[809\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[777\]
+ net991 vssd1 vssd1 vccd1 vccd1 _04916_ sky130_fd_sc_hd__mux2_1
XANTENNA__09942__S net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold16 team_03_WB.instance_to_wrap.core.register_file.registers_state\[940\] vssd1
+ vssd1 vccd1 vccd1 net1509 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_89_Right_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold27 team_03_WB.instance_to_wrap.core.register_file.registers_state\[938\] vssd1
+ vssd1 vccd1 vccd1 net1520 sky130_fd_sc_hd__dlygate4sd3_1
X_07925_ net1087 net892 team_03_WB.instance_to_wrap.core.register_file.registers_state\[23\]
+ vssd1 vssd1 vccd1 vccd1 _03867_ sky130_fd_sc_hd__o21a_1
Xhold38 team_03_WB.instance_to_wrap.core.register_file.registers_state\[986\] vssd1
+ vssd1 vccd1 vccd1 net1531 sky130_fd_sc_hd__dlygate4sd3_1
Xhold49 team_03_WB.instance_to_wrap.core.register_file.registers_state\[984\] vssd1
+ vssd1 vccd1 vccd1 net1542 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout476_A net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07856_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[795\] net804
+ _03792_ net1120 vssd1 vssd1 vccd1 vccd1 _03798_ sky130_fd_sc_hd__o211a_1
XANTENNA__10701__B1 net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14857__Q net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09243__A _04119_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07787_ net1086 team_03_WB.instance_to_wrap.core.register_file.registers_state\[843\]
+ net795 team_03_WB.instance_to_wrap.core.register_file.registers_state\[875\] net1150
+ vssd1 vssd1 vccd1 vccd1 _03729_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout643_A net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout264_X net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1385_A net1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09526_ net577 _05467_ vssd1 vssd1 vccd1 vccd1 _05468_ sky130_fd_sc_hd__or2_1
XFILLER_0_79_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08658__C1 net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_515 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_135_Left_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09457_ _05137_ _05398_ net556 vssd1 vssd1 vccd1 vccd1 _05399_ sky130_fd_sc_hd__mux2_1
XFILLER_0_164_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout431_X net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1173_X net1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout908_A _06285_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout529_X net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11712__S net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08408_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[1017\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[985\]
+ net992 vssd1 vssd1 vccd1 vccd1 _04350_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_98_Right_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07881__A0 _03821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_762 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10480__A2 net1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09388_ _05321_ _05325_ _05329_ vssd1 vssd1 vccd1 vccd1 _05330_ sky130_fd_sc_hd__and3_1
XANTENNA__08146__X _04088_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08293__S net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07050__X _02992_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_244 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_795 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08339_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[53\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[21\]
+ net968 vssd1 vssd1 vccd1 vccd1 _04281_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_163_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1438_X net1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11013__A net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07633__B1 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11350_ net497 net626 _06727_ net401 net1886 vssd1 vssd1 vccd1 vccd1 _02105_ sky130_fd_sc_hd__a32o_1
XFILLER_0_160_940 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10301_ team_03_WB.instance_to_wrap.core.pc.current_pc\[16\] _06142_ vssd1 vssd1
+ vccd1 vccd1 _06143_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout898_X net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11281_ net710 _06518_ net828 vssd1 vssd1 vccd1 vccd1 _06708_ sky130_fd_sc_hd__and3_1
X_13020_ net1413 vssd1 vssd1 vccd1 vccd1 _00784_ sky130_fd_sc_hd__inv_2
X_10232_ _06071_ _06072_ _03864_ vssd1 vssd1 vccd1 vccd1 _06074_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_120_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07397__C1 net1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_1_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11193__B1 net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07936__A1 net1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10163_ _04862_ team_03_WB.instance_to_wrap.core.pc.current_pc\[12\] net674 vssd1
+ vssd1 vccd1 vccd1 _06005_ sky130_fd_sc_hd__mux2_1
Xfanout1003 net1008 vssd1 vssd1 vccd1 vccd1 net1003 sky130_fd_sc_hd__clkbuf_4
Xfanout1014 _02869_ vssd1 vssd1 vccd1 vccd1 net1014 sky130_fd_sc_hd__buf_8
Xfanout1025 _06286_ vssd1 vssd1 vccd1 vccd1 net1025 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_50_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1036 net1038 vssd1 vssd1 vccd1 vccd1 net1036 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_50_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input37_A gpio_in[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1047 net1048 vssd1 vssd1 vccd1 vccd1 net1047 sky130_fd_sc_hd__clkbuf_4
X_14971_ clknet_leaf_81_wb_clk_i _02723_ _01336_ vssd1 vssd1 vccd1 vccd1 net223 sky130_fd_sc_hd__dfrtp_1
X_10094_ _05833_ _05834_ _05841_ _05937_ vssd1 vssd1 vccd1 vccd1 _05938_ sky130_fd_sc_hd__and4_1
Xfanout1058 net1059 vssd1 vssd1 vccd1 vccd1 net1058 sky130_fd_sc_hd__clkbuf_4
Xfanout1069 _02790_ vssd1 vssd1 vccd1 vccd1 net1069 sky130_fd_sc_hd__buf_4
XFILLER_0_22_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13922_ clknet_leaf_170_wb_clk_i _01686_ _00287_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[276\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08897__C1 net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08361__A1 net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13853_ clknet_leaf_24_wb_clk_i _01617_ _00218_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[207\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_159_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12804_ net1366 vssd1 vssd1 vccd1 vccd1 _00568_ sky130_fd_sc_hd__inv_2
XANTENNA__11248__A1 net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13784_ clknet_leaf_19_wb_clk_i _01548_ _00149_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[138\]
+ sky130_fd_sc_hd__dfrtp_1
X_10996_ net714 net702 _06422_ vssd1 vssd1 vccd1 vccd1 _06570_ sky130_fd_sc_hd__or3b_1
XANTENNA__08113__A1 net1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_172 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07879__Y _03821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12735_ net1286 vssd1 vssd1 vccd1 vccd1 _00499_ sky130_fd_sc_hd__inv_2
XFILLER_0_38_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_167_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12666_ net1375 vssd1 vssd1 vccd1 vccd1 _00430_ sky130_fd_sc_hd__inv_2
XANTENNA__07872__B1 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07401__A net1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_154_255 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14405_ clknet_leaf_11_wb_clk_i _02169_ _00770_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[759\]
+ sky130_fd_sc_hd__dfrtp_1
X_11617_ _06691_ net385 net349 net2182 vssd1 vssd1 vccd1 vccd1 _01915_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_137_3180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_423 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09074__C1 net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09613__A1 _03280_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_3191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12597_ net1292 vssd1 vssd1 vccd1 vccd1 _00361_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_96_2338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07624__A0 _03563_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_96_2349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14336_ clknet_leaf_190_wb_clk_i _02100_ _00701_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[690\]
+ sky130_fd_sc_hd__dfrtp_1
X_11548_ net1948 net483 _06789_ net502 vssd1 vssd1 vccd1 vccd1 _01969_ sky130_fd_sc_hd__a22o_1
XFILLER_0_41_927 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08821__C1 net1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_133_3099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold508 team_03_WB.instance_to_wrap.core.register_file.registers_state\[869\] vssd1
+ vssd1 vccd1 vccd1 net2001 sky130_fd_sc_hd__dlygate4sd3_1
Xhold519 team_03_WB.instance_to_wrap.core.register_file.registers_state\[613\] vssd1
+ vssd1 vccd1 vccd1 net2012 sky130_fd_sc_hd__dlygate4sd3_1
X_14267_ clknet_leaf_123_wb_clk_i _02031_ _00632_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[621\]
+ sky130_fd_sc_hd__dfrtp_1
X_11479_ net515 net643 _06603_ net394 net2012 vssd1 vssd1 vccd1 vccd1 _02023_ sky130_fd_sc_hd__a32o_1
XFILLER_0_0_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_1902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_686 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07547__S net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13218_ net1287 vssd1 vssd1 vccd1 vccd1 _00982_ sky130_fd_sc_hd__inv_2
X_14198_ clknet_leaf_150_wb_clk_i _01962_ _00563_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[552\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11069__S net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_2652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07927__A1 net1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_2663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13149_ net1382 vssd1 vssd1 vccd1 vccd1 _00913_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_163_3730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1208 team_03_WB.instance_to_wrap.core.register_file.registers_state\[220\] vssd1
+ vssd1 vccd1 vccd1 net2701 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12689__A net1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1219 team_03_WB.instance_to_wrap.core.register_file.registers_state\[765\] vssd1
+ vssd1 vccd1 vccd1 net2712 sky130_fd_sc_hd__dlygate4sd3_1
X_07710_ net1197 team_03_WB.instance_to_wrap.core.register_file.registers_state\[333\]
+ net778 team_03_WB.instance_to_wrap.core.register_file.registers_state\[365\] net1134
+ vssd1 vssd1 vccd1 vccd1 _03652_ sky130_fd_sc_hd__o221a_1
X_08690_ _04626_ _04631_ net873 vssd1 vssd1 vccd1 vccd1 _04632_ sky130_fd_sc_hd__mux2_1
XANTENNA__11487__B2 net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08378__S net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07641_ _03578_ _03579_ _03581_ net1132 net1164 vssd1 vssd1 vccd1 vccd1 _03583_ sky130_fd_sc_hd__o221a_1
XFILLER_0_73_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07560__C1 net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07572_ net1120 _03507_ _03508_ _03510_ _03513_ vssd1 vssd1 vccd1 vccd1 _03514_ sky130_fd_sc_hd__o32a_1
XFILLER_0_76_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09213__D _05146_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_50_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_50_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_09311_ _04679_ _05252_ vssd1 vssd1 vccd1 vccd1 _05253_ sky130_fd_sc_hd__nor2_1
XFILLER_0_146_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09242_ _03391_ _05153_ vssd1 vssd1 vccd1 vccd1 _05184_ sky130_fd_sc_hd__xor2_1
XFILLER_0_111_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_157_3589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_118_2806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09173_ net433 net427 net589 net546 vssd1 vssd1 vccd1 vccd1 _05115_ sky130_fd_sc_hd__o31a_1
XFILLER_0_146_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09065__C1 net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08124_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[922\] net793
+ net1014 _04065_ vssd1 vssd1 vccd1 vccd1 _04066_ sky130_fd_sc_hd__o211a_1
XFILLER_0_142_962 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08055_ net1186 team_03_WB.instance_to_wrap.core.register_file.registers_state\[214\]
+ net771 team_03_WB.instance_to_wrap.core.register_file.registers_state\[246\] net745
+ vssd1 vssd1 vccd1 vccd1 _03997_ sky130_fd_sc_hd__o221a_1
XANTENNA__10672__A _05429_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1133_A net1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07006_ net608 _02940_ _02947_ vssd1 vssd1 vccd1 vccd1 _02948_ sky130_fd_sc_hd__or3_1
XANTENNA__09238__A _04323_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08142__A net1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07918__A1 net1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08040__B1 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1300_A net1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10922__B1 _06401_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1019_X net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout760_A net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout381_X net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08957_ net1244 team_03_WB.instance_to_wrap.core.register_file.registers_state\[73\]
+ net986 team_03_WB.instance_to_wrap.core.register_file.registers_state\[105\] net929
+ vssd1 vssd1 vccd1 vccd1 _04899_ sky130_fd_sc_hd__o221a_1
XANTENNA__10611__S net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07908_ net1091 team_03_WB.instance_to_wrap.core.register_file.registers_state\[655\]
+ vssd1 vssd1 vccd1 vccd1 _03850_ sky130_fd_sc_hd__and2_1
X_08888_ _02948_ _02949_ net526 vssd1 vssd1 vccd1 vccd1 _04830_ sky130_fd_sc_hd__or3b_2
XANTENNA__11478__B2 net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08288__S net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08343__A1 net1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07839_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[554\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[522\]
+ net760 vssd1 vssd1 vccd1 vccd1 _03781_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout646_X net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11008__A net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10850_ _06394_ _06447_ vssd1 vssd1 vccd1 vccd1 _06449_ sky130_fd_sc_hd__nand2_2
XFILLER_0_6_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07529__S0 net1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09509_ _05350_ _05366_ net568 vssd1 vssd1 vccd1 vccd1 _05451_ sky130_fd_sc_hd__mux2_1
XFILLER_0_149_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10781_ _06381_ _06390_ vssd1 vssd1 vccd1 vccd1 _06391_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout813_X net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_734 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12520_ net1297 vssd1 vssd1 vccd1 vccd1 _00284_ sky130_fd_sc_hd__inv_2
XFILLER_0_82_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11650__A1 _06616_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07854__B1 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07859__C net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_117_Right_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_23_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12451_ net1371 vssd1 vssd1 vccd1 vccd1 _00215_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_43_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_43_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_726 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11402_ net279 net2492 net396 vssd1 vssd1 vccd1 vccd1 _02078_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08751__S net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08803__C1 net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12382_ net1386 vssd1 vssd1 vccd1 vccd1 _00146_ sky130_fd_sc_hd__inv_2
XFILLER_0_34_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14121_ clknet_leaf_75_wb_clk_i _01885_ _00486_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[475\]
+ sky130_fd_sc_hd__dfrtp_1
X_11333_ net281 net709 net695 vssd1 vssd1 vccd1 vccd1 _06719_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_10_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_160_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_91_2246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14052_ clknet_leaf_35_wb_clk_i _01816_ _00417_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[406\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_120_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11264_ net495 net624 _06699_ net408 net2131 vssd1 vssd1 vccd1 vccd1 _02163_ sky130_fd_sc_hd__a32o_1
XANTENNA__07909__A1 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13003_ net1281 vssd1 vssd1 vccd1 vccd1 _00767_ sky130_fd_sc_hd__inv_2
XANTENNA__11705__A2 net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10215_ _06028_ _06056_ _06026_ vssd1 vssd1 vccd1 vccd1 _06057_ sky130_fd_sc_hd__a21o_1
X_11195_ net2264 net414 _06678_ net510 vssd1 vssd1 vccd1 vccd1 _02211_ sky130_fd_sc_hd__a22o_1
XANTENNA__08582__A1 net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10146_ _03109_ _05985_ vssd1 vssd1 vccd1 vccd1 _05988_ sky130_fd_sc_hd__or2_1
XFILLER_0_118_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_49 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14954_ clknet_leaf_88_wb_clk_i _02706_ _01319_ vssd1 vssd1 vccd1 vccd1 net237 sky130_fd_sc_hd__dfrtp_1
X_10077_ _03352_ _04475_ net312 vssd1 vssd1 vccd1 vccd1 _05921_ sky130_fd_sc_hd__mux2_1
XANTENNA__11469__B2 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09531__B1 net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_2197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13905_ clknet_leaf_144_wb_clk_i _01669_ _00270_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[259\]
+ sky130_fd_sc_hd__dfrtp_1
X_14885_ clknet_leaf_67_wb_clk_i _02648_ _01250_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.pc.current_pc\[14\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__11563__D net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload2_A clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13836_ clknet_leaf_18_wb_clk_i _01600_ _00201_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[190\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_67_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09611__A _03280_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_139_3220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1131 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_139_3231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10979_ net266 net2053 net520 vssd1 vssd1 vccd1 vccd1 _02306_ sky130_fd_sc_hd__mux2_1
X_13767_ clknet_leaf_106_wb_clk_i _01531_ _00132_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[121\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_167_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09860__C_N _05718_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10444__A2 _06136_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_63_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12718_ net1269 vssd1 vssd1 vccd1 vccd1 _00482_ sky130_fd_sc_hd__inv_2
X_13698_ clknet_leaf_173_wb_clk_i _01462_ _00063_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[52\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_135_3139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10907__D net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_789 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12649_ net1260 vssd1 vssd1 vccd1 vccd1 _00413_ sky130_fd_sc_hd__inv_2
XFILLER_0_143_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_288 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_152_3486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_113_2703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_152_3497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07785__B _03726_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold305 team_03_WB.instance_to_wrap.core.register_file.registers_state\[403\] vssd1
+ vssd1 vccd1 vccd1 net1798 sky130_fd_sc_hd__dlygate4sd3_1
X_14319_ clknet_leaf_134_wb_clk_i _02083_ _00684_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[673\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold316 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[18\] vssd1 vssd1 vccd1
+ vccd1 net1809 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold327 team_03_WB.instance_to_wrap.core.register_file.registers_state\[902\] vssd1
+ vssd1 vccd1 vccd1 net1820 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold338 team_03_WB.instance_to_wrap.core.register_file.registers_state\[407\] vssd1
+ vssd1 vccd1 vccd1 net1831 sky130_fd_sc_hd__dlygate4sd3_1
Xhold349 team_03_WB.instance_to_wrap.core.register_file.registers_state\[168\] vssd1
+ vssd1 vccd1 vccd1 net1842 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08248__S1 net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11875__X _06813_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09860_ _05706_ _05801_ _05718_ _05697_ vssd1 vssd1 vccd1 vccd1 _05802_ sky130_fd_sc_hd__or4bb_1
Xfanout807 net810 vssd1 vssd1 vccd1 vccd1 net807 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10904__A0 net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout818 net819 vssd1 vssd1 vccd1 vccd1 net818 sky130_fd_sc_hd__clkbuf_8
Xfanout829 net831 vssd1 vssd1 vccd1 vccd1 net829 sky130_fd_sc_hd__clkbuf_4
X_08811_ net1065 _04751_ _04752_ vssd1 vssd1 vccd1 vccd1 _04753_ sky130_fd_sc_hd__a21o_1
X_09791_ _05731_ _05732_ vssd1 vssd1 vccd1 vccd1 _05733_ sky130_fd_sc_hd__nor2_1
Xhold1005 team_03_WB.instance_to_wrap.core.register_file.registers_state\[205\] vssd1
+ vssd1 vccd1 vccd1 net2498 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1016 team_03_WB.instance_to_wrap.core.register_file.registers_state\[325\] vssd1
+ vssd1 vccd1 vccd1 net2509 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13308__A net1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08742_ _04682_ _04683_ net857 vssd1 vssd1 vccd1 vccd1 _04684_ sky130_fd_sc_hd__o21a_1
Xhold1027 team_03_WB.instance_to_wrap.core.register_file.registers_state\[646\] vssd1
+ vssd1 vccd1 vccd1 net2520 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1038 team_03_WB.instance_to_wrap.core.register_file.registers_state\[724\] vssd1
+ vssd1 vccd1 vccd1 net2531 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1049 team_03_WB.instance_to_wrap.core.register_file.registers_state\[359\] vssd1
+ vssd1 vccd1 vccd1 net2542 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08325__A1 net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08673_ net1057 team_03_WB.instance_to_wrap.core.register_file.registers_state\[583\]
+ net1011 team_03_WB.instance_to_wrap.core.register_file.registers_state\[615\] net946
+ vssd1 vssd1 vccd1 vccd1 _04615_ sky130_fd_sc_hd__a221o_1
XFILLER_0_17_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07624_ _03563_ _03565_ net610 vssd1 vssd1 vccd1 vccd1 _03566_ sky130_fd_sc_hd__mux2_2
XFILLER_0_16_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1075 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10683__A2 net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11880__A1 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08089__A0 _04029_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07555_ net1187 team_03_WB.instance_to_wrap.core.register_file.registers_state\[88\]
+ net771 team_03_WB.instance_to_wrap.core.register_file.registers_state\[120\] net729
+ vssd1 vssd1 vccd1 vccd1 _03497_ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout341_A _06806_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09825__B2 net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout439_A _06819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1083_A net1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13043__A net1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07836__B1 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07486_ _03425_ _03427_ net610 vssd1 vssd1 vccd1 vccd1 _03428_ sky130_fd_sc_hd__mux2_2
XFILLER_0_76_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09225_ _05166_ vssd1 vssd1 vccd1 vccd1 _05167_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_hold1289_A team_03_WB.instance_to_wrap.CPU_DAT_O\[3\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_17_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_372 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout606_A _06294_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_161_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_146_1003 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09156_ _05096_ _05097_ vssd1 vssd1 vccd1 vccd1 _05098_ sky130_fd_sc_hd__nor2_1
XFILLER_0_161_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10199__A1 _02774_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08487__S1 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11396__B1 net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08107_ net1172 team_03_WB.instance_to_wrap.core.register_file.registers_state\[602\]
+ vssd1 vssd1 vccd1 vccd1 _04049_ sky130_fd_sc_hd__or2_1
XFILLER_0_161_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09087_ net1240 team_03_WB.instance_to_wrap.core.register_file.registers_state\[717\]
+ net982 team_03_WB.instance_to_wrap.core.register_file.registers_state\[749\] net941
+ vssd1 vssd1 vccd1 vccd1 _05029_ sky130_fd_sc_hd__o221a_1
XFILLER_0_142_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08800__A2 net1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1136_X net1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1057 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08038_ net1086 team_03_WB.instance_to_wrap.core.register_file.registers_state\[305\]
+ net890 net1041 vssd1 vssd1 vccd1 vccd1 _03980_ sky130_fd_sc_hd__o31a_1
Xhold850 team_03_WB.instance_to_wrap.core.register_file.registers_state\[767\] vssd1
+ vssd1 vccd1 vccd1 net2343 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout975_A net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout596_X net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold861 team_03_WB.instance_to_wrap.core.register_file.registers_state\[256\] vssd1
+ vssd1 vccd1 vccd1 net2354 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08013__B1 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold872 team_03_WB.instance_to_wrap.core.register_file.registers_state\[145\] vssd1
+ vssd1 vccd1 vccd1 net2365 sky130_fd_sc_hd__dlygate4sd3_1
Xhold883 team_03_WB.instance_to_wrap.core.register_file.registers_state\[272\] vssd1
+ vssd1 vccd1 vccd1 net2376 sky130_fd_sc_hd__dlygate4sd3_1
Xhold894 team_03_WB.instance_to_wrap.core.register_file.registers_state\[488\] vssd1
+ vssd1 vccd1 vccd1 net2387 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10000_ _05885_ net1854 net290 vssd1 vssd1 vccd1 vccd1 _02714_ sky130_fd_sc_hd__mux2_1
X_09989_ _05874_ net2734 net288 vssd1 vssd1 vccd1 vccd1 _02725_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout763_X net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07772__C1 net1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10341__S net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_212 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10929__D_N team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[8\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_16_wb_clk_i_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout930_X net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11320__A0 _06505_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11951_ net628 _06728_ net459 net364 net2113 vssd1 vssd1 vccd1 vccd1 _01592_ sky130_fd_sc_hd__a32o_1
XFILLER_0_118_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_168_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10902_ team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[13\] net311 net310 net317
+ vssd1 vssd1 vccd1 vccd1 _06494_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_28_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14670_ clknet_leaf_82_wb_clk_i _02434_ _01035_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.ADR_I\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_28_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11882_ net644 _06691_ net478 net374 net2140 vssd1 vssd1 vccd1 vccd1 _01659_ sky130_fd_sc_hd__a32o_1
XFILLER_0_98_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13621_ net1428 vssd1 vssd1 vccd1 vccd1 _01385_ sky130_fd_sc_hd__inv_2
X_10833_ net686 _05517_ _06401_ vssd1 vssd1 vccd1 vccd1 _06435_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_45_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_45_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10764_ net525 _06375_ _06376_ net530 net1761 vssd1 vssd1 vccd1 vccd1 _02436_ sky130_fd_sc_hd__a32o_1
XFILLER_0_149_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13552_ net1416 vssd1 vssd1 vccd1 vccd1 _01316_ sky130_fd_sc_hd__inv_2
XFILLER_0_82_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12503_ net1386 vssd1 vssd1 vccd1 vccd1 _00267_ sky130_fd_sc_hd__inv_2
X_13483_ net1404 vssd1 vssd1 vccd1 vccd1 _01247_ sky130_fd_sc_hd__inv_2
XFILLER_0_82_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09029__C1 net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10695_ _05583_ _06311_ vssd1 vssd1 vccd1 vccd1 _06334_ sky130_fd_sc_hd__nand2_1
XFILLER_0_125_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10864__X _06463_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12792__A net1376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12434_ net1338 vssd1 vssd1 vccd1 vccd1 _00198_ sky130_fd_sc_hd__inv_2
XFILLER_0_164_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_164_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_770 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_3036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12365_ net1332 vssd1 vssd1 vccd1 vccd1 _00129_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_130_3047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14104_ clknet_leaf_185_wb_clk_i _01868_ _00469_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[458\]
+ sky130_fd_sc_hd__dfrtp_1
X_11316_ _06623_ net2619 net405 vssd1 vssd1 vccd1 vccd1 _02129_ sky130_fd_sc_hd__mux2_1
X_15084_ net1470 vssd1 vssd1 vccd1 vccd1 la_data_out[20] sky130_fd_sc_hd__buf_2
XFILLER_0_121_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12296_ net1293 vssd1 vssd1 vccd1 vccd1 _00060_ sky130_fd_sc_hd__inv_2
XFILLER_0_120_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14035_ clknet_leaf_108_wb_clk_i _01799_ _00400_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[389\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08004__B1 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11247_ net277 net715 net830 vssd1 vssd1 vccd1 vccd1 _06691_ sky130_fd_sc_hd__and3_1
XANTENNA_clkbuf_leaf_55_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_120_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10898__C1 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11178_ net710 _06517_ net694 vssd1 vssd1 vccd1 vccd1 _06669_ sky130_fd_sc_hd__or3_1
XFILLER_0_38_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10129_ _05970_ vssd1 vssd1 vccd1 vccd1 _05971_ sky130_fd_sc_hd__inv_2
XANTENNA__10901__A3 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13128__A net1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10104__X _05948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14937_ clknet_leaf_52_wb_clk_i _02692_ _01302_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_O\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11311__A0 _06454_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11293__D net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12967__A net1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_2551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_106_2562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14868_ clknet_leaf_59_wb_clk_i net1700 _01233_ vssd1 vssd1 vccd1 vccd1 net124 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_77_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08883__C _04807_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09341__A _04207_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13819_ clknet_leaf_158_wb_clk_i _01583_ _00184_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[173\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_206 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14799_ clknet_leaf_88_wb_clk_i _02563_ _01164_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_I\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_07340_ net1172 team_03_WB.instance_to_wrap.core.register_file.registers_state\[60\]
+ net880 vssd1 vssd1 vccd1 vccd1 _03282_ sky130_fd_sc_hd__and3_1
XANTENNA__10417__A2 net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_462 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_161_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_156_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_154_3537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_169_1047 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07271_ net1136 _03209_ _03210_ _03212_ net1121 vssd1 vssd1 vccd1 vccd1 _03213_ sky130_fd_sc_hd__a311o_1
XFILLER_0_116_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_14_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_14_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09010_ net850 _04944_ _04951_ vssd1 vssd1 vccd1 vccd1 _04952_ sky130_fd_sc_hd__and3_1
XFILLER_0_170_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_171_854 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_171_3884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_94_wb_clk_i_A clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_131_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11378__B1 net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_171_3895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08469__S1 net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold102 team_03_WB.instance_to_wrap.CPU_DAT_I\[23\] vssd1 vssd1 vccd1 vccd1 net1595
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold113 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[16\] vssd1 vssd1 vccd1
+ vccd1 net1606 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09991__A0 _05876_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold124 team_03_WB.instance_to_wrap.ADR_I\[25\] vssd1 vssd1 vccd1 vccd1 net1617 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10050__B1 net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08794__A1 net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold135 team_03_WB.instance_to_wrap.ADR_I\[23\] vssd1 vssd1 vccd1 vccd1 net1628 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold146 _02607_ vssd1 vssd1 vccd1 vccd1 net1639 sky130_fd_sc_hd__dlygate4sd3_1
Xhold157 team_03_WB.instance_to_wrap.CPU_DAT_O\[27\] vssd1 vssd1 vccd1 vccd1 net1650
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold168 team_03_WB.instance_to_wrap.CPU_DAT_I\[7\] vssd1 vssd1 vccd1 vccd1 net1661
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08123__C net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09912_ _05706_ _05730_ net319 _05853_ vssd1 vssd1 vccd1 vccd1 _05854_ sky130_fd_sc_hd__or4_1
XFILLER_0_1_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold179 net234 vssd1 vssd1 vccd1 vccd1 net1672 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout604 net605 vssd1 vssd1 vccd1 vccd1 net604 sky130_fd_sc_hd__buf_2
Xfanout615 net616 vssd1 vssd1 vccd1 vccd1 net615 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08546__A1 net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout626 net628 vssd1 vssd1 vccd1 vccd1 net626 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08546__B2 net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09843_ _05260_ _05262_ vssd1 vssd1 vccd1 vccd1 _05785_ sky130_fd_sc_hd__xnor2_1
Xfanout637 net638 vssd1 vssd1 vccd1 vccd1 net637 sky130_fd_sc_hd__clkbuf_4
Xfanout648 net659 vssd1 vssd1 vccd1 vccd1 net648 sky130_fd_sc_hd__buf_2
XANTENNA_fanout291_A net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout659 _06457_ vssd1 vssd1 vccd1 vccd1 net659 sky130_fd_sc_hd__clkbuf_8
XANTENNA__08641__S1 net1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07754__C1 net1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout389_A _06778_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13038__A net1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09774_ net666 _05715_ _03208_ _04646_ vssd1 vssd1 vccd1 vccd1 _05716_ sky130_fd_sc_hd__o2bb2a_1
X_06986_ _02822_ _02806_ _02801_ vssd1 vssd1 vccd1 vccd1 _02928_ sky130_fd_sc_hd__and3b_1
XANTENNA__11484__C _06550_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09950__S net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08725_ net928 _04666_ net1067 vssd1 vssd1 vccd1 vccd1 _04667_ sky130_fd_sc_hd__o21a_1
XANTENNA__07506__C1 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1298_A net1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08656_ _04596_ _04597_ net856 vssd1 vssd1 vccd1 vccd1 _04598_ sky130_fd_sc_hd__o21a_1
XFILLER_0_95_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_152_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07607_ net1204 team_03_WB.instance_to_wrap.core.register_file.registers_state\[729\]
+ net787 team_03_WB.instance_to_wrap.core.register_file.registers_state\[761\] net753
+ vssd1 vssd1 vccd1 vccd1 _03549_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_1_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08587_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[893\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[861\]
+ net966 vssd1 vssd1 vccd1 vccd1 _04529_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout344_X net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout723_A _02863_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1086_X net1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10408__A2 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07538_ _03476_ _03479_ net818 vssd1 vssd1 vccd1 vccd1 _03480_ sky130_fd_sc_hd__o21a_1
XANTENNA__08077__A3 net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_12_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11005__B net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07469_ net1116 _03409_ _03410_ vssd1 vssd1 vccd1 vccd1 _03411_ sky130_fd_sc_hd__or3_1
XANTENNA_fanout511_X net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1253_X net1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout609_X net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11720__S net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09208_ net608 _05147_ vssd1 vssd1 vccd1 vccd1 _05150_ sky130_fd_sc_hd__nor2_1
XFILLER_0_63_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10480_ net121 net1028 net906 net1677 vssd1 vssd1 vccd1 vccd1 _02629_ sky130_fd_sc_hd__a22o_1
XFILLER_0_106_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08154__X _04096_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09139_ net583 _05079_ vssd1 vssd1 vccd1 vccd1 _05081_ sky130_fd_sc_hd__nand2_1
XANTENNA__07037__A1 net1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10041__B1 net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08785__A1 net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12150_ net1579 vssd1 vssd1 vccd1 vccd1 _02403_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout880_X net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_442 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11101_ _06505_ net2658 net416 vssd1 vssd1 vccd1 vccd1 _02253_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout978_X net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07993__C1 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12081_ _06785_ net475 net441 net2123 vssd1 vssd1 vccd1 vccd1 _01466_ sky130_fd_sc_hd__a22o_1
XFILLER_0_130_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold680 team_03_WB.instance_to_wrap.core.register_file.registers_state\[274\] vssd1
+ vssd1 vccd1 vccd1 net2173 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_120_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold691 team_03_WB.instance_to_wrap.core.register_file.registers_state\[234\] vssd1
+ vssd1 vccd1 vccd1 net2184 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08537__A1 net1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11032_ net701 net712 net297 vssd1 vssd1 vccd1 vccd1 _06591_ sky130_fd_sc_hd__or3b_1
XANTENNA__11541__B1 net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_139_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12983_ net1392 vssd1 vssd1 vccd1 vccd1 _00747_ sky130_fd_sc_hd__inv_2
XFILLER_0_99_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_169_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14722_ clknet_leaf_46_wb_clk_i _02486_ _01087_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.decoder.inst\[19\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__08476__S net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11934_ net265 net2767 net369 vssd1 vssd1 vccd1 vccd1 _01608_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_178_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_178_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_14653_ clknet_leaf_166_wb_clk_i _02417_ _01018_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1007\]
+ sky130_fd_sc_hd__dfstp_1
X_11865_ net296 net1995 net378 vssd1 vssd1 vccd1 vccd1 _01675_ sky130_fd_sc_hd__mux2_1
XFILLER_0_169_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13604_ net1329 vssd1 vssd1 vccd1 vccd1 _01368_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_107_wb_clk_i clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_107_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_10816_ _06419_ _06420_ _06421_ vssd1 vssd1 vccd1 vccd1 _06422_ sky130_fd_sc_hd__o21ba_2
X_11796_ net2090 _06626_ net329 vssd1 vssd1 vccd1 vccd1 _01742_ sky130_fd_sc_hd__mux2_1
X_14584_ clknet_leaf_3_wb_clk_i _02348_ _00949_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[938\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_60_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07276__A1 net1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13535_ net1316 vssd1 vssd1 vccd1 vccd1 _01299_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10747_ team_03_WB.instance_to_wrap.core.pc.current_pc\[8\] _05718_ net604 vssd1
+ vssd1 vccd1 vccd1 _06366_ sky130_fd_sc_hd__mux2_1
XANTENNA__10594__X _06303_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_523 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13466_ net1340 vssd1 vssd1 vccd1 vccd1 _01230_ sky130_fd_sc_hd__inv_2
X_10678_ _02766_ _06319_ vssd1 vssd1 vccd1 vccd1 _06320_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_42_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07028__A1 net1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12021__A1 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12417_ net1290 vssd1 vssd1 vccd1 vccd1 _00181_ sky130_fd_sc_hd__inv_2
XFILLER_0_51_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13397_ net1431 vssd1 vssd1 vccd1 vccd1 _01161_ sky130_fd_sc_hd__inv_2
XFILLER_0_112_228 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07579__A2 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_874 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09973__A0 _03458_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10032__B1 net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput207 net207 vssd1 vssd1 vccd1 vccd1 gpio_out[10] sky130_fd_sc_hd__buf_2
XANTENNA__08776__A1 net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput218 net218 vssd1 vssd1 vccd1 vccd1 gpio_out[21] sky130_fd_sc_hd__buf_2
XFILLER_0_11_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput229 net229 vssd1 vssd1 vccd1 vccd1 gpio_out[32] sky130_fd_sc_hd__clkbuf_4
X_12348_ net1419 vssd1 vssd1 vccd1 vccd1 _00112_ sky130_fd_sc_hd__inv_2
XFILLER_0_65_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_178_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10583__B2 _02921_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_58_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15067_ net1453 vssd1 vssd1 vccd1 vccd1 la_data_out[3] sky130_fd_sc_hd__buf_2
XANTENNA__10770__A team_03_WB.instance_to_wrap.core.decoder.inst\[10\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12279_ net1386 vssd1 vssd1 vccd1 vccd1 _00043_ sky130_fd_sc_hd__inv_2
XFILLER_0_120_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08528__A1 net1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14018_ clknet_leaf_175_wb_clk_i _01782_ _00383_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[372\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10335__A1 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_147_3385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11077__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06840_ team_03_WB.instance_to_wrap.core.decoder.inst\[26\] vssd1 vssd1 vccd1 vccd1
+ _02783_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_147_3396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10886__A2 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11805__S net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08510_ net1227 team_03_WB.instance_to_wrap.core.register_file.registers_state\[607\]
+ net952 team_03_WB.instance_to_wrap.core.register_file.registers_state\[639\] net916
+ vssd1 vssd1 vccd1 vccd1 _04452_ sky130_fd_sc_hd__o221a_1
X_09490_ _05332_ _05430_ _05315_ _05324_ vssd1 vssd1 vccd1 vccd1 _05432_ sky130_fd_sc_hd__o211a_1
XANTENNA__08386__S net992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10929__B _05846_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07503__A2 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08441_ _04382_ vssd1 vssd1 vccd1 vccd1 _04383_ sky130_fd_sc_hd__inv_2
XFILLER_0_148_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_19_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_2857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_2868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08372_ net1049 team_03_WB.instance_to_wrap.core.register_file.registers_state\[662\]
+ net1000 team_03_WB.instance_to_wrap.core.register_file.registers_state\[694\] net920
+ vssd1 vssd1 vccd1 vccd1 _04314_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_173_3924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_173_3935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07323_ _03262_ _03264_ net812 vssd1 vssd1 vccd1 vccd1 _03265_ sky130_fd_sc_hd__a21o_1
XFILLER_0_45_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_143_320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07254_ net809 _03194_ _03195_ vssd1 vssd1 vccd1 vccd1 _03196_ sky130_fd_sc_hd__or3_1
XANTENNA__10810__A2 _05583_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08216__B1 net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07185_ net1084 team_03_WB.instance_to_wrap.core.register_file.registers_state\[659\]
+ net792 team_03_WB.instance_to_wrap.core.register_file.registers_state\[691\] vssd1
+ vssd1 vccd1 vccd1 _03127_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_30_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout304_A _05925_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08767__A1 net1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1046_A net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09964__A0 _05886_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10574__B2 _05884_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11771__B1 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1213_A team_03_WB.instance_to_wrap.core.decoder.inst\[17\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08519__A1 net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout401 _06718_ vssd1 vssd1 vccd1 vccd1 net401 sky130_fd_sc_hd__buf_4
Xfanout412 _06635_ vssd1 vssd1 vccd1 vccd1 net412 sky130_fd_sc_hd__buf_6
Xfanout423 _06560_ vssd1 vssd1 vccd1 vccd1 net423 sky130_fd_sc_hd__buf_4
Xfanout434 net437 vssd1 vssd1 vccd1 vccd1 net434 sky130_fd_sc_hd__buf_2
XANTENNA_fanout294_X net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout673_A net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_6_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout445 net446 vssd1 vssd1 vccd1 vccd1 net445 sky130_fd_sc_hd__buf_8
Xfanout456 net457 vssd1 vssd1 vccd1 vccd1 net456 sky130_fd_sc_hd__buf_2
X_09826_ _05764_ _05767_ _05758_ vssd1 vssd1 vccd1 vccd1 _05768_ sky130_fd_sc_hd__and3b_2
Xfanout467 net472 vssd1 vssd1 vccd1 vccd1 net467 sky130_fd_sc_hd__clkbuf_2
Xfanout478 net480 vssd1 vssd1 vccd1 vccd1 net478 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout1001_X net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout489 _06680_ vssd1 vssd1 vccd1 vccd1 net489 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09533__X _05475_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12079__A1 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout840_A net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09757_ _03243_ _04922_ net540 vssd1 vssd1 vccd1 vccd1 _05699_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout461_X net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06969_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[933\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[901\]
+ net787 vssd1 vssd1 vccd1 vccd1 _02911_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_5_wb_clk_i clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_5_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout938_A net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11715__S net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08708_ net557 _04649_ _04594_ vssd1 vssd1 vccd1 vccd1 _04650_ sky130_fd_sc_hd__o21ai_1
XANTENNA__08296__S net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09688_ net320 _05462_ _05467_ net322 _05629_ vssd1 vssd1 vccd1 vccd1 _05630_ sky130_fd_sc_hd__a221o_1
XFILLER_0_115_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08639_ net1054 team_03_WB.instance_to_wrap.core.register_file.registers_state\[966\]
+ net1007 team_03_WB.instance_to_wrap.core.register_file.registers_state\[998\] net1077
+ vssd1 vssd1 vccd1 vccd1 _04581_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_81_2031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout726_X net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1370_X net1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_2042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11650_ net2210 _06616_ net345 vssd1 vssd1 vccd1 vccd1 _01883_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10601_ net1751 team_03_WB.instance_to_wrap.CPU_DAT_O\[28\] net840 vssd1 vssd1 vccd1
+ vccd1 _02527_ sky130_fd_sc_hd__mux2_1
XANTENNA__07258__A1 net1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11054__A2 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11581_ net278 net2461 net448 vssd1 vssd1 vccd1 vccd1 _01948_ sky130_fd_sc_hd__mux2_1
XANTENNA__10855__A net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13231__A net1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10532_ net165 net1032 net1024 net1661 vssd1 vssd1 vccd1 vccd1 _02578_ sky130_fd_sc_hd__a22o_1
X_13320_ net1306 vssd1 vssd1 vccd1 vccd1 _01084_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08550__S0 net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_876 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10463_ _06134_ _06276_ vssd1 vssd1 vccd1 vccd1 _06277_ sky130_fd_sc_hd__nand2_1
XFILLER_0_122_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13251_ net1358 vssd1 vssd1 vccd1 vccd1 _01015_ sky130_fd_sc_hd__inv_2
XFILLER_0_33_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11389__C net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08044__B _03985_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12202_ net1618 vssd1 vssd1 vccd1 vccd1 _02351_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__09708__X _05650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13182_ net1410 vssd1 vssd1 vccd1 vccd1 _00946_ sky130_fd_sc_hd__inv_2
X_10394_ _06080_ _06081_ _06083_ vssd1 vssd1 vccd1 vccd1 _06221_ sky130_fd_sc_hd__and3_1
XANTENNA_input67_A wbs_adr_i[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11762__B1 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07966__C1 net1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12133_ net1544 vssd1 vssd1 vccd1 vccd1 _02420_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_102_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07430__A1 net1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09707__B1 net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07981__A2 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12064_ _06519_ net2717 net355 vssd1 vssd1 vccd1 vccd1 _01482_ sky130_fd_sc_hd__mux2_1
XANTENNA__11514__A0 net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08060__A net1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07718__C1 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11015_ net704 _06468_ net827 vssd1 vssd1 vccd1 vccd1 _06581_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_53_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10868__A2 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08930__A1 net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07733__A2 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout990 net994 vssd1 vssd1 vccd1 vccd1 net990 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_5_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_25 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_142_3282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_142_3293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12310__A net1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12966_ net1293 vssd1 vssd1 vccd1 vccd1 _00730_ sky130_fd_sc_hd__inv_2
XANTENNA__08143__C1 net1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10749__B net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14705_ clknet_leaf_33_wb_clk_i _02469_ _01070_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.control_logic.instruction\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_16_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11917_ _06618_ net2762 net368 vssd1 vssd1 vccd1 vccd1 _01625_ sky130_fd_sc_hd__mux2_1
XANTENNA__08694__B1 net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12897_ net1272 vssd1 vssd1 vccd1 vccd1 _00661_ sky130_fd_sc_hd__inv_2
XFILLER_0_68_760 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14636_ clknet_leaf_15_wb_clk_i _02400_ _01001_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[990\]
+ sky130_fd_sc_hd__dfstp_1
X_11848_ net278 net2085 net375 vssd1 vssd1 vccd1 vccd1 _01692_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_145_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11045__A2 net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14567_ clknet_leaf_97_wb_clk_i _02331_ _00932_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[921\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_32_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11779_ net2748 _06612_ net327 vssd1 vssd1 vccd1 vccd1 _01759_ sky130_fd_sc_hd__mux2_1
XANTENNA__10253__A0 _04235_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13518_ net1318 vssd1 vssd1 vccd1 vccd1 _01282_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14498_ clknet_leaf_177_wb_clk_i _02262_ _00863_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[852\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08235__A net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_1136 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload11 clknet_leaf_186_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload11/Y sky130_fd_sc_hd__clkinv_4
X_13449_ net1407 vssd1 vssd1 vccd1 vccd1 _01213_ sky130_fd_sc_hd__inv_2
Xclkload22 clknet_leaf_10_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload22/X sky130_fd_sc_hd__clkbuf_4
Xclkload33 clknet_leaf_179_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload33/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__11299__C net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_75_wb_clk_i clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_75_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__09097__S1 net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload44 clknet_leaf_24_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload44/Y sky130_fd_sc_hd__clkinv_2
XFILLER_0_140_334 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload55 clknet_leaf_15_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload55/Y sky130_fd_sc_hd__clkinv_2
XFILLER_0_51_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_1955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkload66 clknet_leaf_45_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload66/Y sky130_fd_sc_hd__inv_6
XFILLER_0_2_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkload77 clknet_leaf_57_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload77/Y sky130_fd_sc_hd__clkinv_2
XANTENNA__09410__A2 net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_1966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload88 clknet_leaf_70_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload88/Y sky130_fd_sc_hd__clkinv_4
XANTENNA__11753__B1 net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_149_3425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload99 clknet_leaf_146_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload99/Y sky130_fd_sc_hd__clkinv_1
X_15119_ net1488 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[24] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_149_3436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08990_ net1045 team_03_WB.instance_to_wrap.core.register_file.registers_state\[330\]
+ net995 team_03_WB.instance_to_wrap.core.register_file.registers_state\[362\] net1210
+ vssd1 vssd1 vccd1 vccd1 _04932_ sky130_fd_sc_hd__a221o_1
XANTENNA__09066__A net1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07941_ net822 _03876_ net720 vssd1 vssd1 vccd1 vccd1 _03883_ sky130_fd_sc_hd__o21ai_1
XANTENNA__11505__A0 _06623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_166_3783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07872_ net1200 team_03_WB.instance_to_wrap.core.register_file.registers_state\[219\]
+ net781 team_03_WB.instance_to_wrap.core.register_file.registers_state\[251\] net751
+ vssd1 vssd1 vccd1 vccd1 _03814_ sky130_fd_sc_hd__o221a_1
XANTENNA__07185__B1 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09611_ _03280_ _04532_ vssd1 vssd1 vccd1 vccd1 _05553_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_3_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06823_ team_03_WB.instance_to_wrap.core.pc.current_pc\[31\] vssd1 vssd1 vccd1 vccd1
+ _02766_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_123_2908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13316__A net1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09513__B _05453_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09542_ _05482_ _05483_ net565 vssd1 vssd1 vccd1 vccd1 _05484_ sky130_fd_sc_hd__mux2_1
XANTENNA__09005__S net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09473_ _05413_ _05414_ net553 vssd1 vssd1 vccd1 vccd1 _05415_ sky130_fd_sc_hd__mux2_1
XANTENNA__11284__A2 net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11481__D net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10492__B1 net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08424_ net1063 _04363_ _04364_ vssd1 vssd1 vccd1 vccd1 _04366_ sky130_fd_sc_hd__or3_1
XFILLER_0_136_607 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08355_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[54\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[22\]
+ net972 vssd1 vssd1 vccd1 vccd1 _04297_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout421_A _06560_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1163_A net1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07306_ net1185 team_03_WB.instance_to_wrap.core.register_file.registers_state\[605\]
+ net768 team_03_WB.instance_to_wrap.core.register_file.registers_state\[637\] net728
+ vssd1 vssd1 vccd1 vccd1 _03248_ sky130_fd_sc_hd__o221a_1
XANTENNA__13051__A net1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout519_A _06395_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload5 clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload5/Y sky130_fd_sc_hd__clkinv_8
XFILLER_0_11_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08286_ _04224_ _04225_ _04226_ _04227_ net861 net920 vssd1 vssd1 vccd1 vccd1 _04228_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_116_342 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_876 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11992__A0 net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07237_ net1131 _03172_ _03173_ net1139 vssd1 vssd1 vccd1 vccd1 _03179_ sky130_fd_sc_hd__a31o_1
XFILLER_0_131_301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1330_A net1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout307_X net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1049_X net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07984__A net1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07168_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[51\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[19\]
+ net763 vssd1 vssd1 vccd1 vccd1 _03110_ sky130_fd_sc_hd__mux2_1
XANTENNA__07099__S0 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout790_A _02851_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11744__B1 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08799__B net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout888_A net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07099_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[929\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[897\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[801\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[769\]
+ net780 net1134 vssd1 vssd1 vccd1 vccd1 _03041_ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout1216_X net1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07195__S net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07963__A2 net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1207 net1209 vssd1 vssd1 vccd1 vccd1 net1207 sky130_fd_sc_hd__buf_6
XFILLER_0_79_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1218 net1225 vssd1 vssd1 vccd1 vccd1 net1218 sky130_fd_sc_hd__buf_4
XFILLER_0_121_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1229 net1238 vssd1 vssd1 vccd1 vccd1 net1229 sky130_fd_sc_hd__clkbuf_2
Xfanout264 _06537_ vssd1 vssd1 vccd1 vccd1 net264 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_31_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout275 _06446_ vssd1 vssd1 vccd1 vccd1 net275 sky130_fd_sc_hd__buf_2
XANTENNA__08373__C1 net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout286 _05946_ vssd1 vssd1 vccd1 vccd1 net286 sky130_fd_sc_hd__buf_4
X_09809_ _02923_ _04565_ net667 _05750_ vssd1 vssd1 vccd1 vccd1 _05751_ sky130_fd_sc_hd__a22o_1
Xfanout297 _06499_ vssd1 vssd1 vccd1 vccd1 net297 sky130_fd_sc_hd__buf_2
XANTENNA_fanout843_X net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1041 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12820_ net1313 vssd1 vssd1 vccd1 vccd1 _00584_ sky130_fd_sc_hd__inv_2
XFILLER_0_69_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12751_ net1337 vssd1 vssd1 vccd1 vccd1 _00515_ sky130_fd_sc_hd__inv_2
XANTENNA__11391__D net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_1084 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10483__B1 net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11702_ _06744_ net384 net340 net1999 vssd1 vssd1 vccd1 vccd1 _01832_ sky130_fd_sc_hd__a22o_1
XFILLER_0_96_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12682_ net1279 vssd1 vssd1 vccd1 vccd1 _00446_ sky130_fd_sc_hd__inv_2
XFILLER_0_166_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14421_ clknet_leaf_114_wb_clk_i _02185_ _00786_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[775\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_108_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08428__B1 net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11633_ _06707_ net385 net349 net2277 vssd1 vssd1 vccd1 vccd1 _01899_ sky130_fd_sc_hd__a22o_1
XFILLER_0_166_286 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08979__A1 net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14352_ clknet_leaf_156_wb_clk_i _02116_ _00717_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[706\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07597__C net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11564_ net2325 net484 _06796_ net508 vssd1 vssd1 vccd1 vccd1 _01960_ sky130_fd_sc_hd__a22o_1
XANTENNA__11983__A0 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13303_ net1321 vssd1 vssd1 vccd1 vccd1 _01067_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_98_2380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10515_ net152 net1032 net1024 net1716 vssd1 vssd1 vccd1 vccd1 _02595_ sky130_fd_sc_hd__a22o_1
XANTENNA__07651__A1 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_2391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14283_ clknet_leaf_42_wb_clk_i _02047_ _00648_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[637\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11495_ _06616_ net2608 net391 vssd1 vssd1 vccd1 vccd1 _02011_ sky130_fd_sc_hd__mux2_1
XFILLER_0_162_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09928__A0 _05868_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_811 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10446_ _06032_ _06055_ vssd1 vssd1 vccd1 vccd1 _06263_ sky130_fd_sc_hd__xor2_1
X_13234_ net1398 vssd1 vssd1 vccd1 vccd1 _00998_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_1056 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07939__C1 net1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_2299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_855 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07403__A1 net1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10377_ _05986_ _05987_ _06087_ vssd1 vssd1 vccd1 vccd1 _06207_ sky130_fd_sc_hd__or3_1
XFILLER_0_21_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13165_ net1276 vssd1 vssd1 vccd1 vccd1 _00929_ sky130_fd_sc_hd__inv_2
XANTENNA__12305__A net1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12116_ _02776_ team_03_WB.instance_to_wrap.READ_I team_03_WB.instance_to_wrap.wb.curr_state\[0\]
+ _02797_ net2774 vssd1 vssd1 vccd1 vccd1 _00008_ sky130_fd_sc_hd__a32o_1
X_13096_ net1297 vssd1 vssd1 vccd1 vccd1 _00860_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_72_1852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_3322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12047_ _06616_ net2605 net358 vssd1 vssd1 vccd1 vccd1 _01499_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_144_3333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07833__S net1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_68 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10710__A1 net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_161_3680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_122_wb_clk_i clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_122_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_1_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12040__A net1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13998_ clknet_leaf_128_wb_clk_i _01762_ _00363_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[352\]
+ sky130_fd_sc_hd__dfrtp_1
X_12949_ net1275 vssd1 vssd1 vccd1 vccd1 _00713_ sky130_fd_sc_hd__inv_2
XANTENNA__11266__A2 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08667__B1 net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_146_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11018__A2 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_315 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14619_ clknet_leaf_120_wb_clk_i _02383_ _00984_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[973\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__07890__A1 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11090__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08140_ net1207 _02820_ vssd1 vssd1 vccd1 vccd1 _04082_ sky130_fd_sc_hd__nand2_1
XFILLER_0_16_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_wire591_A _04861_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09631__A2 _04415_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07642__A1 net1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload100 clknet_leaf_147_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload100/Y sky130_fd_sc_hd__clkinv_4
X_08071_ net1183 team_03_WB.instance_to_wrap.core.register_file.registers_state\[566\]
+ net876 vssd1 vssd1 vccd1 vccd1 _04013_ sky130_fd_sc_hd__and3_1
Xclkload111 clknet_leaf_118_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload111/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_3_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload122 clknet_leaf_135_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload122/X sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_116_2756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_2767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07022_ net1196 net883 team_03_WB.instance_to_wrap.core.register_file.registers_state\[643\]
+ vssd1 vssd1 vccd1 vccd1 _02964_ sky130_fd_sc_hd__a21o_1
Xclkload133 clknet_leaf_123_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload133/Y sky130_fd_sc_hd__inv_6
Xclkload144 clknet_leaf_78_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload144/X sky130_fd_sc_hd__clkbuf_8
Xclkload155 clknet_leaf_85_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload155/Y sky130_fd_sc_hd__clkinv_2
XFILLER_0_114_879 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload166 clknet_leaf_126_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload166/Y sky130_fd_sc_hd__bufinv_16
XTAP_TAPCELL_ROW_168_3823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload177 clknet_leaf_93_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload177/Y sky130_fd_sc_hd__inv_8
XTAP_TAPCELL_ROW_168_3834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_343 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08973_ net1209 _04911_ _04914_ net853 vssd1 vssd1 vccd1 vccd1 _04915_ sky130_fd_sc_hd__o31a_1
Xhold17 team_03_WB.instance_to_wrap.core.register_file.registers_state\[937\] vssd1
+ vssd1 vccd1 vccd1 net1510 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_46_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07924_ net613 _03864_ _03865_ vssd1 vssd1 vccd1 vccd1 _03866_ sky130_fd_sc_hd__o21a_2
Xhold28 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1011\] vssd1
+ vssd1 vccd1 vccd1 net1521 sky130_fd_sc_hd__dlygate4sd3_1
Xhold39 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1021\] vssd1
+ vssd1 vccd1 vccd1 net1532 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1009_A net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07855_ net1120 _03795_ _03796_ net1136 vssd1 vssd1 vccd1 vccd1 _03797_ sky130_fd_sc_hd__a211o_1
XANTENNA__10701__A1 _06316_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout371_A _06813_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout469_A net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07786_ _03680_ _03681_ _03725_ _03726_ vssd1 vssd1 vccd1 vccd1 _03728_ sky130_fd_sc_hd__o22a_1
XFILLER_0_78_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07044__A net1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09525_ _05464_ _05465_ net567 vssd1 vssd1 vccd1 vccd1 _05467_ sky130_fd_sc_hd__mux2_1
XANTENNA__08658__B1 net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1280_A net1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12885__A net1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout636_A net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1378_A net1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08122__A2 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_376 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_3_5_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_5_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_66_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09456_ net552 _04080_ _04770_ _05135_ vssd1 vssd1 vccd1 vccd1 _05398_ sky130_fd_sc_hd__o31ai_1
XANTENNA__06883__A team_03_WB.instance_to_wrap.core.decoder.inst\[28\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08407_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[953\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[921\]
+ net991 vssd1 vssd1 vccd1 vccd1 _04349_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout424_X net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09387_ _05327_ _05328_ vssd1 vssd1 vccd1 vccd1 _05329_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout803_A net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1166_X net1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08338_ _04274_ _04279_ net872 vssd1 vssd1 vccd1 vccd1 _04280_ sky130_fd_sc_hd__mux2_1
XANTENNA__11965__B1 net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_824 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07094__C1 net1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07633__A1 net1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11013__B net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08269_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[55\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[23\]
+ net964 vssd1 vssd1 vccd1 vccd1 _04211_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10300_ team_03_WB.instance_to_wrap.core.pc.current_pc\[15\] team_03_WB.instance_to_wrap.core.pc.current_pc\[14\]
+ _06141_ vssd1 vssd1 vccd1 vccd1 _06142_ sky130_fd_sc_hd__and3_1
XFILLER_0_160_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11280_ net512 net644 _06707_ net411 net2475 vssd1 vssd1 vccd1 vccd1 _02155_ sky130_fd_sc_hd__a32o_1
XFILLER_0_15_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout793_X net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10231_ _03864_ _06071_ _06072_ vssd1 vssd1 vccd1 vccd1 _06073_ sky130_fd_sc_hd__and3_1
XFILLER_0_113_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11193__A1 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10162_ _06003_ vssd1 vssd1 vccd1 vccd1 _06004_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_7_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout960_X net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07492__S0 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1004 net1005 vssd1 vssd1 vccd1 vccd1 net1004 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10940__A1 team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[6\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1015 _02821_ vssd1 vssd1 vccd1 vccd1 net1015 sky130_fd_sc_hd__buf_4
XFILLER_0_100_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1026 _06286_ vssd1 vssd1 vccd1 vccd1 net1026 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_50_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1037 net1038 vssd1 vssd1 vccd1 vccd1 net1037 sky130_fd_sc_hd__clkbuf_2
X_14970_ clknet_leaf_94_wb_clk_i _02722_ _01335_ vssd1 vssd1 vccd1 vccd1 net222 sky130_fd_sc_hd__dfrtp_1
X_10093_ _05611_ _05676_ _05811_ _05931_ vssd1 vssd1 vccd1 vccd1 _05937_ sky130_fd_sc_hd__and4bb_1
XTAP_TAPCELL_ROW_50_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1048 net1049 vssd1 vssd1 vccd1 vccd1 net1048 sky130_fd_sc_hd__buf_2
Xfanout1059 net1060 vssd1 vssd1 vccd1 vccd1 net1059 sky130_fd_sc_hd__buf_4
XANTENNA__08346__C1 net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_156_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13921_ clknet_leaf_174_wb_clk_i _01685_ _00286_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[275\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08897__B1 net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1135 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08992__S0 net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13852_ clknet_leaf_149_wb_clk_i _01616_ _00217_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[206\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_16_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12803_ net1354 vssd1 vssd1 vccd1 vccd1 _00567_ sky130_fd_sc_hd__inv_2
XANTENNA__11248__A2 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13783_ clknet_leaf_113_wb_clk_i _01547_ _00148_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[137\]
+ sky130_fd_sc_hd__dfrtp_1
X_10995_ net491 net647 _06569_ net420 net2104 vssd1 vssd1 vccd1 vccd1 _02302_ sky130_fd_sc_hd__a32o_1
XFILLER_0_85_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_48_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12734_ net1392 vssd1 vssd1 vccd1 vccd1 _00498_ sky130_fd_sc_hd__inv_2
XANTENNA__08484__S net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_184 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09614__A1_N team_03_WB.instance_to_wrap.core.decoder.inst\[29\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1060 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07872__A1 net1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12665_ net1365 vssd1 vssd1 vccd1 vccd1 _00429_ sky130_fd_sc_hd__inv_2
XFILLER_0_84_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14404_ clknet_leaf_29_wb_clk_i _02168_ _00769_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[758\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_936 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11616_ _06690_ net381 net347 net2251 vssd1 vssd1 vccd1 vccd1 _01916_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_137_3181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09613__A2 _04532_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12596_ net1304 vssd1 vssd1 vccd1 vccd1 _00360_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_137_3192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11956__B1 net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_2339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14335_ clknet_leaf_171_wb_clk_i _02099_ _00700_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[689\]
+ sky130_fd_sc_hd__dfrtp_1
X_11547_ net630 _06657_ vssd1 vssd1 vccd1 vccd1 _06789_ sky130_fd_sc_hd__and2_1
XFILLER_0_41_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold509 team_03_WB.instance_to_wrap.core.register_file.registers_state\[685\] vssd1
+ vssd1 vccd1 vccd1 net2002 sky130_fd_sc_hd__dlygate4sd3_1
X_14266_ clknet_leaf_142_wb_clk_i _02030_ _00631_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[620\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11971__A3 net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08513__A net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11478_ net2638 net393 _06774_ net509 vssd1 vssd1 vccd1 vccd1 _02024_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_74_1903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10762__B _06294_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11708__B1 net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_698 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13217_ net1260 vssd1 vssd1 vccd1 vccd1 _00981_ sky130_fd_sc_hd__inv_2
X_10429_ _06248_ _06249_ team_03_WB.instance_to_wrap.core.pc.current_pc\[10\] net682
+ vssd1 vssd1 vccd1 vccd1 _02644_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_122_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14197_ clknet_leaf_107_wb_clk_i _01961_ _00562_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[551\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_111_2653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07927__A2 net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_2664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11723__A3 net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_23 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07129__A net1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13148_ net1419 vssd1 vssd1 vccd1 vccd1 _00912_ sky130_fd_sc_hd__inv_2
XFILLER_0_20_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_163_3720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_163_3731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13079_ net1391 vssd1 vssd1 vccd1 vccd1 _00843_ sky130_fd_sc_hd__inv_2
XFILLER_0_40_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1209 team_03_WB.instance_to_wrap.core.register_file.registers_state\[81\] vssd1
+ vssd1 vccd1 vccd1 net2702 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_174_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11487__A2 net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_164_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11085__S net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07155__A3 net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07640_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[430\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[398\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[302\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[270\]
+ net777 net1131 vssd1 vssd1 vccd1 vccd1 _03582_ sky130_fd_sc_hd__mux4_1
XANTENNA__07560__B1 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07571_ net750 _03511_ _03512_ net1167 vssd1 vssd1 vccd1 vccd1 _03513_ sky130_fd_sc_hd__a31o_1
X_09310_ net583 _05251_ vssd1 vssd1 vccd1 vccd1 _05252_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_76_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07312__B1 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10998__B2 net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09241_ _05176_ _05182_ _05177_ vssd1 vssd1 vccd1 vccd1 _05183_ sky130_fd_sc_hd__or3b_1
XFILLER_0_29_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_145_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_560 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_90_wb_clk_i clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_90_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_118_2807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09172_ _05110_ _05113_ net555 vssd1 vssd1 vccd1 vccd1 _05114_ sky130_fd_sc_hd__mux2_1
XANTENNA__09065__B1 net999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11947__B1 net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08123_ net1087 team_03_WB.instance_to_wrap.core.register_file.registers_state\[954\]
+ net892 vssd1 vssd1 vccd1 vccd1 _04065_ sky130_fd_sc_hd__or3_1
XFILLER_0_161_749 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08812__B1 net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08054_ net1188 team_03_WB.instance_to_wrap.core.register_file.registers_state\[86\]
+ net771 team_03_WB.instance_to_wrap.core.register_file.registers_state\[118\] net738
+ vssd1 vssd1 vccd1 vccd1 _03996_ sky130_fd_sc_hd__o221a_1
XFILLER_0_142_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11962__A3 net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07005_ _02945_ _02946_ vssd1 vssd1 vccd1 vccd1 _02947_ sky130_fd_sc_hd__and2b_1
XFILLER_0_3_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_838 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_674 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1126_A net1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07039__A net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08040__A1 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold1234_A team_03_WB.instance_to_wrap.core.register_file.registers_state\[9\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08956_ net945 _04896_ _04897_ vssd1 vssd1 vccd1 vccd1 _04898_ sky130_fd_sc_hd__o21a_1
XFILLER_0_138_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07907_ net1187 team_03_WB.instance_to_wrap.core.register_file.registers_state\[687\]
+ net877 vssd1 vssd1 vccd1 vccd1 _03849_ sky130_fd_sc_hd__and3_1
XANTENNA__11478__A2 net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08887_ net565 _04827_ vssd1 vssd1 vccd1 vccd1 _04829_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout753_A net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout374_X net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07146__A3 net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07838_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[938\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[906\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[810\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[778\]
+ net760 net1127 vssd1 vssd1 vccd1 vccd1 _03780_ sky130_fd_sc_hd__mux4_1
XANTENNA__07551__B1 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout920_A net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11008__B net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07769_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[908\] net796
+ _03703_ net1118 vssd1 vssd1 vccd1 vccd1 _03711_ sky130_fd_sc_hd__o211a_1
XFILLER_0_6_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1283_X net1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout639_X net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09508_ net573 _05449_ vssd1 vssd1 vccd1 vccd1 _05450_ sky130_fd_sc_hd__or2_1
XANTENNA__07529__S1 net1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10780_ _06389_ _06380_ vssd1 vssd1 vccd1 vccd1 _06390_ sky130_fd_sc_hd__and2b_2
XFILLER_0_39_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07502__A net1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09439_ _05379_ _05380_ net557 vssd1 vssd1 vccd1 vccd1 _05381_ sky130_fd_sc_hd__mux2_1
XANTENNA__07854__A1 net1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout806_X net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_519 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11024__A net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07221__B net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12450_ net1359 vssd1 vssd1 vccd1 vccd1 _00214_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_43_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_576 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11938__A0 net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_738 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11401_ _06413_ net2576 net397 vssd1 vssd1 vccd1 vccd1 _02079_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08803__B1 net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12381_ net1383 vssd1 vssd1 vccd1 vccd1 _00145_ sky130_fd_sc_hd__inv_2
XFILLER_0_151_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09071__A3 net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07648__S net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14120_ clknet_leaf_8_wb_clk_i _01884_ _00485_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[474\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09429__A net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11953__A3 net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11332_ net1042 _06449_ net650 net694 vssd1 vssd1 vccd1 vccd1 _06718_ sky130_fd_sc_hd__or4_4
XFILLER_0_132_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07082__A2 _03023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_160_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_91_2236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14051_ clknet_leaf_30_wb_clk_i _01815_ _00416_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[405\]
+ sky130_fd_sc_hd__dfrtp_1
X_11263_ net1249 net838 _06477_ net671 vssd1 vssd1 vccd1 vccd1 _06699_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_91_2247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_45_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11166__B2 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08567__C1 net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13002_ net1286 vssd1 vssd1 vccd1 vccd1 _00766_ sky130_fd_sc_hd__inv_2
X_10214_ _06032_ _06055_ _06030_ vssd1 vssd1 vccd1 vccd1 _06056_ sky130_fd_sc_hd__o21ai_1
X_11194_ net655 net705 net267 net697 vssd1 vssd1 vccd1 vccd1 _06678_ sky130_fd_sc_hd__and4_1
XANTENNA__10913__A1 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10145_ _03109_ _05985_ vssd1 vssd1 vccd1 vccd1 _05987_ sky130_fd_sc_hd__nor2_1
XFILLER_0_27_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08319__C1 net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10076_ _05342_ net314 _05919_ net581 _02937_ vssd1 vssd1 vccd1 vccd1 _05920_ sky130_fd_sc_hd__o2111a_1
X_14953_ clknet_leaf_95_wb_clk_i _02705_ _01318_ vssd1 vssd1 vccd1 vccd1 net236 sky130_fd_sc_hd__dfrtp_1
XANTENNA__11469__A2 net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13904_ clknet_leaf_160_wb_clk_i _01668_ _00269_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[258\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_89_2198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14884_ clknet_leaf_67_wb_clk_i _02647_ _01249_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.pc.current_pc\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_159_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13835_ clknet_leaf_34_wb_clk_i _01599_ _00200_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[189\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_159_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_600 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09611__B _04532_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_139_3221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09295__B1 net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13766_ clknet_leaf_73_wb_clk_i _01530_ _00131_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[120\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_174_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_139_3232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10978_ _06551_ _06554_ _06556_ _06391_ vssd1 vssd1 vccd1 vccd1 _06557_ sky130_fd_sc_hd__o211a_4
XFILLER_0_70_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09834__A2 _05436_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07412__A net1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12717_ net1331 vssd1 vssd1 vccd1 vccd1 _00481_ sky130_fd_sc_hd__inv_2
XANTENNA__11641__A2 net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13697_ clknet_leaf_181_wb_clk_i _01461_ _00062_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[51\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12648_ net1297 vssd1 vssd1 vccd1 vccd1 _00412_ sky130_fd_sc_hd__inv_2
XANTENNA__09047__B1 net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11929__A0 _06505_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_84_wb_clk_i_A clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_170_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_154_Left_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_749 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_535 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12579_ net1374 vssd1 vssd1 vccd1 vccd1 _00343_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_152_3487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_152_3498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_2704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14318_ clknet_leaf_124_wb_clk_i _02082_ _00683_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[672\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_382 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11944__A3 net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold306 team_03_WB.instance_to_wrap.core.register_file.registers_state\[683\] vssd1
+ vssd1 vccd1 vccd1 net1799 sky130_fd_sc_hd__dlygate4sd3_1
Xhold317 _02517_ vssd1 vssd1 vccd1 vccd1 net1810 sky130_fd_sc_hd__dlygate4sd3_1
Xhold328 team_03_WB.instance_to_wrap.CPU_DAT_I\[12\] vssd1 vssd1 vccd1 vccd1 net1821
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold339 team_03_WB.instance_to_wrap.core.register_file.registers_state\[549\] vssd1
+ vssd1 vccd1 vccd1 net1832 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14249_ clknet_leaf_117_wb_clk_i _02013_ _00614_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[603\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_68 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout808 net810 vssd1 vssd1 vccd1 vccd1 net808 sky130_fd_sc_hd__buf_4
Xfanout819 net820 vssd1 vssd1 vccd1 vccd1 net819 sky130_fd_sc_hd__clkbuf_8
XANTENNA__09770__A1 net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08810_ net1221 _04749_ _04750_ vssd1 vssd1 vccd1 vccd1 _04752_ sky130_fd_sc_hd__and3_1
XANTENNA__11808__S net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09770__B2 net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09790_ _05246_ _05250_ _05269_ net595 vssd1 vssd1 vccd1 vccd1 _05732_ sky130_fd_sc_hd__a31o_1
XFILLER_0_84_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1006 team_03_WB.instance_to_wrap.core.register_file.registers_state\[39\] vssd1
+ vssd1 vccd1 vccd1 net2499 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_163_Left_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1017 team_03_WB.instance_to_wrap.core.register_file.registers_state\[544\] vssd1
+ vssd1 vccd1 vccd1 net2510 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_84_32 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08741_ net1239 team_03_WB.instance_to_wrap.core.register_file.registers_state\[131\]
+ net980 team_03_WB.instance_to_wrap.core.register_file.registers_state\[163\] net942
+ vssd1 vssd1 vccd1 vccd1 _04683_ sky130_fd_sc_hd__o221a_1
Xhold1028 team_03_WB.instance_to_wrap.core.register_file.registers_state\[657\] vssd1
+ vssd1 vccd1 vccd1 net2521 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1039 team_03_WB.instance_to_wrap.core.register_file.registers_state\[536\] vssd1
+ vssd1 vccd1 vccd1 net2532 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_139_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1390 net1392 vssd1 vssd1 vccd1 vccd1 net1390 sky130_fd_sc_hd__buf_4
XFILLER_0_139_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08672_ net930 _04612_ _04613_ vssd1 vssd1 vccd1 vccd1 _04614_ sky130_fd_sc_hd__a21o_1
XANTENNA__07533__B1 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07623_ _03278_ _03564_ vssd1 vssd1 vccd1 vccd1 _03565_ sky130_fd_sc_hd__and2b_1
XPHY_EDGE_ROW_5_Right_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07554_ _03493_ _03495_ net812 vssd1 vssd1 vccd1 vccd1 _03496_ sky130_fd_sc_hd__a21o_1
X_07485_ _03426_ vssd1 vssd1 vccd1 vccd1 _03427_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07836__A1 net1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11632__A2 net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout334_A _06809_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1076_A net1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09948__S net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_172_Left_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09224_ _05164_ _05165_ vssd1 vssd1 vccd1 vccd1 _05166_ sky130_fd_sc_hd__nor2_1
XFILLER_0_63_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_173_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09155_ net432 net425 _04267_ net547 vssd1 vssd1 vccd1 vccd1 _05097_ sky130_fd_sc_hd__o31a_1
XFILLER_0_16_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout501_A net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1243_A net1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11396__A1 net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_287 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08106_ net1087 team_03_WB.instance_to_wrap.core.register_file.registers_state\[634\]
+ net892 vssd1 vssd1 vccd1 vccd1 _04048_ sky130_fd_sc_hd__or3_1
XANTENNA__09249__A _04294_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09086_ net1240 team_03_WB.instance_to_wrap.core.register_file.registers_state\[589\]
+ net982 team_03_WB.instance_to_wrap.core.register_file.registers_state\[621\] net927
+ vssd1 vssd1 vccd1 vccd1 _05028_ sky130_fd_sc_hd__o221a_1
XFILLER_0_71_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_142_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08037_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[401\] net792
+ _03978_ vssd1 vssd1 vccd1 vccd1 _03979_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout1031_X net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1069 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1410_A net1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold840 team_03_WB.instance_to_wrap.core.register_file.registers_state\[590\] vssd1
+ vssd1 vccd1 vccd1 net2333 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_31_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08549__C1 net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1129_X net1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold851 team_03_WB.instance_to_wrap.core.register_file.registers_state\[807\] vssd1
+ vssd1 vccd1 vccd1 net2344 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12106__C _06293_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold862 team_03_WB.instance_to_wrap.core.register_file.registers_state\[762\] vssd1
+ vssd1 vccd1 vccd1 net2355 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08013__A1 net1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold873 team_03_WB.instance_to_wrap.core.register_file.registers_state\[514\] vssd1
+ vssd1 vccd1 vccd1 net2366 sky130_fd_sc_hd__dlygate4sd3_1
Xhold884 team_03_WB.instance_to_wrap.core.register_file.registers_state\[863\] vssd1
+ vssd1 vccd1 vccd1 net2377 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08440__X _04382_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11699__A2 net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout491_X net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold895 team_03_WB.instance_to_wrap.core.register_file.registers_state\[112\] vssd1
+ vssd1 vccd1 vccd1 net2388 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout968_A net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11718__S net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10622__S net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09988_ _05873_ net1769 net288 vssd1 vssd1 vccd1 vccd1 _02726_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_129_wb_clk_i_A clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_15095__1481 vssd1 vssd1 vccd1 vccd1 _15095__1481/HI net1481 sky130_fd_sc_hd__conb_1
XANTENNA__10108__C1 _03060_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08939_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[811\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[779\]
+ net961 vssd1 vssd1 vccd1 vccd1 _04881_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_150_Right_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08316__A2 net999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11019__A net1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11950_ net628 _06727_ net460 net364 net2539 vssd1 vssd1 vccd1 vccd1 _01593_ sky130_fd_sc_hd__a32o_1
XANTENNA__06895__X _02837_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09712__A net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10901_ net313 net309 net316 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[13\]
+ vssd1 vssd1 vccd1 vccd1 _06493_ sky130_fd_sc_hd__o31a_1
XFILLER_0_54_1127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11881_ net619 _06690_ net452 net372 net2199 vssd1 vssd1 vccd1 vccd1 _01660_ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout923_X net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13620_ net1425 vssd1 vssd1 vccd1 vccd1 _01384_ sky130_fd_sc_hd__inv_2
XANTENNA__13234__A net1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10832_ _06434_ net2464 net518 vssd1 vssd1 vccd1 vccd1 _02330_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_45_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_167 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_2095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07232__A net1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13551_ net1420 vssd1 vssd1 vccd1 vccd1 _01315_ sky130_fd_sc_hd__inv_2
XANTENNA__07288__C1 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10763_ _05798_ net604 vssd1 vssd1 vccd1 vccd1 _06376_ sky130_fd_sc_hd__nand2_1
XANTENNA__11623__A2 net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_165_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10296__C _06136_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12502_ net1258 vssd1 vssd1 vccd1 vccd1 _00266_ sky130_fd_sc_hd__inv_2
XFILLER_0_82_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10831__B1 _06401_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09029__B1 net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13482_ net1405 vssd1 vssd1 vccd1 vccd1 _01246_ sky130_fd_sc_hd__inv_2
XANTENNA__08762__S net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input97_A wbs_adr_i[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10694_ team_03_WB.instance_to_wrap.core.pc.current_pc\[28\] _06316_ net602 vssd1
+ vssd1 vccd1 vccd1 _06333_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_124_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_152_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12433_ net1271 vssd1 vssd1 vccd1 vccd1 _00197_ sky130_fd_sc_hd__inv_2
XFILLER_0_63_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12364_ net1313 vssd1 vssd1 vccd1 vccd1 _00128_ sky130_fd_sc_hd__inv_2
XANTENNA__08252__A1 net1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_1_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_3037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_544 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_130_3048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14103_ clknet_leaf_112_wb_clk_i _01867_ _00468_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[457\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_168_wb_clk_i_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_11315_ _06622_ net2642 net407 vssd1 vssd1 vccd1 vccd1 _02130_ sky130_fd_sc_hd__mux2_1
X_15083_ net1469 vssd1 vssd1 vccd1 vccd1 la_data_out[19] sky130_fd_sc_hd__buf_2
XANTENNA__07460__C1 net1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12295_ net1368 vssd1 vssd1 vccd1 vccd1 _00059_ sky130_fd_sc_hd__inv_2
XANTENNA__11139__B2 net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09446__X _05388_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14034_ clknet_leaf_165_wb_clk_i _01798_ _00399_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[388\]
+ sky130_fd_sc_hd__dfrtp_1
X_11246_ net497 net626 _06690_ net409 net2355 vssd1 vssd1 vccd1 vccd1 _02172_ sky130_fd_sc_hd__a32o_1
XANTENNA__07212__C1 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11177_ net2219 net415 _06668_ net512 vssd1 vssd1 vccd1 vccd1 _02219_ sky130_fd_sc_hd__a22o_1
XFILLER_0_59_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10128_ _05966_ _05967_ _03279_ vssd1 vssd1 vccd1 vccd1 _05970_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_59_1027 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12103__A3 net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14936_ clknet_leaf_52_wb_clk_i _02691_ _01301_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_O\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_10059_ net28 net1037 net910 net2772 vssd1 vssd1 vccd1 vccd1 _02672_ sky130_fd_sc_hd__o22a_1
XANTENNA__08937__S net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07515__B1 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_171_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_29_wb_clk_i clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_29_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_106_2552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14867_ clknet_leaf_59_wb_clk_i net1641 _01232_ vssd1 vssd1 vccd1 vccd1 net123 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_106_2563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10768__A _05142_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_159_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13818_ clknet_leaf_144_wb_clk_i _01582_ _00183_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[172\]
+ sky130_fd_sc_hd__dfrtp_1
X_14798_ clknet_leaf_89_wb_clk_i _02562_ _01163_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_I\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07142__A net1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07279__C1 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_666 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11614__A2 net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13749_ clknet_leaf_105_wb_clk_i _01513_ _00114_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[103\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_154_3527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10822__A0 net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_154_3538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09768__S net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07270_ net1112 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1001\]
+ net902 _03211_ net1158 vssd1 vssd1 vccd1 vccd1 _03212_ sky130_fd_sc_hd__o311a_1
XFILLER_0_73_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08491__A1 net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_171_822 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_171_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_171_3885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11378__A1 net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08779__C1 net1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08243__A1 net1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold103 _02594_ vssd1 vssd1 vccd1 vccd1 net1596 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10050__A1 net6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold114 team_03_WB.instance_to_wrap.core.register_file.registers_state\[30\] vssd1
+ vssd1 vccd1 vccd1 net1607 sky130_fd_sc_hd__dlygate4sd3_1
Xhold125 team_03_WB.instance_to_wrap.core.register_file.registers_state\[941\] vssd1
+ vssd1 vccd1 vccd1 net1618 sky130_fd_sc_hd__dlygate4sd3_1
Xhold136 _02626_ vssd1 vssd1 vccd1 vccd1 net1629 sky130_fd_sc_hd__dlygate4sd3_1
Xhold147 team_03_WB.instance_to_wrap.ADR_I\[28\] vssd1 vssd1 vccd1 vccd1 net1640 sky130_fd_sc_hd__dlygate4sd3_1
Xhold158 team_03_WB.instance_to_wrap.core.register_file.registers_state\[31\] vssd1
+ vssd1 vccd1 vccd1 net1651 sky130_fd_sc_hd__dlygate4sd3_1
X_09911_ _05757_ _05769_ vssd1 vssd1 vccd1 vccd1 _05853_ sky130_fd_sc_hd__nand2_1
XFILLER_0_111_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold169 _02578_ vssd1 vssd1 vccd1 vccd1 net1662 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10950__B net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08701__A net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout605 _06295_ vssd1 vssd1 vccd1 vccd1 net605 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09743__A1 _05073_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout616 net617 vssd1 vssd1 vccd1 vccd1 net616 sky130_fd_sc_hd__buf_2
XANTENNA__10889__A0 net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_42 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09842_ _05077_ _05783_ _05781_ _05776_ vssd1 vssd1 vccd1 vccd1 _05784_ sky130_fd_sc_hd__o211a_2
Xfanout627 net628 vssd1 vssd1 vccd1 vccd1 net627 sky130_fd_sc_hd__clkbuf_4
Xfanout638 _06458_ vssd1 vssd1 vccd1 vccd1 net638 sky130_fd_sc_hd__clkbuf_4
Xfanout649 net652 vssd1 vssd1 vccd1 vccd1 net649 sky130_fd_sc_hd__buf_4
XANTENNA__07317__A net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09773_ net539 _05713_ vssd1 vssd1 vccd1 vccd1 _05715_ sky130_fd_sc_hd__nand2_1
XFILLER_0_77_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06985_ net1022 _02814_ _02827_ team_03_WB.instance_to_wrap.core.decoder.inst\[14\]
+ vssd1 vssd1 vccd1 vccd1 _02927_ sky130_fd_sc_hd__or4b_4
XANTENNA__11484__D net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout284_A net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08724_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[676\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[644\]
+ net985 vssd1 vssd1 vccd1 vccd1 _04666_ sky130_fd_sc_hd__mux2_1
XANTENNA__07506__B1 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07601__S0 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08655_ net1245 team_03_WB.instance_to_wrap.core.register_file.registers_state\[135\]
+ net990 team_03_WB.instance_to_wrap.core.register_file.registers_state\[167\] net946
+ vssd1 vssd1 vccd1 vccd1 _04597_ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout451_A net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1193_A net1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout549_A _03105_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07606_ net1112 team_03_WB.instance_to_wrap.core.register_file.registers_state\[825\]
+ net902 vssd1 vssd1 vccd1 vccd1 _03548_ sky130_fd_sc_hd__or3_1
X_08586_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[1021\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[989\]
+ net967 vssd1 vssd1 vccd1 vccd1 _04528_ sky130_fd_sc_hd__mux2_1
XFILLER_0_113_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1122 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07809__A1 net1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07537_ net815 _03477_ _03478_ vssd1 vssd1 vccd1 vccd1 _03479_ sky130_fd_sc_hd__and3_1
XFILLER_0_147_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1360_A net1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout337_X net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1079_X net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_338 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07468_ net1184 team_03_WB.instance_to_wrap.core.register_file.registers_state\[597\]
+ net769 team_03_WB.instance_to_wrap.core.register_file.registers_state\[629\] net728
+ vssd1 vssd1 vccd1 vccd1 _03410_ sky130_fd_sc_hd__o221a_1
XANTENNA__11005__C net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09207_ _03866_ _03947_ _04072_ _05147_ net608 vssd1 vssd1 vccd1 vccd1 _05149_ sky130_fd_sc_hd__a41o_1
XANTENNA__10617__S net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout504_X net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07399_ net1146 _03338_ _03340_ net1114 vssd1 vssd1 vccd1 vccd1 _03341_ sky130_fd_sc_hd__o211a_1
XFILLER_0_91_488 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1246_X net1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09138_ net584 _05079_ vssd1 vssd1 vccd1 vccd1 _05080_ sky130_fd_sc_hd__nand2_1
XFILLER_0_32_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12030__A2 net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10041__A1 net16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07442__C1 net1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09069_ net1209 _05010_ _05005_ vssd1 vssd1 vccd1 vccd1 _05011_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout1413_X net1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11100_ _06626_ net2479 net418 vssd1 vssd1 vccd1 vccd1 _02254_ sky130_fd_sc_hd__mux2_1
XANTENNA__07993__B1 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12080_ _06784_ net478 net441 net1960 vssd1 vssd1 vccd1 vccd1 _01467_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout873_X net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold670 team_03_WB.instance_to_wrap.core.register_file.registers_state\[791\] vssd1
+ vssd1 vccd1 vccd1 net2163 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold681 team_03_WB.instance_to_wrap.core.register_file.registers_state\[743\] vssd1
+ vssd1 vccd1 vccd1 net2174 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09734__A1 net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold692 team_03_WB.instance_to_wrap.core.register_file.registers_state\[642\] vssd1
+ vssd1 vccd1 vccd1 net2185 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_498 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11031_ net2552 net422 _06590_ net514 vssd1 vssd1 vccd1 vccd1 _02287_ sky130_fd_sc_hd__a22o_1
XANTENNA__11541__A1 net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12097__A2 net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12982_ net1258 vssd1 vssd1 vccd1 vccd1 _00746_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_86_2146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10859__Y _06458_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14721_ clknet_leaf_44_wb_clk_i _02485_ _01086_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.decoder.inst\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input12_A DAT_I[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11933_ _06629_ net2773 net370 vssd1 vssd1 vccd1 vccd1 _01609_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14652_ clknet_leaf_151_wb_clk_i _02416_ _01017_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1006\]
+ sky130_fd_sc_hd__dfstp_1
X_11864_ net270 net2055 net375 vssd1 vssd1 vccd1 vccd1 _01676_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08058__A net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13603_ net1316 vssd1 vssd1 vccd1 vccd1 _01367_ sky130_fd_sc_hd__inv_2
XFILLER_0_68_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10815_ net686 _05454_ _06401_ vssd1 vssd1 vccd1 vccd1 _06421_ sky130_fd_sc_hd__a21o_1
XFILLER_0_95_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14583_ clknet_leaf_80_wb_clk_i _02347_ _00948_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[937\]
+ sky130_fd_sc_hd__dfstp_1
X_11795_ net2447 _06625_ net329 vssd1 vssd1 vccd1 vccd1 _01743_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_316 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11911__S net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10804__B1 _06401_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13534_ net1317 vssd1 vssd1 vccd1 vccd1 _01298_ sky130_fd_sc_hd__inv_2
X_10746_ net524 _06364_ _06365_ net529 net1611 vssd1 vssd1 vccd1 vccd1 _02443_ sky130_fd_sc_hd__a32o_1
XFILLER_0_40_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08473__A1 net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_147_wb_clk_i clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_147_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_13465_ net1341 vssd1 vssd1 vccd1 vccd1 _01229_ sky130_fd_sc_hd__inv_2
XANTENNA__07681__C1 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10677_ team_03_WB.instance_to_wrap.core.pc.current_pc\[30\] _06318_ vssd1 vssd1
+ vccd1 vccd1 _06319_ sky130_fd_sc_hd__nand2_1
XFILLER_0_82_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08505__B net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12416_ net1402 vssd1 vssd1 vccd1 vccd1 _00180_ sky130_fd_sc_hd__inv_2
XFILLER_0_35_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13396_ net1428 vssd1 vssd1 vccd1 vccd1 _01160_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput208 net208 vssd1 vssd1 vccd1 vccd1 gpio_out[11] sky130_fd_sc_hd__buf_2
XFILLER_0_133_590 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12347_ net1362 vssd1 vssd1 vccd1 vccd1 _00111_ sky130_fd_sc_hd__inv_2
XFILLER_0_105_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput219 net219 vssd1 vssd1 vccd1 vccd1 gpio_out[22] sky130_fd_sc_hd__buf_2
XANTENNA__10583__A2 net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15066_ net1452 vssd1 vssd1 vccd1 vccd1 la_data_out[2] sky130_fd_sc_hd__buf_2
XFILLER_0_26_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12278_ net1280 vssd1 vssd1 vccd1 vccd1 _00042_ sky130_fd_sc_hd__inv_2
X_14017_ clknet_leaf_177_wb_clk_i _01781_ _00382_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[371\]
+ sky130_fd_sc_hd__dfrtp_1
X_11229_ _06536_ net2535 net488 vssd1 vssd1 vccd1 vccd1 _02182_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09904__X _05846_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_147_3386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_147_3397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_58 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12088__A2 net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09352__A _04178_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11296__B1 net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14919_ clknet_leaf_44_wb_clk_i _02674_ _01284_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_O\[6\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__11835__A2 net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08440_ net851 _04368_ _04381_ vssd1 vssd1 vccd1 vccd1 _04382_ sky130_fd_sc_hd__o21ba_4
XTAP_TAPCELL_ROW_19_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_121_2858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_2869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08371_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[566\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[534\]
+ net965 vssd1 vssd1 vccd1 vccd1 _04313_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07303__C net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10785__X _06395_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_173_3925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_173_3936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07322_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[157\] net768
+ net728 _03263_ vssd1 vssd1 vccd1 vccd1 _03264_ sky130_fd_sc_hd__a211o_1
XFILLER_0_45_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_945 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08464__A1 net1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10945__B net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_711 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_171_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07253_ net1176 team_03_WB.instance_to_wrap.core.register_file.registers_state\[200\]
+ net774 team_03_WB.instance_to_wrap.core.register_file.registers_state\[232\] net741
+ vssd1 vssd1 vccd1 vccd1 _03195_ sky130_fd_sc_hd__o221a_1
XFILLER_0_143_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15094__1480 vssd1 vssd1 vccd1 vccd1 _15094__1480/HI net1480 sky130_fd_sc_hd__conb_1
XFILLER_0_147_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11122__A net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_888 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07184_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[563\] net763
+ net726 _03125_ vssd1 vssd1 vccd1 vccd1 _03126_ sky130_fd_sc_hd__o211a_1
XFILLER_0_14_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08216__A1 net1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12012__A2 net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_207 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_3_3_0_wb_clk_i_X clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08134__C _03280_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07424__C1 net1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10574__A2 net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11771__A1 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10680__B net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout499_A net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout402 _06718_ vssd1 vssd1 vccd1 vccd1 net402 sky130_fd_sc_hd__clkbuf_8
Xfanout413 _06635_ vssd1 vssd1 vccd1 vccd1 net413 sky130_fd_sc_hd__buf_4
Xfanout424 net426 vssd1 vssd1 vccd1 vccd1 net424 sky130_fd_sc_hd__buf_2
Xfanout435 net437 vssd1 vssd1 vccd1 vccd1 net435 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07727__B1 net1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11523__B2 net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08924__C1 net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout446 _06816_ vssd1 vssd1 vccd1 vccd1 net446 sky130_fd_sc_hd__buf_4
X_09825_ _04834_ _05568_ _05765_ net595 _05766_ vssd1 vssd1 vccd1 vccd1 _05767_ sky130_fd_sc_hd__o221a_1
Xfanout457 net481 vssd1 vssd1 vccd1 vccd1 net457 sky130_fd_sc_hd__buf_2
XANTENNA_input4_A DAT_I[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout468 net471 vssd1 vssd1 vccd1 vccd1 net468 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout666_A net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout479 net480 vssd1 vssd1 vccd1 vccd1 net479 sky130_fd_sc_hd__clkbuf_2
XANTENNA__12888__A net1376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09756_ _05236_ _05661_ vssd1 vssd1 vccd1 vccd1 _05698_ sky130_fd_sc_hd__xor2_1
X_06968_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[805\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[773\]
+ net789 vssd1 vssd1 vccd1 vccd1 _02910_ sky130_fd_sc_hd__mux2_1
XANTENNA__06950__A1 net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08707_ _04621_ _04648_ vssd1 vssd1 vccd1 vccd1 _04649_ sky130_fd_sc_hd__nor2_1
X_09687_ _04829_ _05513_ _05627_ _05628_ vssd1 vssd1 vccd1 vccd1 _05629_ sky130_fd_sc_hd__a211o_1
XANTENNA__11826__A2 net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06899_ _02837_ net690 vssd1 vssd1 vccd1 vccd1 _02841_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout833_A _06387_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout454_X net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1196_X net1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08638_ net1054 team_03_WB.instance_to_wrap.core.register_file.registers_state\[838\]
+ net1007 team_03_WB.instance_to_wrap.core.register_file.registers_state\[870\] net1215
+ vssd1 vssd1 vccd1 vccd1 _04580_ sky130_fd_sc_hd__a221o_1
XFILLER_0_68_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10201__A _02990_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_2032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_2043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11039__B1 net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08569_ net858 _04509_ _04510_ vssd1 vssd1 vccd1 vccd1 _04511_ sky130_fd_sc_hd__or3_1
XANTENNA_fanout621_X net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1086 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1363_X net1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout719_X net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10600_ net2114 net1808 net841 vssd1 vssd1 vccd1 vccd1 _02528_ sky130_fd_sc_hd__mux2_1
X_11580_ net302 net2525 net450 vssd1 vssd1 vccd1 vccd1 _01949_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_967 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10855__B net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07510__A net1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10531_ net166 net1034 net1026 net1725 vssd1 vssd1 vccd1 vccd1 _02579_ sky130_fd_sc_hd__a22o_1
XANTENNA__08550__S1 net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10347__S net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11032__A net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13250_ net1289 vssd1 vssd1 vccd1 vccd1 _01014_ sky130_fd_sc_hd__inv_2
X_10462_ team_03_WB.instance_to_wrap.core.pc.current_pc\[3\] team_03_WB.instance_to_wrap.core.pc.current_pc\[2\]
+ vssd1 vssd1 vccd1 vccd1 _06276_ sky130_fd_sc_hd__or2_1
XFILLER_0_10_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout990_X net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12201_ net1517 vssd1 vssd1 vccd1 vccd1 _02352_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__11211__A0 _06468_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13181_ net1383 vssd1 vssd1 vccd1 vccd1 _00945_ sky130_fd_sc_hd__inv_2
X_10393_ team_03_WB.instance_to_wrap.core.pc.current_pc\[16\] _06142_ vssd1 vssd1
+ vccd1 vccd1 _06220_ sky130_fd_sc_hd__nor2_1
XANTENNA__10871__A net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10565__A2 net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07966__B1 net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12132_ net1521 vssd1 vssd1 vccd1 vccd1 _02421_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_36_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10590__B _05914_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12063_ _06628_ net2490 net358 vssd1 vssd1 vccd1 vccd1 _01483_ sky130_fd_sc_hd__mux2_1
X_11014_ net493 net647 _06580_ net420 net2072 vssd1 vssd1 vccd1 vccd1 _02294_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_53_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout980 net981 vssd1 vssd1 vccd1 vccd1 net980 sky130_fd_sc_hd__clkbuf_4
Xfanout991 net993 vssd1 vssd1 vccd1 vccd1 net991 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_5_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_37 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11278__B1 net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input15_X net15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_142_3283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11817__A2 net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12965_ net1349 vssd1 vssd1 vccd1 vccd1 _00729_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_142_3294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_103_2500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_251 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14704_ clknet_leaf_32_wb_clk_i _02468_ _01069_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.control_logic.instruction\[1\]
+ sky130_fd_sc_hd__dfrtp_4
X_11916_ _06617_ net2557 net368 vssd1 vssd1 vccd1 vccd1 _01626_ sky130_fd_sc_hd__mux2_1
XANTENNA__10111__A _04807_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08694__A1 net1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12896_ net1402 vssd1 vssd1 vccd1 vccd1 _00660_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_16_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14635_ clknet_leaf_50_wb_clk_i _02399_ _01000_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[989\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_142_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11847_ net302 net2043 net377 vssd1 vssd1 vccd1 vccd1 _01693_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_772 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14566_ clknet_leaf_72_wb_clk_i _02330_ _00931_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[920\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08446__A1 net1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11778_ net2370 _06611_ net328 vssd1 vssd1 vccd1 vccd1 _01760_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_166_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13517_ net1307 vssd1 vssd1 vccd1 vccd1 _01281_ sky130_fd_sc_hd__inv_2
X_10729_ net1985 net528 net523 _06356_ vssd1 vssd1 vccd1 vccd1 _02451_ sky130_fd_sc_hd__a22o_1
XFILLER_0_153_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14497_ clknet_leaf_179_wb_clk_i _02261_ _00862_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[851\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_83_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13448_ net1407 vssd1 vssd1 vccd1 vccd1 _01212_ sky130_fd_sc_hd__inv_2
Xclkload12 clknet_leaf_187_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload12/Y sky130_fd_sc_hd__clkinv_2
XFILLER_0_67_1148 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkload23 clknet_leaf_12_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload23/Y sky130_fd_sc_hd__inv_8
XANTENNA__11299__D _06463_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload34 clknet_leaf_180_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload34/Y sky130_fd_sc_hd__bufinv_16
XANTENNA__11202__A0 net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07406__C1 net1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload45 clknet_leaf_25_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload45/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_141_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload56 clknet_leaf_34_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload56/X sky130_fd_sc_hd__clkbuf_4
X_13379_ net1430 vssd1 vssd1 vccd1 vccd1 _01143_ sky130_fd_sc_hd__inv_2
Xclkload67 clknet_leaf_47_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload67/Y sky130_fd_sc_hd__clkinvlp_4
XTAP_TAPCELL_ROW_77_1956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload78 clknet_leaf_58_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload78/Y sky130_fd_sc_hd__clkinv_4
XTAP_TAPCELL_ROW_77_1967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_149_3426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15118_ net915 vssd1 vssd1 vccd1 vccd1 net250 sky130_fd_sc_hd__clkbuf_1
Xclkload89 clknet_leaf_71_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload89/Y sky130_fd_sc_hd__clkinv_4
XANTENNA__09347__A _04148_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_149_3437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15049_ net1490 vssd1 vssd1 vccd1 vccd1 gpio_oeb[1] sky130_fd_sc_hd__buf_2
X_07940_ _03880_ _03881_ net822 vssd1 vssd1 vccd1 vccd1 _03882_ sky130_fd_sc_hd__o21a_1
XFILLER_0_167_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_166_3773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_166_3784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_44_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_44_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08906__C1 net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07871_ net1200 team_03_WB.instance_to_wrap.core.register_file.registers_state\[91\]
+ net781 team_03_WB.instance_to_wrap.core.register_file.registers_state\[123\] net737
+ vssd1 vssd1 vccd1 vccd1 _03813_ sky130_fd_sc_hd__o221a_1
XANTENNA__07185__A1 net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09610_ _05551_ vssd1 vssd1 vccd1 vccd1 _05552_ sky130_fd_sc_hd__inv_2
X_06822_ net1143 vssd1 vssd1 vccd1 vccd1 _02765_ sky130_fd_sc_hd__inv_2
XANTENNA__12501__A net1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_2909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06932__B2 net1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09541_ _05398_ _05401_ net556 vssd1 vssd1 vccd1 vccd1 _05483_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09472_ net542 _04296_ _05087_ vssd1 vssd1 vccd1 vccd1 _05414_ sky130_fd_sc_hd__a21oi_1
X_08423_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[442\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[410\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[314\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[282\]
+ net954 net1072 vssd1 vssd1 vccd1 vccd1 _04365_ sky130_fd_sc_hd__mux4_1
XFILLER_0_65_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08354_ net438 net426 _04295_ vssd1 vssd1 vccd1 vccd1 _04296_ sky130_fd_sc_hd__or3_2
XFILLER_0_46_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10675__B _06316_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07305_ net1185 team_03_WB.instance_to_wrap.core.register_file.registers_state\[733\]
+ net768 team_03_WB.instance_to_wrap.core.register_file.registers_state\[765\] net743
+ vssd1 vssd1 vccd1 vccd1 _03247_ sky130_fd_sc_hd__o221a_1
XFILLER_0_46_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload6 clknet_leaf_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload6/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_62_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08285_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[631\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[599\]
+ net963 vssd1 vssd1 vccd1 vccd1 _04227_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout414_A _06635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1156_A net1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09956__S net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07236_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[904\] net796
+ _03171_ net1154 vssd1 vssd1 vccd1 vccd1 _03178_ sky130_fd_sc_hd__o211a_1
XFILLER_0_6_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_143_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10691__A net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07167_ _03108_ vssd1 vssd1 vccd1 vccd1 _03109_ sky130_fd_sc_hd__inv_2
XFILLER_0_70_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07099__S1 net1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_711 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07098_ net1165 _03038_ vssd1 vssd1 vccd1 vccd1 _03040_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout783_A net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07048__Y _02990_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1208 net1209 vssd1 vssd1 vccd1 vccd1 net1208 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout1111_X net1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1219 net1220 vssd1 vssd1 vccd1 vccd1 net1219 sky130_fd_sc_hd__buf_4
XANTENNA_fanout1209_X net1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input7_X net7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout950_A net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07176__A1 net1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout265 _06528_ vssd1 vssd1 vccd1 vccd1 net265 sky130_fd_sc_hd__buf_2
Xfanout276 _06434_ vssd1 vssd1 vccd1 vccd1 net276 sky130_fd_sc_hd__buf_2
XANTENNA__11726__S net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout669_X net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09808_ _02923_ _04565_ net540 vssd1 vssd1 vccd1 vccd1 _05750_ sky130_fd_sc_hd__o21ai_1
Xfanout287 net290 vssd1 vssd1 vccd1 vccd1 net287 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10630__S net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10180__B1 _03242_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout298 _06495_ vssd1 vssd1 vccd1 vccd1 net298 sky130_fd_sc_hd__buf_2
Xclkbuf_4_15__f_wb_clk_i clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_15__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_158_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09739_ _03790_ _04953_ _05680_ net667 vssd1 vssd1 vccd1 vccd1 _05681_ sky130_fd_sc_hd__a22o_1
XFILLER_0_119_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout836_X net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08125__B1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11027__A net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12750_ net1270 vssd1 vssd1 vccd1 vccd1 _00514_ sky130_fd_sc_hd__inv_2
XANTENNA__07479__A2 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_901 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11701_ _06743_ net386 net341 net1950 vssd1 vssd1 vccd1 vccd1 _01833_ sky130_fd_sc_hd__a22o_1
XFILLER_0_55_1096 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12681_ net1260 vssd1 vssd1 vccd1 vccd1 _00445_ sky130_fd_sc_hd__inv_2
XANTENNA__11680__B1 net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13242__A net1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14420_ clknet_leaf_123_wb_clk_i _02184_ _00785_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[774\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_77_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_166_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_154_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11632_ _06706_ net379 net346 net2515 vssd1 vssd1 vccd1 vccd1 _01900_ sky130_fd_sc_hd__a22o_1
XANTENNA__08428__A1 net1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14351_ clknet_leaf_136_wb_clk_i _02115_ _00716_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[705\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11432__B1 net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10077__S net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11563_ net636 net706 _06527_ net697 vssd1 vssd1 vccd1 vccd1 _06796_ sky130_fd_sc_hd__and4_1
XANTENNA__07100__B2 net1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13302_ net1322 vssd1 vssd1 vccd1 vccd1 _01066_ sky130_fd_sc_hd__inv_2
XFILLER_0_107_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10514_ net153 net1031 net1023 net1997 vssd1 vssd1 vccd1 vccd1 _02596_ sky130_fd_sc_hd__a22o_1
X_14282_ clknet_leaf_7_wb_clk_i _02046_ _00647_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[636\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_98_2381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11494_ _06615_ net2749 net388 vssd1 vssd1 vccd1 vccd1 _02012_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_98_2392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13233_ net1269 vssd1 vssd1 vccd1 vccd1 _00997_ sky130_fd_sc_hd__inv_2
X_10445_ team_03_WB.instance_to_wrap.core.pc.current_pc\[7\] net682 _06260_ _06262_
+ vssd1 vssd1 vccd1 vccd1 _02641_ sky130_fd_sc_hd__o22a_1
XFILLER_0_27_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_823 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10538__A2 net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_55_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13164_ net1314 vssd1 vssd1 vccd1 vccd1 _00928_ sky130_fd_sc_hd__inv_2
XFILLER_0_32_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_55_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08061__C1 net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10376_ team_03_WB.instance_to_wrap.core.pc.current_pc\[18\] _06144_ team_03_WB.instance_to_wrap.core.pc.current_pc\[19\]
+ vssd1 vssd1 vccd1 vccd1 _06206_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_27_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08071__A net1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12115_ _06287_ _06289_ vssd1 vssd1 vccd1 vccd1 _00007_ sky130_fd_sc_hd__nand2_1
X_13095_ net1400 vssd1 vssd1 vccd1 vccd1 _00859_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_72_1853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_16 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12046_ _06615_ net2716 net356 vssd1 vssd1 vccd1 vccd1 _01500_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_144_3323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_3334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10171__B1 _03758_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_161_3681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13997_ clknet_leaf_187_wb_clk_i _01761_ _00362_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[351\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12040__B net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_322 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12948_ net1313 vssd1 vssd1 vccd1 vccd1 _00712_ sky130_fd_sc_hd__inv_2
XFILLER_0_88_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08667__A1 net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08945__S net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09630__A net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_162_wb_clk_i clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_162_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_75_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12879_ net1363 vssd1 vssd1 vccd1 vccd1 _00643_ sky130_fd_sc_hd__inv_2
X_14618_ clknet_leaf_148_wb_clk_i _02382_ _00983_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[972\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_139_980 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11423__A0 net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14549_ clknet_leaf_107_wb_clk_i _02313_ _00914_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[903\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_28_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_674 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08070_ net1088 net893 team_03_WB.instance_to_wrap.core.register_file.registers_state\[534\]
+ vssd1 vssd1 vccd1 vccd1 _04012_ sky130_fd_sc_hd__o21a_1
XANTENNA__08533__X _04475_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload101 clknet_leaf_148_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload101/X sky130_fd_sc_hd__clkbuf_4
Xclkload112 clknet_leaf_119_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload112/Y sky130_fd_sc_hd__inv_6
XTAP_TAPCELL_ROW_116_2757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload123 clknet_leaf_136_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload123/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_114_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07021_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[515\] net801
+ net731 _02962_ vssd1 vssd1 vccd1 vccd1 _02963_ sky130_fd_sc_hd__o211a_1
Xclkload134 clknet_leaf_125_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload134/Y sky130_fd_sc_hd__clkinv_8
Xclkload145 clknet_leaf_79_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload145/Y sky130_fd_sc_hd__clkinvlp_4
XTAP_TAPCELL_ROW_116_2768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08278__S0 net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload156 clknet_leaf_110_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload156/X sky130_fd_sc_hd__clkbuf_8
XANTENNA__10529__A2 net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload167 clknet_leaf_127_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload167/Y sky130_fd_sc_hd__inv_6
XANTENNA__11726__A1 _06483_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_168_3824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload178 clknet_leaf_94_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload178/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_113_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_355 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08972_ net945 _04913_ _04912_ net1067 vssd1 vssd1 vccd1 vccd1 _04914_ sky130_fd_sc_hd__o211a_1
X_07923_ net611 _03844_ _03863_ vssd1 vssd1 vccd1 vccd1 _03865_ sky130_fd_sc_hd__or3_1
Xhold18 team_03_WB.instance_to_wrap.core.register_file.registers_state\[936\] vssd1
+ vssd1 vccd1 vccd1 net1511 sky130_fd_sc_hd__dlygate4sd3_1
Xhold29 team_03_WB.instance_to_wrap.core.register_file.registers_state\[975\] vssd1
+ vssd1 vccd1 vccd1 net1522 sky130_fd_sc_hd__dlygate4sd3_1
X_07854_ net1202 team_03_WB.instance_to_wrap.core.register_file.registers_state\[987\]
+ net784 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1019\] net1167
+ vssd1 vssd1 vccd1 vccd1 _03796_ sky130_fd_sc_hd__o221a_1
XFILLER_0_39_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09016__S net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07785_ _03725_ _03726_ vssd1 vssd1 vccd1 vccd1 _03727_ sky130_fd_sc_hd__or2_2
XANTENNA_fanout364_A _06815_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09524_ _05465_ vssd1 vssd1 vccd1 vccd1 _05466_ sky130_fd_sc_hd__inv_2
XFILLER_0_149_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08855__S net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09455_ _05393_ _05396_ net567 vssd1 vssd1 vccd1 vccd1 _05397_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout531_A net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_232 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06883__B team_03_WB.instance_to_wrap.core.decoder.inst\[27\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout629_A net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1273_A net1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08406_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[825\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[793\]
+ net993 vssd1 vssd1 vccd1 vccd1 _04348_ sky130_fd_sc_hd__mux2_1
XANTENNA__13062__A net1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09386_ _04267_ _05326_ vssd1 vssd1 vccd1 vccd1 _05328_ sky130_fd_sc_hd__and2_1
XFILLER_0_4_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_49_Left_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08337_ _04275_ _04276_ _04278_ _04277_ net920 net861 vssd1 vssd1 vccd1 vccd1 _04279_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_4_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1061_X net1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11965__A1 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout417_X net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_419 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1159_X net1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08268_ net548 _04179_ _04209_ vssd1 vssd1 vccd1 vccd1 _04210_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_6_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11013__C net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout998_A net999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07219_ net1170 team_03_WB.instance_to_wrap.core.register_file.registers_state\[978\]
+ net757 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1010\] net1149
+ vssd1 vssd1 vccd1 vccd1 _03161_ sky130_fd_sc_hd__o221a_1
XFILLER_0_46_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10625__S net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12406__A net1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08199_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[819\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[787\]
+ net957 vssd1 vssd1 vccd1 vccd1 _04141_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1326_X net1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11717__A1 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_368 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10230_ net589 net674 vssd1 vssd1 vccd1 vccd1 _06072_ sky130_fd_sc_hd__or2_1
XANTENNA_clkbuf_leaf_35_wb_clk_i_A clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_132_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout786_X net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10161_ _06000_ _06001_ _03679_ vssd1 vssd1 vccd1 vccd1 _06003_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_7_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07492__S1 net1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10940__A2 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1005 net1008 vssd1 vssd1 vccd1 vccd1 net1005 sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_EDGE_ROW_58_Left_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1027 net1028 vssd1 vssd1 vccd1 vccd1 net1027 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_50_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10092_ _05563_ _05647_ _05933_ _05935_ vssd1 vssd1 vccd1 vccd1 _05936_ sky130_fd_sc_hd__nand4_1
Xfanout1038 _05905_ vssd1 vssd1 vccd1 vccd1 net1038 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_50_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07149__A1 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1049 net1060 vssd1 vssd1 vccd1 vccd1 net1049 sky130_fd_sc_hd__buf_4
XANTENNA__08346__B1 net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13920_ clknet_leaf_2_wb_clk_i _01684_ _00285_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[274\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08897__A1 net1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13851_ clknet_leaf_145_wb_clk_i _01615_ _00216_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[205\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08992__S1 net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1147 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15073__1459 vssd1 vssd1 vccd1 vccd1 _15073__1459/HI net1459 sky130_fd_sc_hd__conb_1
X_12802_ net1296 vssd1 vssd1 vccd1 vccd1 _00566_ sky130_fd_sc_hd__inv_2
X_13782_ clknet_leaf_154_wb_clk_i _01546_ _00147_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[136\]
+ sky130_fd_sc_hd__dfrtp_1
X_10994_ net1044 net836 _06418_ net670 vssd1 vssd1 vccd1 vccd1 _06569_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_48_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12733_ net1389 vssd1 vssd1 vccd1 vccd1 _00497_ sky130_fd_sc_hd__inv_2
XANTENNA__07857__C1 net1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_67_Left_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_1072 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12664_ net1375 vssd1 vssd1 vccd1 vccd1 _00428_ sky130_fd_sc_hd__inv_2
XFILLER_0_32_49 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08066__A net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11405__A0 _06430_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14403_ clknet_leaf_34_wb_clk_i _02167_ _00768_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[757\]
+ sky130_fd_sc_hd__dfrtp_1
X_11615_ _06689_ net385 net349 net2220 vssd1 vssd1 vccd1 vccd1 _01917_ sky130_fd_sc_hd__a22o_1
XFILLER_0_143_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09074__A1 net1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_74_wb_clk_i_A clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_26_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12595_ net1255 vssd1 vssd1 vccd1 vccd1 _00359_ sky130_fd_sc_hd__inv_2
XANTENNA__09074__B2 net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_3182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_3193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11956__A1 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07085__B1 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14334_ clknet_leaf_118_wb_clk_i _02098_ _00699_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[688\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11546_ net513 net641 _06656_ net485 net1926 vssd1 vssd1 vccd1 vccd1 _01970_ sky130_fd_sc_hd__a32o_1
XFILLER_0_53_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10085__A_N _05757_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14265_ clknet_leaf_155_wb_clk_i _02029_ _00630_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[619\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_64_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11477_ net636 net705 _06527_ net829 vssd1 vssd1 vccd1 vccd1 _06774_ sky130_fd_sc_hd__and4_1
XANTENNA__11220__A _06456_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_1904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13216_ net1403 vssd1 vssd1 vccd1 vccd1 _00980_ sky130_fd_sc_hd__inv_2
X_10428_ net285 _06139_ _06246_ net682 vssd1 vssd1 vccd1 vccd1 _06249_ sky130_fd_sc_hd__o31a_1
XFILLER_0_111_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08034__C1 net1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_164_Right_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14196_ clknet_leaf_124_wb_clk_i _01960_ _00561_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[550\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_76_Left_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_111_2654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13147_ net1362 vssd1 vssd1 vccd1 vccd1 _00911_ sky130_fd_sc_hd__inv_2
X_10359_ _06191_ _06192_ team_03_WB.instance_to_wrap.core.pc.current_pc\[23\] net679
+ vssd1 vssd1 vccd1 vccd1 _02657_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_111_2665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_35 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09184__X _05126_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07844__S net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_163_3721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13078_ net1260 vssd1 vssd1 vccd1 vccd1 _00842_ sky130_fd_sc_hd__inv_2
X_12029_ net620 _06595_ net452 net359 net2172 vssd1 vssd1 vccd1 vccd1 _01516_ sky130_fd_sc_hd__a32o_1
XFILLER_0_164_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_164_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11892__B1 net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12986__A net1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07560__A1 net1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07570_ net1106 team_03_WB.instance_to_wrap.core.register_file.registers_state\[696\]
+ net903 vssd1 vssd1 vccd1 vccd1 _03512_ sky130_fd_sc_hd__or3_1
XANTENNA__10777__Y _06387_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_85_Left_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07312__A1 net1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10998__A2 net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09240_ _04323_ _05179_ vssd1 vssd1 vccd1 vccd1 _05182_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_173_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_146_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_173_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_118_2808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09171_ _05111_ _05112_ vssd1 vssd1 vccd1 vccd1 _05113_ sky130_fd_sc_hd__nor2_1
XFILLER_0_111_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09065__A1 net1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11947__A1 net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08122_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[794\] net793
+ net1041 _04063_ vssd1 vssd1 vccd1 vccd1 _04064_ sky130_fd_sc_hd__o211a_1
XFILLER_0_83_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_wire587_X net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_994 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08812__A1 net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08273__C1 net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_142_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08053_ _03992_ _03994_ net812 vssd1 vssd1 vccd1 vccd1 _03995_ sky130_fd_sc_hd__a21o_1
XFILLER_0_25_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_141_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07004_ team_03_WB.instance_to_wrap.core.decoder.inst\[13\] _02929_ _02827_ _02836_
+ vssd1 vssd1 vccd1 vccd1 _02946_ sky130_fd_sc_hd__or4b_1
XFILLER_0_24_491 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_141_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_131_Right_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_686 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07918__A3 net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1021_A net1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10922__A2 _05706_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1119_A net1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_119_wb_clk_i_A clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_08955_ net1245 team_03_WB.instance_to_wrap.core.register_file.registers_state\[169\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[137\] net991 net929
+ vssd1 vssd1 vccd1 vccd1 _04897_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout579_A _02993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07906_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[527\] net771
+ net745 _03847_ vssd1 vssd1 vccd1 vccd1 _03848_ sky130_fd_sc_hd__a211o_1
X_08886_ _04827_ vssd1 vssd1 vccd1 vccd1 _04828_ sky130_fd_sc_hd__inv_2
XFILLER_0_98_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07837_ _03777_ _03778_ vssd1 vssd1 vccd1 vccd1 _03779_ sky130_fd_sc_hd__and2_1
XANTENNA__11883__B1 net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12896__A net1402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout746_A net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout367_X net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07768_ net1194 team_03_WB.instance_to_wrap.core.register_file.registers_state\[844\]
+ vssd1 vssd1 vccd1 vccd1 _03710_ sky130_fd_sc_hd__or2_1
XFILLER_0_168_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09507_ _05353_ _05374_ net563 vssd1 vssd1 vccd1 vccd1 _05449_ sky130_fd_sc_hd__mux2_1
XANTENNA__09270__A net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_163 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11635__B1 net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07699_ _03638_ _03640_ net610 vssd1 vssd1 vccd1 vccd1 _03641_ sky130_fd_sc_hd__mux2_2
XANTENNA_fanout534_X net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09438_ _04593_ _04621_ vssd1 vssd1 vccd1 vccd1 _05380_ sky130_fd_sc_hd__nor2_1
XFILLER_0_137_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11024__B net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09369_ _05310_ vssd1 vssd1 vccd1 vccd1 _05311_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout701_X net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11400_ net280 net2622 net396 vssd1 vssd1 vccd1 vccd1 _02080_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12380_ net1411 vssd1 vssd1 vccd1 vccd1 _00144_ sky130_fd_sc_hd__inv_2
XANTENNA__08803__A1 net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11331_ _06633_ net2779 net406 vssd1 vssd1 vccd1 vccd1 _02114_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_158_wb_clk_i_A clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11040__A net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14050_ clknet_leaf_175_wb_clk_i _01814_ _00415_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[404\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_132_3090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11262_ net490 net618 _06698_ net408 net2134 vssd1 vssd1 vccd1 vccd1 _02164_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_91_2237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_2248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08567__B1 net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13001_ net1254 vssd1 vssd1 vccd1 vccd1 _00765_ sky130_fd_sc_hd__inv_2
XANTENNA__11166__A2 net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10213_ _06037_ _06053_ _06035_ vssd1 vssd1 vccd1 vccd1 _06055_ sky130_fd_sc_hd__a21oi_1
X_11193_ net505 net654 _06677_ net414 net1915 vssd1 vssd1 vccd1 vccd1 _02212_ sky130_fd_sc_hd__a32o_1
XANTENNA__08662__S0 net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07517__X _03459_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input42_A gpio_in[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10144_ _03109_ _05985_ vssd1 vssd1 vccd1 vccd1 _05986_ sky130_fd_sc_hd__and2_1
XANTENNA__08319__B1 net999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10075_ _05346_ _05347_ _05386_ _05341_ vssd1 vssd1 vccd1 vccd1 _05919_ sky130_fd_sc_hd__a211o_1
X_14952_ clknet_leaf_103_wb_clk_i _02704_ _01317_ vssd1 vssd1 vccd1 vccd1 net235 sky130_fd_sc_hd__dfrtp_1
XANTENNA__09531__A2 _04354_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13903_ clknet_leaf_144_wb_clk_i _01667_ _00268_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[257\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11874__A0 net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_2199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14883_ clknet_leaf_81_wb_clk_i _02646_ _01248_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.pc.current_pc\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10103__B net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11914__S net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13834_ clknet_leaf_3_wb_clk_i _01598_ _00199_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[188\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_67_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_67_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10429__B2 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11626__B1 net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13765_ clknet_leaf_11_wb_clk_i _01529_ _00130_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[119\]
+ sky130_fd_sc_hd__dfrtp_1
X_10977_ net692 _06552_ _06553_ _06555_ vssd1 vssd1 vccd1 vccd1 _06556_ sky130_fd_sc_hd__a31o_1
XANTENNA__09295__A1 net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_139_3222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_139_3233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12716_ net1311 vssd1 vssd1 vccd1 vccd1 _00480_ sky130_fd_sc_hd__inv_2
X_13696_ clknet_leaf_190_wb_clk_i _01460_ _00061_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[50\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12647_ net1369 vssd1 vssd1 vccd1 vccd1 _00411_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_156_3580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07839__S net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12578_ net1350 vssd1 vssd1 vccd1 vccd1 _00342_ sky130_fd_sc_hd__inv_2
XFILLER_0_41_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_430 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_152_3488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11529_ net658 _06641_ vssd1 vssd1 vccd1 vccd1 _06783_ sky130_fd_sc_hd__nor2_1
X_14317_ clknet_leaf_183_wb_clk_i _02081_ _00682_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[671\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_152_3499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_2705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold307 team_03_WB.instance_to_wrap.core.register_file.registers_state\[296\] vssd1
+ vssd1 vccd1 vccd1 net1800 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_394 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_236 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold318 net189 vssd1 vssd1 vccd1 vccd1 net1811 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_151_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold329 _02583_ vssd1 vssd1 vccd1 vccd1 net1822 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08007__C1 net1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14248_ clknet_leaf_10_wb_clk_i _02012_ _00613_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[602\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_269 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08558__B1 net1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14179_ clknet_leaf_32_wb_clk_i _01943_ _00544_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[533\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout809 net810 vssd1 vssd1 vccd1 vccd1 net809 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_0_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11096__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08740_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[3\] net1004
+ net926 _04681_ vssd1 vssd1 vccd1 vccd1 _04682_ sky130_fd_sc_hd__o211a_1
Xhold1007 team_03_WB.instance_to_wrap.core.register_file.registers_state\[516\] vssd1
+ vssd1 vccd1 vccd1 net2500 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_84_44 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1018 team_03_WB.instance_to_wrap.core.register_file.registers_state\[485\] vssd1
+ vssd1 vccd1 vccd1 net2511 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10117__B1 _03065_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1029 team_03_WB.instance_to_wrap.core.register_file.registers_state\[162\] vssd1
+ vssd1 vccd1 vccd1 net2522 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11865__A0 net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1380 net1381 vssd1 vssd1 vccd1 vccd1 net1380 sky130_fd_sc_hd__buf_4
Xfanout1391 net1392 vssd1 vssd1 vccd1 vccd1 net1391 sky130_fd_sc_hd__buf_2
X_08671_ net1057 team_03_WB.instance_to_wrap.core.register_file.registers_state\[679\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[647\] net1011 net946
+ vssd1 vssd1 vccd1 vccd1 _04613_ sky130_fd_sc_hd__o221a_1
XFILLER_0_139_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13605__A net1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07622_ team_03_WB.instance_to_wrap.core.decoder.inst\[25\] net1020 vssd1 vssd1 vccd1
+ vccd1 _03564_ sky130_fd_sc_hd__nand2_1
XFILLER_0_89_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07162__X _03104_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11880__A3 net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11617__B1 net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07553_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[152\] net783
+ net734 _03494_ vssd1 vssd1 vccd1 vccd1 _03495_ sky130_fd_sc_hd__a211o_1
XFILLER_0_88_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07484_ net1162 net1019 net684 vssd1 vssd1 vccd1 vccd1 _03426_ sky130_fd_sc_hd__a21o_1
XFILLER_0_119_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09223_ _04503_ _05163_ vssd1 vssd1 vccd1 vccd1 _05165_ sky130_fd_sc_hd__and2_1
XFILLER_0_29_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout327_A _06810_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13340__A net1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09154_ net432 net424 _04354_ net542 vssd1 vssd1 vccd1 vccd1 _05096_ sky130_fd_sc_hd__o31a_1
XANTENNA__09589__A2 _02804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08246__C1 net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08105_ _04045_ _04046_ net820 vssd1 vssd1 vccd1 vccd1 _04047_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_71_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11396__A2 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09085_ _05021_ _05026_ net873 vssd1 vssd1 vccd1 vccd1 _05027_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1236_A net1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15072__1458 vssd1 vssd1 vccd1 vccd1 _15072__1458/HI net1458 sky130_fd_sc_hd__conb_1
XFILLER_0_47_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09964__S net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08036_ net1086 team_03_WB.instance_to_wrap.core.register_file.registers_state\[433\]
+ net890 net1014 vssd1 vssd1 vccd1 vccd1 _03978_ sky130_fd_sc_hd__o31a_1
XFILLER_0_114_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput90 wbs_adr_i[30] vssd1 vssd1 vccd1 vccd1 net90 sky130_fd_sc_hd__buf_1
XANTENNA__10970__Y _06550_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold830 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[0\] vssd1 vssd1 vccd1
+ vccd1 net2323 sky130_fd_sc_hd__dlygate4sd3_1
Xhold841 team_03_WB.instance_to_wrap.core.register_file.registers_state\[872\] vssd1
+ vssd1 vccd1 vccd1 net2334 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout696_A _06561_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold852 team_03_WB.instance_to_wrap.core.register_file.registers_state\[497\] vssd1
+ vssd1 vccd1 vccd1 net2345 sky130_fd_sc_hd__dlygate4sd3_1
Xhold863 team_03_WB.instance_to_wrap.core.register_file.registers_state\[472\] vssd1
+ vssd1 vccd1 vccd1 net2356 sky130_fd_sc_hd__dlygate4sd3_1
Xhold874 team_03_WB.instance_to_wrap.core.register_file.registers_state\[788\] vssd1
+ vssd1 vccd1 vccd1 net2367 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1024_X net1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06889__A team_03_WB.instance_to_wrap.core.decoder.inst\[12\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1403_A net1408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold885 team_03_WB.instance_to_wrap.core.register_file.registers_state\[164\] vssd1
+ vssd1 vccd1 vccd1 net2378 sky130_fd_sc_hd__dlygate4sd3_1
Xhold896 team_03_WB.instance_to_wrap.core.register_file.registers_state\[889\] vssd1
+ vssd1 vccd1 vccd1 net2389 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09265__A _05041_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09987_ _05872_ net1695 net290 vssd1 vssd1 vccd1 vccd1 _02727_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout484_X net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout863_A net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07772__A1 net1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08938_ net1217 _04879_ _04878_ net1211 vssd1 vssd1 vccd1 vccd1 _04880_ sky130_fd_sc_hd__o211a_1
XFILLER_0_157_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10659__A1 team_03_WB.instance_to_wrap.CPU_DAT_O\[2\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_99_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11019__B net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08869_ _04770_ _04809_ _04810_ vssd1 vssd1 vccd1 vccd1 _04811_ sky130_fd_sc_hd__or3_1
XANTENNA_fanout651_X net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout749_X net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1393_X net1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10900_ net691 _05659_ net586 vssd1 vssd1 vccd1 vccd1 _06492_ sky130_fd_sc_hd__o21a_1
X_11880_ net640 _06689_ net475 net373 net2142 vssd1 vssd1 vccd1 vccd1 _01661_ sky130_fd_sc_hd__a32o_1
XFILLER_0_169_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_28_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10831_ _06431_ _06433_ _06401_ vssd1 vssd1 vccd1 vccd1 _06434_ sky130_fd_sc_hd__a21oi_4
XANTENNA_fanout916_X net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_179 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11035__A net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13550_ net1420 vssd1 vssd1 vccd1 vccd1 _01314_ sky130_fd_sc_hd__inv_2
XANTENNA__07288__B1 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10762_ _02775_ _06294_ vssd1 vssd1 vccd1 vccd1 _06375_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_11_Right_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_165_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12501_ net1291 vssd1 vssd1 vccd1 vccd1 _00265_ sky130_fd_sc_hd__inv_2
XFILLER_0_48_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13481_ net1407 vssd1 vssd1 vccd1 vccd1 _01245_ sky130_fd_sc_hd__inv_2
XANTENNA__09029__A1 net1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10693_ net1699 net527 net522 _06332_ vssd1 vssd1 vccd1 vccd1 _02463_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_62_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_134_3130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12432_ net1412 vssd1 vssd1 vccd1 vccd1 _00196_ sky130_fd_sc_hd__inv_2
XFILLER_0_30_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12033__B1 net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08344__A net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_350 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12363_ net1288 vssd1 vssd1 vccd1 vccd1 _00127_ sky130_fd_sc_hd__inv_2
XFILLER_0_164_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10595__B1 net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_3038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14102_ clknet_leaf_176_wb_clk_i _01866_ _00467_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[456\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_130_3049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11314_ _06479_ net2594 net404 vssd1 vssd1 vccd1 vccd1 _02131_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_556 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15082_ net1468 vssd1 vssd1 vccd1 vccd1 la_data_out[18] sky130_fd_sc_hd__buf_2
XANTENNA__07460__B1 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12294_ net1337 vssd1 vssd1 vccd1 vccd1 _00058_ sky130_fd_sc_hd__inv_2
XANTENNA__11139__A2 net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14033_ clknet_leaf_143_wb_clk_i _01797_ _00398_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[387\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11909__S net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11245_ net1247 net836 net278 net670 vssd1 vssd1 vccd1 vccd1 _06690_ sky130_fd_sc_hd__and4_1
XPHY_EDGE_ROW_20_Right_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07394__S net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09752__A2 net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11176_ net641 _06667_ vssd1 vssd1 vccd1 vccd1 _06668_ sky130_fd_sc_hd__nor2_1
XFILLER_0_98_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10127_ _05968_ vssd1 vssd1 vccd1 vccd1 _05969_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09504__A2 _04444_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11847__A0 net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14935_ clknet_leaf_53_wb_clk_i _02690_ _01300_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_O\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_10058_ net29 net1039 net911 team_03_WB.instance_to_wrap.CPU_DAT_O\[5\] vssd1 vssd1
+ vccd1 vccd1 _02673_ sky130_fd_sc_hd__a22o_1
XANTENNA__07515__A1 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11644__S net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08712__B1 net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14866_ clknet_leaf_60_wb_clk_i _02630_ _01231_ vssd1 vssd1 vccd1 vccd1 net122 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_106_2553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10768__B net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07423__A net1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13817_ clknet_leaf_162_wb_clk_i _01581_ _00182_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[171\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_158_3620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14797_ clknet_leaf_87_wb_clk_i _02561_ _01162_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_I\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_69_wb_clk_i clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_69_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__07279__B1 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_831 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_678 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13748_ clknet_leaf_131_wb_clk_i _01512_ _00113_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[102\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_174_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_154_3528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_154_3539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13679_ clknet_leaf_134_wb_clk_i _01443_ _00044_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[33\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_14_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12024__B1 net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11378__A2 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_171_3886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08779__B1 net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_372 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10586__B1 net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold104 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1002\] vssd1
+ vssd1 vccd1 vccd1 net1597 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10050__A2 net1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold115 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1020\] vssd1
+ vssd1 vccd1 vccd1 net1608 sky130_fd_sc_hd__dlygate4sd3_1
Xhold126 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[21\] vssd1 vssd1 vccd1
+ vccd1 net1619 sky130_fd_sc_hd__dlygate4sd3_1
Xhold137 team_03_WB.instance_to_wrap.core.register_file.registers_state\[15\] vssd1
+ vssd1 vccd1 vccd1 net1630 sky130_fd_sc_hd__dlygate4sd3_1
Xhold148 _02631_ vssd1 vssd1 vccd1 vccd1 net1641 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09910_ net314 _05851_ _05429_ vssd1 vssd1 vccd1 vccd1 _05852_ sky130_fd_sc_hd__or3b_2
XFILLER_0_10_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold159 team_03_WB.instance_to_wrap.core.register_file.registers_state\[16\] vssd1
+ vssd1 vccd1 vccd1 net1652 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_10 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout606 _06294_ vssd1 vssd1 vccd1 vccd1 net606 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_42_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09841_ _02992_ _05671_ _05782_ vssd1 vssd1 vccd1 vccd1 _05783_ sky130_fd_sc_hd__o21ai_1
Xfanout617 _02842_ vssd1 vssd1 vccd1 vccd1 net617 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_1_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08400__C1 net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout628 net631 vssd1 vssd1 vccd1 vccd1 net628 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07754__A1 net1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout639 net641 vssd1 vssd1 vccd1 vccd1 net639 sky130_fd_sc_hd__clkbuf_4
X_09772_ net536 _05713_ vssd1 vssd1 vccd1 vccd1 _05714_ sky130_fd_sc_hd__nor2_1
X_06984_ _02828_ _02829_ _02925_ vssd1 vssd1 vccd1 vccd1 _02926_ sky130_fd_sc_hd__or3_2
XPHY_EDGE_ROW_13_Left_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08723_ net940 _04664_ vssd1 vssd1 vccd1 vccd1 _04665_ sky130_fd_sc_hd__or2_1
XANTENNA__11838__B1 net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07506__A1 net1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout277_A _06430_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08654_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[7\] net1009
+ net930 _04595_ vssd1 vssd1 vccd1 vccd1 _04596_ sky130_fd_sc_hd__o211a_1
XANTENNA__10510__B1 net1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07601__S1 net1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07605_ net1205 team_03_WB.instance_to_wrap.core.register_file.registers_state\[697\]
+ net887 vssd1 vssd1 vccd1 vccd1 _03547_ sky130_fd_sc_hd__and3_1
XFILLER_0_77_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08585_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[957\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[925\]
+ net967 vssd1 vssd1 vccd1 vccd1 _04527_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout444_A net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1186_A net1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07536_ net1103 team_03_WB.instance_to_wrap.core.register_file.registers_state\[198\]
+ net799 team_03_WB.instance_to_wrap.core.register_file.registers_state\[230\] net732
+ vssd1 vssd1 vccd1 vccd1 _03478_ sky130_fd_sc_hd__a221o_1
XANTENNA__08467__C1 net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1134 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07467_ net1184 team_03_WB.instance_to_wrap.core.register_file.registers_state\[725\]
+ net769 team_03_WB.instance_to_wrap.core.register_file.registers_state\[757\] net744
+ vssd1 vssd1 vccd1 vccd1 _03409_ sky130_fd_sc_hd__o221a_1
XFILLER_0_14_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout611_A net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_957 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1353_A net1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout709_A net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11005__D net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09206_ _03866_ _04072_ _05147_ net608 vssd1 vssd1 vccd1 vccd1 _05148_ sky130_fd_sc_hd__a31o_1
XPHY_EDGE_ROW_22_Left_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_40_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12015__B1 net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07690__B1 net1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07398_ net1123 _03335_ _03339_ net1138 vssd1 vssd1 vccd1 vccd1 _03340_ sky130_fd_sc_hd__a211o_1
XFILLER_0_63_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09137_ net526 _02944_ _02948_ _02952_ vssd1 vssd1 vccd1 vccd1 _05079_ sky130_fd_sc_hd__and4_1
XFILLER_0_17_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1141_X net1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10577__B1 net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1239_X net1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10041__A2 net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07442__B1 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09068_ net1064 _05009_ _05008_ vssd1 vssd1 vccd1 vccd1 _05010_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout980_A net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07993__A1 net1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout699_X net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11729__S net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08019_ net1161 _03953_ _03952_ net1146 vssd1 vssd1 vccd1 vccd1 _03961_ sky130_fd_sc_hd__o211a_1
XANTENNA__10633__S net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold660 team_03_WB.instance_to_wrap.core.register_file.registers_state\[399\] vssd1
+ vssd1 vccd1 vccd1 net2153 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_38_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold671 team_03_WB.instance_to_wrap.core.register_file.registers_state\[368\] vssd1
+ vssd1 vccd1 vccd1 net2164 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_38_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11030_ net637 _06589_ vssd1 vssd1 vccd1 vccd1 _06590_ sky130_fd_sc_hd__nor2_1
Xhold682 team_03_WB.instance_to_wrap.core.register_file.registers_state\[817\] vssd1
+ vssd1 vccd1 vccd1 net2175 sky130_fd_sc_hd__dlygate4sd3_1
Xhold693 team_03_WB.instance_to_wrap.core.register_file.registers_state\[113\] vssd1
+ vssd1 vccd1 vccd1 net2186 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07745__A1 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout866_X net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11541__A2 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08942__B1 net1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11829__B1 net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12981_ net1275 vssd1 vssd1 vccd1 vccd1 _00745_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_86_2136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14720_ clknet_leaf_50_wb_clk_i _02484_ _01085_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.decoder.inst\[17\]
+ sky130_fd_sc_hd__dfrtp_4
X_11932_ _06519_ net2743 net367 vssd1 vssd1 vccd1 vccd1 _01610_ sky130_fd_sc_hd__mux2_1
XANTENNA__10501__B1 net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11863_ _06682_ net456 net375 net1899 vssd1 vssd1 vccd1 vccd1 _01677_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_64_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14651_ clknet_leaf_121_wb_clk_i _02415_ _01016_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1005\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_157_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_157_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10814_ team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[27\] _05865_ net318 _06403_
+ net686 vssd1 vssd1 vccd1 vccd1 _06420_ sky130_fd_sc_hd__a41o_1
XFILLER_0_67_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13602_ net1304 vssd1 vssd1 vccd1 vccd1 _01366_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_0_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11794_ net2353 _06624_ net329 vssd1 vssd1 vccd1 vccd1 _01744_ sky130_fd_sc_hd__mux2_1
X_14582_ clknet_leaf_151_wb_clk_i _02346_ _00947_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[936\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_156_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_101_2450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10804__A1 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10745_ _05706_ net604 vssd1 vssd1 vccd1 vccd1 _06365_ sky130_fd_sc_hd__nand2_1
X_13533_ net1307 vssd1 vssd1 vccd1 vccd1 _01297_ sky130_fd_sc_hd__inv_2
XFILLER_0_27_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_60_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12006__A0 net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13464_ net1341 vssd1 vssd1 vccd1 vccd1 _01228_ sky130_fd_sc_hd__inv_2
XANTENNA__07681__B1 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10676_ team_03_WB.instance_to_wrap.core.pc.current_pc\[29\] _06317_ vssd1 vssd1
+ vccd1 vccd1 _06318_ sky130_fd_sc_hd__or2_1
XFILLER_0_42_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12415_ net1351 vssd1 vssd1 vccd1 vccd1 _00179_ sky130_fd_sc_hd__inv_2
XFILLER_0_51_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13395_ net1406 vssd1 vssd1 vccd1 vccd1 _01159_ sky130_fd_sc_hd__inv_2
XANTENNA__09422__A1 _04816_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07028__A3 net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10568__B1 net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12021__A3 net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10032__A2 net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12346_ net1377 vssd1 vssd1 vccd1 vccd1 _00110_ sky130_fd_sc_hd__inv_2
XANTENNA__07433__B1 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput209 net209 vssd1 vssd1 vccd1 vccd1 gpio_out[12] sky130_fd_sc_hd__buf_2
Xclkbuf_leaf_187_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_187_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08630__C1 net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15065_ net1451 vssd1 vssd1 vccd1 vccd1 la_data_out[1] sky130_fd_sc_hd__buf_2
Xclkbuf_leaf_116_wb_clk_i clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_116_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_12277_ net1271 vssd1 vssd1 vccd1 vccd1 _00041_ sky130_fd_sc_hd__inv_2
X_14016_ clknet_leaf_192_wb_clk_i _01780_ _00381_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[370\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09725__A2 _04893_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11228_ _06532_ net2338 net489 vssd1 vssd1 vccd1 vccd1 _02183_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_147_3387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11159_ net1043 net839 net299 net669 vssd1 vssd1 vccd1 vccd1 _06657_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_108_2604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_147_3398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13155__A net1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14918_ clknet_leaf_44_wb_clk_i _02673_ _01283_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_O\[5\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_125_2951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11296__A1 net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08249__A net1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11008__C_N net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15071__1457 vssd1 vssd1 vccd1 vccd1 _15071__1457/HI net1457 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_19_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14849_ clknet_leaf_82_wb_clk_i net1655 _01214_ vssd1 vssd1 vccd1 vccd1 net104 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_77_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_2859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09779__S net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08370_ _04310_ _04311_ net1219 vssd1 vssd1 vccd1 vccd1 _04312_ sky130_fd_sc_hd__o21a_1
XANTENNA__11048__B2 net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08449__C1 net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_173_3926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14982__Q team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[1\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07321_ net1185 team_03_WB.instance_to_wrap.core.register_file.registers_state\[189\]
+ vssd1 vssd1 vccd1 vccd1 _03263_ sky130_fd_sc_hd__and2_1
XFILLER_0_74_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07252_ net1176 team_03_WB.instance_to_wrap.core.register_file.registers_state\[72\]
+ net774 team_03_WB.instance_to_wrap.core.register_file.registers_state\[104\] net726
+ vssd1 vssd1 vccd1 vccd1 _03194_ sky130_fd_sc_hd__o221a_1
XFILLER_0_6_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_144_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11122__B net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07183_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[531\] net792
+ vssd1 vssd1 vccd1 vccd1 _03125_ sky130_fd_sc_hd__or2_1
XFILLER_0_131_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_30_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_30_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08134__D _03314_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10961__B net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11776__C net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout403 _06718_ vssd1 vssd1 vccd1 vccd1 net403 sky130_fd_sc_hd__clkbuf_4
Xfanout414 _06635_ vssd1 vssd1 vccd1 vccd1 net414 sky130_fd_sc_hd__clkbuf_8
Xfanout425 net426 vssd1 vssd1 vccd1 vccd1 net425 sky130_fd_sc_hd__buf_1
Xfanout436 net437 vssd1 vssd1 vccd1 vccd1 net436 sky130_fd_sc_hd__buf_2
XANTENNA__11523__A2 net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout394_A net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08924__B1 net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09824_ _05073_ _05688_ vssd1 vssd1 vccd1 vccd1 _05766_ sky130_fd_sc_hd__nand2_1
Xfanout447 _06801_ vssd1 vssd1 vccd1 vccd1 net447 sky130_fd_sc_hd__buf_6
XANTENNA_fanout1101_A net1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout458 net460 vssd1 vssd1 vccd1 vccd1 net458 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10731__B1 net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout469 net471 vssd1 vssd1 vccd1 vccd1 net469 sky130_fd_sc_hd__clkbuf_4
Xclkbuf_4_14__f_wb_clk_i clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_14__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
X_09755_ net582 _05276_ _05687_ _05696_ vssd1 vssd1 vccd1 vccd1 _05697_ sky130_fd_sc_hd__a31o_2
X_06967_ net1167 _02907_ _02908_ vssd1 vssd1 vccd1 vccd1 _02909_ sky130_fd_sc_hd__and3_1
XANTENNA__10689__A _05563_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout561_A net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12079__A3 net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06950__A2 _02888_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08706_ net435 net430 _04647_ net546 vssd1 vssd1 vccd1 vccd1 _04648_ sky130_fd_sc_hd__o31a_1
X_09686_ _03988_ _04178_ _04820_ _03985_ net1020 vssd1 vssd1 vccd1 vccd1 _05628_ sky130_fd_sc_hd__a32o_1
X_06898_ team_03_WB.instance_to_wrap.core.control_logic.instruction\[4\] _02815_ _02828_
+ _02831_ vssd1 vssd1 vccd1 vccd1 _02840_ sky130_fd_sc_hd__or4_1
XANTENNA__08159__A net1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1103 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08637_ _04573_ _04578_ net873 vssd1 vssd1 vccd1 vccd1 _04579_ sky130_fd_sc_hd__mux2_1
XFILLER_0_139_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout826_A _02819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07360__C1 net1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout447_X net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_2033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1189_X net1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11039__A1 net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_2044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08568_ net1235 team_03_WB.instance_to_wrap.core.register_file.registers_state\[221\]
+ net966 team_03_WB.instance_to_wrap.core.register_file.registers_state\[253\] net938
+ vssd1 vssd1 vccd1 vccd1 _04510_ sky130_fd_sc_hd__o221a_1
XFILLER_0_37_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_30_Left_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_1098 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07519_ net1102 team_03_WB.instance_to_wrap.core.register_file.registers_state\[838\]
+ net799 team_03_WB.instance_to_wrap.core.register_file.registers_state\[870\] net1156
+ vssd1 vssd1 vccd1 vccd1 _03461_ sky130_fd_sc_hd__a221o_1
XFILLER_0_147_650 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10628__S net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08499_ net1067 _04438_ _04439_ vssd1 vssd1 vccd1 vccd1 _04441_ sky130_fd_sc_hd__or3_1
XANTENNA__09652__B2 net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_979 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10530_ net167 net1031 net1023 net1721 vssd1 vssd1 vccd1 vccd1 _02580_ sky130_fd_sc_hd__a22o_1
XFILLER_0_36_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08860__C1 net1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11032__B net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10461_ _06043_ _06050_ _06274_ vssd1 vssd1 vccd1 vccd1 _06275_ sky130_fd_sc_hd__o21a_1
XFILLER_0_162_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_388 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12200_ net1550 vssd1 vssd1 vccd1 vccd1 _02353_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_161_174 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13180_ net1430 vssd1 vssd1 vccd1 vccd1 _00944_ sky130_fd_sc_hd__inv_2
X_10392_ _06218_ _06219_ team_03_WB.instance_to_wrap.core.pc.current_pc\[17\] net680
+ vssd1 vssd1 vccd1 vccd1 _02651_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__08612__C1 net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10871__B _06468_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout983_X net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07966__A1 net1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12131_ net1593 vssd1 vssd1 vccd1 vccd1 _02422_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__11762__A2 net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12062_ _06627_ net2574 net355 vssd1 vssd1 vccd1 vccd1 _01484_ sky130_fd_sc_hd__mux2_1
Xhold490 team_03_WB.instance_to_wrap.core.register_file.registers_state\[622\] vssd1
+ vssd1 vccd1 vccd1 net1983 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07718__A1 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11013_ net274 net703 net827 vssd1 vssd1 vccd1 vccd1 _06580_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_53_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10722__B1 net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout970 net971 vssd1 vssd1 vccd1 vccd1 net970 sky130_fd_sc_hd__clkbuf_4
Xfanout981 net994 vssd1 vssd1 vccd1 vccd1 net981 sky130_fd_sc_hd__buf_2
Xfanout992 net993 vssd1 vssd1 vccd1 vccd1 net992 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_5_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11278__A1 net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12964_ net1384 vssd1 vssd1 vccd1 vccd1 _00728_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_142_3284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_142_3295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1190 team_03_WB.instance_to_wrap.core.register_file.registers_state\[832\] vssd1
+ vssd1 vccd1 vccd1 net2683 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_103_2501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14703_ clknet_leaf_68_wb_clk_i _02467_ _01068_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.control_logic.instruction\[0\]
+ sky130_fd_sc_hd__dfrtp_4
X_11915_ _06616_ net2450 net370 vssd1 vssd1 vccd1 vccd1 _01627_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_16_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_263 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10111__B net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12895_ net1350 vssd1 vssd1 vccd1 vccd1 _00659_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11922__S net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09900__B _05841_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14634_ clknet_leaf_7_wb_clk_i _02398_ _00999_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[988\]
+ sky130_fd_sc_hd__dfstp_1
X_11846_ net279 net2096 net375 vssd1 vssd1 vccd1 vccd1 _01694_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_784 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07701__A net1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11777_ net2469 _06609_ net327 vssd1 vssd1 vccd1 vccd1 _01761_ sky130_fd_sc_hd__mux2_1
X_14565_ clknet_leaf_39_wb_clk_i _02329_ _00930_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[919\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_166_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10728_ team_03_WB.instance_to_wrap.core.pc.current_pc\[17\] _05632_ net603 vssd1
+ vssd1 vccd1 vccd1 _06356_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_834 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13516_ net1307 vssd1 vssd1 vccd1 vccd1 _01280_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14496_ clknet_leaf_192_wb_clk_i _02260_ _00861_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[850\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_344 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_832 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13447_ net1406 vssd1 vssd1 vccd1 vccd1 _01211_ sky130_fd_sc_hd__inv_2
X_10659_ team_03_WB.instance_to_wrap.core.control_logic.instruction\[2\] team_03_WB.instance_to_wrap.CPU_DAT_O\[2\]
+ net846 vssd1 vssd1 vccd1 vccd1 _02469_ sky130_fd_sc_hd__mux2_1
Xclkload13 clknet_leaf_188_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload13/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_35_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkload24 clknet_leaf_13_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload24/Y sky130_fd_sc_hd__inv_8
Xclkload35 clknet_leaf_181_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload35/Y sky130_fd_sc_hd__inv_4
XFILLER_0_106_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07406__B1 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload46 clknet_leaf_26_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload46/X sky130_fd_sc_hd__clkbuf_8
X_13378_ net1428 vssd1 vssd1 vccd1 vccd1 _01142_ sky130_fd_sc_hd__inv_2
XFILLER_0_106_591 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload57 clknet_leaf_36_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload57/Y sky130_fd_sc_hd__bufinv_16
Xclkload68 clknet_leaf_48_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload68/Y sky130_fd_sc_hd__clkinv_2
XTAP_TAPCELL_ROW_77_1957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07957__A1 net1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload79 clknet_leaf_61_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload79/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_23_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_77_1968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11753__A2 net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15117_ net1487 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[22] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_149_3427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12329_ net1253 vssd1 vssd1 vccd1 vccd1 _00093_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_149_3438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09159__B1 net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15048_ net135 vssd1 vssd1 vccd1 vccd1 net172 sky130_fd_sc_hd__clkbuf_1
XANTENNA__07709__A1 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_166_3774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08906__B1 net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_166_3785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09174__A3 net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07870_ _03808_ _03811_ net823 vssd1 vssd1 vccd1 vccd1 _03812_ sky130_fd_sc_hd__o21ai_1
XANTENNA__06917__C1 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_84_wb_clk_i clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_84_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_09540_ _05394_ _05400_ net561 vssd1 vssd1 vccd1 vccd1 _05482_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_13_wb_clk_i clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_13_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_09471_ net549 net354 _05090_ vssd1 vssd1 vccd1 vccd1 _05413_ sky130_fd_sc_hd__o21ba_1
XANTENNA__07342__C1 net1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08422_ net1228 team_03_WB.instance_to_wrap.core.register_file.registers_state\[474\]
+ net954 team_03_WB.instance_to_wrap.core.register_file.registers_state\[506\] net1210
+ vssd1 vssd1 vccd1 vccd1 _04364_ sky130_fd_sc_hd__o221a_1
XFILLER_0_116_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10492__A2 net1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10956__B net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_721 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08353_ _04294_ vssd1 vssd1 vccd1 vccd1 _04295_ sky130_fd_sc_hd__inv_2
XFILLER_0_50_1131 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10448__S net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07304_ net1089 team_03_WB.instance_to_wrap.core.register_file.registers_state\[829\]
+ net893 vssd1 vssd1 vccd1 vccd1 _03246_ sky130_fd_sc_hd__or3_1
XFILLER_0_132_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_631 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07645__B1 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08284_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[567\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[535\]
+ net963 vssd1 vssd1 vccd1 vccd1 _04226_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11441__B2 net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload7 clknet_leaf_1_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload7/Y sky130_fd_sc_hd__inv_6
XANTENNA__08842__C1 net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_94 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07235_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[648\] net796
+ net746 _03176_ vssd1 vssd1 vccd1 vccd1 _03177_ sky130_fd_sc_hd__o211a_1
XFILLER_0_26_180 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1051_A net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout407_A _06717_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1149_A net1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07166_ team_03_WB.instance_to_wrap.core.decoder.inst\[19\] _02821_ _03107_ vssd1
+ vssd1 vccd1 vccd1 _03108_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_70_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_25_wb_clk_i_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__08442__A net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07984__C net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11744__A2 net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10183__S net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_183 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07097_ net1099 team_03_WB.instance_to_wrap.core.register_file.registers_state\[961\]
+ net801 team_03_WB.instance_to_wrap.core.register_file.registers_state\[993\] net1134
+ vssd1 vssd1 vccd1 vccd1 _03039_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_140_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09972__S net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1209 team_03_WB.instance_to_wrap.core.decoder.inst\[18\] vssd1 vssd1 vccd1
+ vccd1 net1209 sky130_fd_sc_hd__buf_4
XANTENNA_fanout776_A net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout397_X net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1104_X net1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08373__A1 net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout266 _06557_ vssd1 vssd1 vccd1 vccd1 net266 sky130_fd_sc_hd__buf_2
X_09807_ _05268_ _05747_ _05748_ net595 vssd1 vssd1 vccd1 vccd1 _05749_ sky130_fd_sc_hd__a211oi_1
Xfanout277 _06430_ vssd1 vssd1 vccd1 vccd1 net277 sky130_fd_sc_hd__buf_2
Xfanout288 net289 vssd1 vssd1 vccd1 vccd1 net288 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout564_X net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout943_A net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07999_ net813 _03939_ _03940_ net820 vssd1 vssd1 vccd1 vccd1 _03941_ sky130_fd_sc_hd__o211a_1
Xfanout299 _06487_ vssd1 vssd1 vccd1 vccd1 net299 sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_105_Left_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09738_ net540 _05679_ vssd1 vssd1 vccd1 vccd1 _05680_ sky130_fd_sc_hd__nand2_1
XFILLER_0_9_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08125__A1 net1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11027__B net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout731_X net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09873__A1 net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09669_ net594 _05598_ _05599_ _05610_ vssd1 vssd1 vccd1 vccd1 _05611_ sky130_fd_sc_hd__o31ai_2
XFILLER_0_16_1015 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout829_X net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09873__B2 net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11742__S net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_211 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11700_ _06742_ net383 net340 net2051 vssd1 vssd1 vccd1 vccd1 _01834_ sky130_fd_sc_hd__a22o_1
XANTENNA__10483__A2 net1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12680_ net1291 vssd1 vssd1 vccd1 vccd1 _00444_ sky130_fd_sc_hd__inv_2
XFILLER_0_139_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11631_ _06705_ net383 net348 net2518 vssd1 vssd1 vccd1 vccd1 _01901_ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_64_wb_clk_i_A clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09086__C1 net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11043__A net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_145_Right_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11432__A1 net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14350_ clknet_leaf_131_wb_clk_i _02114_ _00715_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[704\]
+ sky130_fd_sc_hd__dfrtp_1
X_11562_ net2431 net485 _06795_ net514 vssd1 vssd1 vccd1 vccd1 _01961_ sky130_fd_sc_hd__a22o_1
XFILLER_0_163_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10513_ net154 net1033 net1025 net1837 vssd1 vssd1 vccd1 vccd1 _02597_ sky130_fd_sc_hd__a22o_1
X_13301_ net1322 vssd1 vssd1 vccd1 vccd1 _01065_ sky130_fd_sc_hd__inv_2
XFILLER_0_80_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14281_ clknet_leaf_116_wb_clk_i _02045_ _00646_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[635\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_135_675 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11493_ _06614_ net2710 net391 vssd1 vssd1 vccd1 vccd1 _02013_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_98_2382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_2393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08623__Y _04565_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13232_ net1413 vssd1 vssd1 vccd1 vccd1 _00996_ sky130_fd_sc_hd__inv_2
XFILLER_0_122_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10444_ net285 _06136_ _06261_ net682 vssd1 vssd1 vccd1 vccd1 _06262_ sky130_fd_sc_hd__o31ai_1
XANTENNA__09448__A net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input72_A wbs_adr_i[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_1085 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07939__A1 net1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13163_ net1287 vssd1 vssd1 vccd1 vccd1 _00927_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_55_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15070__1456 vssd1 vssd1 vccd1 vccd1 _15070__1456/HI net1456 sky130_fd_sc_hd__conb_1
X_10375_ team_03_WB.instance_to_wrap.core.pc.current_pc\[20\] net677 _06203_ _06205_
+ vssd1 vssd1 vccd1 vccd1 _02654_ sky130_fd_sc_hd__o22a_1
XFILLER_0_0_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07403__A3 net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12114_ net1142 net1845 _06292_ net1145 vssd1 vssd1 vccd1 vccd1 _00006_ sky130_fd_sc_hd__a22o_1
XFILLER_0_130_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13094_ net1299 vssd1 vssd1 vccd1 vccd1 _00858_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_72_1854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11917__S net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_1865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12045_ _06614_ net2730 net357 vssd1 vssd1 vccd1 vccd1 _01501_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_144_3324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_28 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12602__A net1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_144_3335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09183__A net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_161_3671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1132 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_161_3682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10122__A _03640_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13996_ clknet_leaf_21_wb_clk_i _01760_ _00361_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[350\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12040__C _06463_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09911__A _05757_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12947_ net1261 vssd1 vssd1 vccd1 vccd1 _00711_ sky130_fd_sc_hd__inv_2
XANTENNA__07324__C1 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_723 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09864__B2 _02945_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11652__S net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11671__A1 net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12878_ net1269 vssd1 vssd1 vccd1 vccd1 _00642_ sky130_fd_sc_hd__inv_2
XFILLER_0_157_244 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09122__S net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14617_ clknet_leaf_176_wb_clk_i _02381_ _00982_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[971\]
+ sky130_fd_sc_hd__dfstp_1
X_11829_ _06663_ net465 net325 net1943 vssd1 vssd1 vccd1 vccd1 _01710_ sky130_fd_sc_hd__a22o_1
XANTENNA__09077__C1 net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_157_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08824__C1 net1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14548_ clknet_leaf_123_wb_clk_i _02312_ _00913_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[902\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_112_Right_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_131_wb_clk_i clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_131_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_126_686 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload102 clknet_leaf_149_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload102/Y sky130_fd_sc_hd__clkinv_2
X_14479_ clknet_leaf_138_wb_clk_i _02243_ _00844_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[833\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkload113 clknet_leaf_121_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload113/Y sky130_fd_sc_hd__clkinv_2
X_07020_ net1099 team_03_WB.instance_to_wrap.core.register_file.registers_state\[547\]
+ net897 vssd1 vssd1 vccd1 vccd1 _02962_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_116_2758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload124 clknet_leaf_137_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload124/Y sky130_fd_sc_hd__inv_6
XFILLER_0_30_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload135 clknet_leaf_128_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload135/Y sky130_fd_sc_hd__clkinv_8
Xclkload146 clknet_leaf_111_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload146/Y sky130_fd_sc_hd__clkinv_2
XANTENNA__11187__B1 net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload157 clknet_leaf_99_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload157/Y sky130_fd_sc_hd__inv_6
XPHY_EDGE_ROW_49_Right_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08278__S1 net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_168_3814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload168 clknet_leaf_129_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload168/Y sky130_fd_sc_hd__clkinvlp_4
XTAP_TAPCELL_ROW_168_3825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload179 clknet_leaf_96_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload179/Y sky130_fd_sc_hd__inv_6
XFILLER_0_51_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08052__B1 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09645__X _05587_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_367 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08971_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[553\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[521\]
+ net988 vssd1 vssd1 vccd1 vccd1 _04913_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_109_wb_clk_i_A clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_07922_ net1237 net1015 _03107_ vssd1 vssd1 vccd1 vccd1 _03864_ sky130_fd_sc_hd__a21oi_4
Xhold19 team_03_WB.instance_to_wrap.core.register_file.registers_state\[969\] vssd1
+ vssd1 vccd1 vccd1 net1512 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09001__C1 net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07158__A2 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1020 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07853_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[955\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[923\]
+ net783 vssd1 vssd1 vccd1 vccd1 _03795_ sky130_fd_sc_hd__mux2_1
XANTENNA__07606__A net1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08201__S net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07563__C1 net1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07784_ _03700_ _03701_ _03722_ net617 vssd1 vssd1 vccd1 vccd1 _03726_ sky130_fd_sc_hd__o211a_2
XPHY_EDGE_ROW_58_Right_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09523_ _05372_ _05376_ net562 vssd1 vssd1 vccd1 vccd1 _05465_ sky130_fd_sc_hd__mux2_1
XFILLER_0_149_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13343__A net1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout357_A _06818_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09881__D_N _05646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09454_ _05394_ _05395_ net555 vssd1 vssd1 vccd1 vccd1 _05396_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout1099_A net1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_412 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09032__S net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08405_ net1208 _04343_ _04346_ vssd1 vssd1 vccd1 vccd1 _04347_ sky130_fd_sc_hd__or3_1
X_09385_ _04267_ _05326_ vssd1 vssd1 vccd1 vccd1 _05327_ sky130_fd_sc_hd__nor2_1
XANTENNA__10870__C1 net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout524_A _06322_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1057 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1266_A net1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_163_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08336_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[1013\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[981\]
+ net969 vssd1 vssd1 vccd1 vccd1 _04278_ sky130_fd_sc_hd__mux2_1
XANTENNA__07618__B1 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08815__C1 net1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11414__B2 net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_962 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08267_ net432 _04079_ _04207_ net543 vssd1 vssd1 vccd1 vccd1 _04209_ sky130_fd_sc_hd__o31a_1
XANTENNA__07094__B2 net1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout312_X net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_148_wb_clk_i_A clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout1054_X net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_67_Right_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07218_ net1171 team_03_WB.instance_to_wrap.core.register_file.registers_state\[850\]
+ net757 team_03_WB.instance_to_wrap.core.register_file.registers_state\[882\] net1123
+ vssd1 vssd1 vccd1 vccd1 _03160_ sky130_fd_sc_hd__o221a_1
X_08198_ net935 _04138_ _04139_ net855 vssd1 vssd1 vccd1 vccd1 _04140_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout893_A net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07149_ net810 _03086_ _03089_ _03090_ vssd1 vssd1 vccd1 vccd1 _03091_ sky130_fd_sc_hd__a22o_1
XFILLER_0_30_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1221_X net1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07397__A2 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_2290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10160_ _03679_ _06000_ _06001_ vssd1 vssd1 vccd1 vccd1 _06002_ sky130_fd_sc_hd__nor3_2
XANTENNA_fanout681_X net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1006 net1008 vssd1 vssd1 vccd1 vccd1 net1006 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11737__S net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10091_ _05583_ _05596_ _05821_ _05934_ vssd1 vssd1 vccd1 vccd1 _05935_ sky130_fd_sc_hd__and4b_1
XANTENNA__10641__S net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1028 net1029 vssd1 vssd1 vccd1 vccd1 net1028 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_50_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1039 net1040 vssd1 vssd1 vccd1 vccd1 net1039 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_50_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08346__A1 net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout946_X net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11350__B1 net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_76_Right_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11038__A net1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13850_ clknet_leaf_141_wb_clk_i _01614_ _00215_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[204\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09731__A net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12801_ net1272 vssd1 vssd1 vccd1 vccd1 _00565_ sky130_fd_sc_hd__inv_2
X_10993_ net2278 net420 _06568_ net499 vssd1 vssd1 vccd1 vccd1 _02303_ sky130_fd_sc_hd__a22o_1
X_13781_ clknet_leaf_126_wb_clk_i _01545_ _00146_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[135\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07306__C1 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07857__B1 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11653__A1 _06619_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12732_ net1418 vssd1 vssd1 vccd1 vccd1 _00496_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_48_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_187_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12663_ net1386 vssd1 vssd1 vccd1 vccd1 _00427_ sky130_fd_sc_hd__inv_2
XFILLER_0_132_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14402_ clknet_leaf_185_wb_clk_i _02166_ _00767_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[756\]
+ sky130_fd_sc_hd__dfrtp_1
X_11614_ _06688_ net379 net346 net2519 vssd1 vssd1 vccd1 vccd1 _01918_ sky130_fd_sc_hd__a22o_1
XANTENNA__10883__Y _06479_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12594_ net1395 vssd1 vssd1 vccd1 vccd1 _00358_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_137_3183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_85_Right_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_137_3194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14333_ clknet_leaf_26_wb_clk_i _02097_ _00698_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[687\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_135_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11545_ net2071 net482 _06788_ net501 vssd1 vssd1 vccd1 vccd1 _01971_ sky130_fd_sc_hd__a22o_1
XANTENNA__08821__A2 net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_196 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14264_ clknet_leaf_3_wb_clk_i _02028_ _00629_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[618\]
+ sky130_fd_sc_hd__dfrtp_1
X_11476_ net2560 net394 _06773_ net514 vssd1 vssd1 vccd1 vccd1 _02025_ sky130_fd_sc_hd__a22o_1
XFILLER_0_111_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11708__A2 net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10427_ net304 net303 _06063_ _06247_ vssd1 vssd1 vccd1 vccd1 _06248_ sky130_fd_sc_hd__a211o_1
XFILLER_0_150_464 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13215_ net1347 vssd1 vssd1 vccd1 vccd1 _00979_ sky130_fd_sc_hd__inv_2
XANTENNA__11220__B _06503_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_1905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14195_ clknet_leaf_99_wb_clk_i _01959_ _00560_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[549\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_110_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10916__B1 net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10358_ net283 _06148_ _06186_ net679 vssd1 vssd1 vccd1 vccd1 _06192_ sky130_fd_sc_hd__o31a_1
XANTENNA__09906__A _05596_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_2655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13146_ net1377 vssd1 vssd1 vccd1 vccd1 _00910_ sky130_fd_sc_hd__inv_2
XANTENNA__08810__A net1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10392__B2 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11647__S net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07793__C1 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13077_ net1275 vssd1 vssd1 vccd1 vccd1 _00841_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_163_3722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10289_ _05963_ _06128_ _06130_ vssd1 vssd1 vccd1 vccd1 _06131_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_57_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_94_Right_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07426__A net1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12028_ _06770_ net466 net361 net2568 vssd1 vssd1 vccd1 vccd1 _01517_ sky130_fd_sc_hd__a22o_1
XFILLER_0_73_13 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11892__A1 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10787__A net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13979_ clknet_leaf_123_wb_clk_i _01743_ _00344_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[333\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_654 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07848__A0 _03788_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09170_ net436 net428 _04922_ net546 vssd1 vssd1 vccd1 vccd1 _05112_ sky130_fd_sc_hd__o31a_1
XFILLER_0_28_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_916 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_118_2809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09696__S0 net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08121_ net1087 team_03_WB.instance_to_wrap.core.register_file.registers_state\[826\]
+ net892 vssd1 vssd1 vccd1 vccd1 _04063_ sky130_fd_sc_hd__or3_1
XFILLER_0_83_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_161_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07076__A1 net1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08273__B1 net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09470__C1 net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_494 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08052_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[150\] net772
+ net738 _03993_ vssd1 vssd1 vccd1 vccd1 _03994_ sky130_fd_sc_hd__a211o_1
XFILLER_0_114_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_1080 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07003_ _02838_ _02928_ _02935_ _02832_ vssd1 vssd1 vccd1 vccd1 _02945_ sky130_fd_sc_hd__o211a_1
XFILLER_0_40_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11580__A0 net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07784__C1 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13338__A net1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08954_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[41\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[9\]
+ net991 vssd1 vssd1 vccd1 vccd1 _04896_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout1014_A _02869_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07336__A team_03_WB.instance_to_wrap.core.decoder.inst\[31\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07905_ net1187 team_03_WB.instance_to_wrap.core.register_file.registers_state\[559\]
+ net877 vssd1 vssd1 vccd1 vccd1 _03847_ sky130_fd_sc_hd__and3_1
X_08885_ net544 _04825_ _04772_ net561 vssd1 vssd1 vccd1 vccd1 _04827_ sky130_fd_sc_hd__a211o_1
XANTENNA__08423__S1 net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07536__C1 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout474_A net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07836_ net1082 team_03_WB.instance_to_wrap.core.register_file.registers_state\[970\]
+ net791 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1002\] net1123
+ vssd1 vssd1 vccd1 vccd1 _03778_ sky130_fd_sc_hd__a221o_1
XANTENNA__11883__A1 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07551__A2 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout641_A _06458_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07767_ net1194 team_03_WB.instance_to_wrap.core.register_file.registers_state\[588\]
+ vssd1 vssd1 vccd1 vccd1 _03709_ sky130_fd_sc_hd__or2_1
XFILLER_0_17_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout739_A net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13073__A net1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09506_ _04778_ _05441_ _05444_ _05446_ vssd1 vssd1 vccd1 vccd1 _05448_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_39_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07698_ net684 _03639_ vssd1 vssd1 vccd1 vccd1 _03640_ sky130_fd_sc_hd__and2b_2
XFILLER_0_78_175 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08500__A1 net1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09437_ _04566_ _04680_ vssd1 vssd1 vccd1 vccd1 _05379_ sky130_fd_sc_hd__nor2_1
XFILLER_0_66_348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10984__X _06562_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout906_A _06285_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout527_X net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1171_X net1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09368_ _05176_ _05181_ _05309_ _05177_ vssd1 vssd1 vccd1 vccd1 _05310_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_23_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11399__A0 net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11024__C net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_286 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_164_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08319_ net1048 team_03_WB.instance_to_wrap.core.register_file.registers_state\[664\]
+ net999 team_03_WB.instance_to_wrap.core.register_file.registers_state\[696\] net929
+ vssd1 vssd1 vccd1 vccd1 _04261_ sky130_fd_sc_hd__a221o_1
XANTENNA__10636__S net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09299_ _04619_ _05238_ vssd1 vssd1 vccd1 vccd1 _05241_ sky130_fd_sc_hd__and2_1
XFILLER_0_90_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_554 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1436_X net1436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_2330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11330_ _06632_ net2688 net406 vssd1 vssd1 vccd1 vccd1 _02115_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout896_X net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_3080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11261_ net709 _06473_ net827 vssd1 vssd1 vccd1 vccd1 _06698_ sky130_fd_sc_hd__and3_1
XANTENNA__11040__B net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_3091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_2238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08567__A1 net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_2249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10212_ _06037_ _06053_ vssd1 vssd1 vccd1 vccd1 _06054_ sky130_fd_sc_hd__nand2_1
X_13000_ net1290 vssd1 vssd1 vccd1 vccd1 _00764_ sky130_fd_sc_hd__inv_2
XFILLER_0_30_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11192_ net1043 net839 _06545_ net669 vssd1 vssd1 vccd1 vccd1 _06677_ sky130_fd_sc_hd__and4_1
XFILLER_0_24_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08662__S1 net1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10143_ _04148_ net672 _05984_ vssd1 vssd1 vccd1 vccd1 _05985_ sky130_fd_sc_hd__o21ai_1
XANTENNA__08319__A1 net1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input35_A gpio_in[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10074_ _05917_ vssd1 vssd1 vccd1 vccd1 _05918_ sky130_fd_sc_hd__inv_2
X_14951_ clknet_leaf_104_wb_clk_i _02703_ _01316_ vssd1 vssd1 vccd1 vccd1 net234 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11323__A0 _06519_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13902_ clknet_leaf_126_wb_clk_i _01666_ _00267_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[256\]
+ sky130_fd_sc_hd__dfrtp_1
X_14882_ clknet_leaf_81_wb_clk_i _02645_ _01247_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.pc.current_pc\[11\]
+ sky130_fd_sc_hd__dfrtp_2
X_13833_ clknet_leaf_71_wb_clk_i _01597_ _00198_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[187\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09819__A1 net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_67_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13764_ clknet_leaf_29_wb_clk_i _01528_ _00129_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[118\]
+ sky130_fd_sc_hd__dfrtp_1
X_10976_ net692 _05142_ _02932_ vssd1 vssd1 vccd1 vccd1 _06555_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_57_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_139_3223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_139_3234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12715_ net1287 vssd1 vssd1 vccd1 vccd1 _00479_ sky130_fd_sc_hd__inv_2
XFILLER_0_31_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13695_ clknet_leaf_21_wb_clk_i _01459_ _00060_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[49\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11930__S net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12646_ net1363 vssd1 vssd1 vccd1 vccd1 _00410_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_156_3570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_156_3581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08805__A net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12577_ net1281 vssd1 vssd1 vccd1 vccd1 _00341_ sky130_fd_sc_hd__inv_2
XFILLER_0_108_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14316_ clknet_leaf_17_wb_clk_i _02080_ _00681_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[670\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_151_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_152_3489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_954 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11528_ net491 net619 _06640_ net482 net1789 vssd1 vssd1 vccd1 vccd1 _01982_ sky130_fd_sc_hd__a32o_1
XFILLER_0_151_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_113_2706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold308 team_03_WB.instance_to_wrap.core.register_file.registers_state\[883\] vssd1
+ vssd1 vccd1 vccd1 net1801 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold319 net111 vssd1 vssd1 vccd1 vccd1 net1812 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14247_ clknet_leaf_107_wb_clk_i _02011_ _00612_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[601\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_150_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11459_ net2437 net392 _06766_ net495 vssd1 vssd1 vccd1 vccd1 _02035_ sky130_fd_sc_hd__a22o_1
XFILLER_0_22_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08102__S0 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14178_ clknet_leaf_185_wb_clk_i _01942_ _00543_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[532\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13158__A net1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13129_ net1253 vssd1 vssd1 vccd1 vccd1 _00893_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1008 team_03_WB.instance_to_wrap.core.register_file.registers_state\[587\] vssd1
+ vssd1 vccd1 vccd1 net2501 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11314__A0 _06479_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12997__A net1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1019 team_03_WB.instance_to_wrap.core.register_file.registers_state\[208\] vssd1
+ vssd1 vccd1 vccd1 net2512 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout1370 net1437 vssd1 vssd1 vccd1 vccd1 net1370 sky130_fd_sc_hd__buf_2
X_08670_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[551\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[519\]
+ net990 vssd1 vssd1 vccd1 vccd1 _04612_ sky130_fd_sc_hd__mux2_1
Xfanout1381 net1393 vssd1 vssd1 vccd1 vccd1 net1381 sky130_fd_sc_hd__clkbuf_4
Xfanout1392 net1393 vssd1 vssd1 vccd1 vccd1 net1392 sky130_fd_sc_hd__buf_4
XANTENNA__09371__A _04382_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14985__Q team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[4\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07621_ net724 _03562_ _03546_ _03538_ vssd1 vssd1 vccd1 vccd1 _03563_ sky130_fd_sc_hd__o2bb2a_4
XFILLER_0_36_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07552_ net1200 team_03_WB.instance_to_wrap.core.register_file.registers_state\[184\]
+ vssd1 vssd1 vccd1 vccd1 _03494_ sky130_fd_sc_hd__and2_1
XANTENNA__12001__S net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10825__C1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07297__A1 net1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07483_ _03407_ _03408_ _03416_ _03424_ vssd1 vssd1 vccd1 vccd1 _03425_ sky130_fd_sc_hd__o22a_4
XFILLER_0_159_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_71 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09222_ _04503_ _05163_ vssd1 vssd1 vccd1 vccd1 _05164_ sky130_fd_sc_hd__nor2_1
XFILLER_0_29_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09153_ net547 _04384_ _05094_ vssd1 vssd1 vccd1 vccd1 _05095_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_146_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09994__A0 _05879_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_792 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08797__A1 net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08104_ net1114 _04042_ _04043_ vssd1 vssd1 vccd1 vccd1 _04046_ sky130_fd_sc_hd__or3_1
XANTENNA__11141__A net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06880__D team_03_WB.instance_to_wrap.core.decoder.inst\[31\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09084_ net1221 _05024_ _05025_ vssd1 vssd1 vccd1 vccd1 _05026_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_142_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08035_ _03974_ _03976_ net1161 vssd1 vssd1 vccd1 vccd1 _03977_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_4_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold820 team_03_WB.instance_to_wrap.core.register_file.registers_state\[803\] vssd1
+ vssd1 vccd1 vccd1 net2313 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput80 wbs_adr_i[21] vssd1 vssd1 vccd1 vccd1 net80 sky130_fd_sc_hd__buf_1
Xinput91 wbs_adr_i[31] vssd1 vssd1 vccd1 vccd1 net91 sky130_fd_sc_hd__buf_1
XANTENNA_fanout1131_A net1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold831 team_03_WB.instance_to_wrap.core.register_file.registers_state\[213\] vssd1
+ vssd1 vccd1 vccd1 net2324 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08549__A1 net1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold842 team_03_WB.instance_to_wrap.core.register_file.registers_state\[557\] vssd1
+ vssd1 vccd1 vccd1 net2335 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1229_A net1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold853 team_03_WB.instance_to_wrap.core.register_file.registers_state\[232\] vssd1
+ vssd1 vccd1 vccd1 net2346 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold864 team_03_WB.instance_to_wrap.core.register_file.registers_state\[319\] vssd1
+ vssd1 vccd1 vccd1 net2357 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold875 team_03_WB.instance_to_wrap.core.register_file.registers_state\[524\] vssd1
+ vssd1 vccd1 vccd1 net2368 sky130_fd_sc_hd__dlygate4sd3_1
Xhold886 team_03_WB.instance_to_wrap.core.register_file.registers_state\[789\] vssd1
+ vssd1 vccd1 vccd1 net2379 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07337__Y _03279_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold897 team_03_WB.instance_to_wrap.core.register_file.registers_state\[135\] vssd1
+ vssd1 vccd1 vccd1 net2390 sky130_fd_sc_hd__dlygate4sd3_1
X_09986_ _05871_ net228 net289 vssd1 vssd1 vccd1 vccd1 _02728_ sky130_fd_sc_hd__mux2_1
XANTENNA__09980__S net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10108__A1 _04770_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08937_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[939\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[907\]
+ net961 vssd1 vssd1 vccd1 vccd1 _04879_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout856_A net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout477_X net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07509__C1 net1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08868_ _02937_ net544 net556 vssd1 vssd1 vccd1 vccd1 _04810_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11019__C _06478_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09281__A net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07819_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[10\] net791
+ net726 _03760_ vssd1 vssd1 vccd1 vccd1 _03761_ sky130_fd_sc_hd__o211a_1
X_08799_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[33\] net983
+ vssd1 vssd1 vccd1 vccd1 _04741_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout644_X net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10830_ team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[24\] net305 _06432_ net691
+ vssd1 vssd1 vccd1 vccd1 _06433_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_79_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_45_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07288__A1 net1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11035__B _06503_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10761_ net524 _06373_ _06374_ net529 net1679 vssd1 vssd1 vccd1 vccd1 _02437_ sky130_fd_sc_hd__a32o_1
XANTENNA__07232__C net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout811_X net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout909_X net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12500_ net1304 vssd1 vssd1 vccd1 vccd1 _00264_ sky130_fd_sc_hd__inv_2
X_13480_ net1406 vssd1 vssd1 vccd1 vccd1 _01244_ sky130_fd_sc_hd__inv_2
X_10692_ net602 _06313_ _06329_ _06331_ vssd1 vssd1 vccd1 vccd1 _06332_ sky130_fd_sc_hd__a31oi_1
XANTENNA__10831__A2 _06433_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_510 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_3120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12431_ net1394 vssd1 vssd1 vccd1 vccd1 _00195_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_134_3131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09985__A0 _05870_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08332__S0 net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11051__A net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12362_ net1285 vssd1 vssd1 vccd1 vccd1 _00126_ sky130_fd_sc_hd__inv_2
XFILLER_0_22_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_130_3039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14101_ clknet_leaf_129_wb_clk_i _01865_ _00466_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[455\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07996__C1 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11313_ _06621_ net2713 net404 vssd1 vssd1 vccd1 vccd1 _02132_ sky130_fd_sc_hd__mux2_1
XANTENNA__07460__A1 net1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15081_ net1467 vssd1 vssd1 vccd1 vccd1 la_data_out[17] sky130_fd_sc_hd__buf_2
XFILLER_0_22_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12293_ net1353 vssd1 vssd1 vccd1 vccd1 _00057_ sky130_fd_sc_hd__inv_2
XFILLER_0_50_568 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14032_ clknet_leaf_160_wb_clk_i _01796_ _00397_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[386\]
+ sky130_fd_sc_hd__dfrtp_1
X_11244_ net512 net640 _06689_ net411 net2038 vssd1 vssd1 vccd1 vccd1 _02173_ sky130_fd_sc_hd__a32o_1
XANTENNA__08360__A net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_18 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07212__A1 net1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11175_ net694 net714 net296 vssd1 vssd1 vccd1 vccd1 _06667_ sky130_fd_sc_hd__or3b_1
XFILLER_0_101_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10126_ _03279_ _05966_ _05967_ vssd1 vssd1 vccd1 vccd1 _05968_ sky130_fd_sc_hd__and3_1
XANTENNA__08960__A1 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07763__A2 net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06971__B1 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11925__S net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14934_ clknet_leaf_51_wb_clk_i _02689_ _01299_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_O\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_10057_ net30 net1036 net909 net2714 vssd1 vssd1 vccd1 vccd1 _02674_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_69_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08173__C1 net1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07263__X _03205_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14865_ clknet_leaf_63_wb_clk_i net1678 _01230_ vssd1 vssd1 vccd1 vccd1 net121 sky130_fd_sc_hd__dfrtp_1
XANTENNA__10093__B_N _05676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_2543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkload0_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13816_ clknet_leaf_19_wb_clk_i _01580_ _00181_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[170\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_158_3610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14796_ clknet_leaf_89_wb_clk_i _02560_ _01161_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_I\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_158_3621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07279__A1 net1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13747_ clknet_leaf_102_wb_clk_i _01511_ _00112_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[101\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07142__C net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10959_ _06538_ _06539_ _06540_ _06399_ vssd1 vssd1 vccd1 vccd1 _06541_ sky130_fd_sc_hd__o211a_4
XANTENNA__11660__S net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_154_3529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08535__A _04476_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13678_ clknet_leaf_124_wb_clk_i _01442_ _00043_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[32\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_14_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_4_2__f_wb_clk_i_A clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_375 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08228__B1 net1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12629_ net1292 vssd1 vssd1 vccd1 vccd1 _00393_ sky130_fd_sc_hd__inv_2
XANTENNA__09425__C1 net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_171_3876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10035__B1 net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09976__A0 _02888_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08779__A1 net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_660 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_171_3887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_38_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_38_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_53_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07987__C1 net1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10586__B2 _03023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold105 team_03_WB.instance_to_wrap.core.register_file.registers_state\[21\] vssd1
+ vssd1 vccd1 vccd1 net1598 sky130_fd_sc_hd__dlygate4sd3_1
Xhold116 team_03_WB.instance_to_wrap.core.register_file.registers_state\[973\] vssd1
+ vssd1 vccd1 vccd1 net1609 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_145_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold127 _02520_ vssd1 vssd1 vccd1 vccd1 net1620 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold138 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[4\] vssd1 vssd1 vccd1
+ vccd1 net1631 sky130_fd_sc_hd__dlygate4sd3_1
Xhold149 team_03_WB.instance_to_wrap.ADR_I\[19\] vssd1 vssd1 vccd1 vccd1 net1642 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08270__A net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_22 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09840_ net568 _05447_ _05439_ net574 vssd1 vssd1 vccd1 vccd1 _05782_ sky130_fd_sc_hd__a211o_1
Xfanout607 net609 vssd1 vssd1 vccd1 vccd1 net607 sky130_fd_sc_hd__clkbuf_4
Xfanout618 net621 vssd1 vssd1 vccd1 vccd1 net618 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08400__B1 net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout629 net631 vssd1 vssd1 vccd1 vccd1 net629 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_0_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08951__A1 net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_13__f_wb_clk_i clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_13__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
X_09771_ _03208_ _04646_ vssd1 vssd1 vccd1 vccd1 _05713_ sky130_fd_sc_hd__nand2_1
XFILLER_0_95_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06983_ _02806_ _02810_ vssd1 vssd1 vccd1 vccd1 _02925_ sky130_fd_sc_hd__nand2_2
XANTENNA__06996__Y _02938_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08722_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[548\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[516\]
+ net977 vssd1 vssd1 vccd1 vccd1 _04664_ sky130_fd_sc_hd__mux2_1
X_08653_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[39\] net990
+ vssd1 vssd1 vccd1 vccd1 _04595_ sky130_fd_sc_hd__or2_1
XFILLER_0_96_719 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07604_ net825 _03545_ net724 vssd1 vssd1 vccd1 vccd1 _03546_ sky130_fd_sc_hd__a21o_1
XANTENNA__11136__A net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08584_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[829\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[797\]
+ net967 vssd1 vssd1 vccd1 vccd1 _04526_ sky130_fd_sc_hd__mux2_1
XFILLER_0_113_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_646 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07535_ net1103 team_03_WB.instance_to_wrap.core.register_file.registers_state\[70\]
+ net799 team_03_WB.instance_to_wrap.core.register_file.registers_state\[102\] net747
+ vssd1 vssd1 vccd1 vccd1 _03477_ sky130_fd_sc_hd__a221o_1
XFILLER_0_165_117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07809__A3 net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_819 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1081_A _02788_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1179_A net1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10813__A2 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07466_ net822 _03401_ net720 vssd1 vssd1 vccd1 vccd1 _03408_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_63_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_174_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09205_ net526 _03491_ _04074_ _05144_ vssd1 vssd1 vccd1 vccd1 _05147_ sky130_fd_sc_hd__and4_2
XTAP_TAPCELL_ROW_40_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_146_375 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07397_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[927\] net791
+ _03334_ net1149 vssd1 vssd1 vccd1 vccd1 _03339_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout604_A net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1346_A net1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09975__S net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09136_ net583 _05076_ vssd1 vssd1 vccd1 vccd1 _05078_ sky130_fd_sc_hd__nand2_1
XFILLER_0_44_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_971 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11774__B1 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07442__A1 net1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09067_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[943\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[911\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[815\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[783\]
+ net985 net921 vssd1 vssd1 vccd1 vccd1 _05009_ sky130_fd_sc_hd__mux4_1
XFILLER_0_20_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1134_X net1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08018_ net729 _03957_ _03959_ net1161 vssd1 vssd1 vccd1 vccd1 _03960_ sky130_fd_sc_hd__a211o_1
Xhold650 team_03_WB.instance_to_wrap.core.register_file.registers_state\[171\] vssd1
+ vssd1 vccd1 vccd1 net2143 sky130_fd_sc_hd__dlygate4sd3_1
Xhold661 team_03_WB.instance_to_wrap.core.ru.prev_busy vssd1 vssd1 vccd1 vccd1 net2154
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout594_X net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout973_A net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold672 team_03_WB.instance_to_wrap.core.register_file.registers_state\[32\] vssd1
+ vssd1 vccd1 vccd1 net2165 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold683 team_03_WB.instance_to_wrap.core.register_file.registers_state\[262\] vssd1
+ vssd1 vccd1 vccd1 net2176 sky130_fd_sc_hd__dlygate4sd3_1
Xhold694 team_03_WB.instance_to_wrap.core.register_file.registers_state\[914\] vssd1
+ vssd1 vccd1 vccd1 net2187 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1301_X net1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09969_ _03241_ net662 vssd1 vssd1 vccd1 vccd1 _05889_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout761_X net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout859_X net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09723__B _04893_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12980_ net1306 vssd1 vssd1 vccd1 vccd1 _00744_ sky130_fd_sc_hd__inv_2
XANTENNA__10869__B _05833_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07083__X _03025_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11931_ _06628_ net2620 net370 vssd1 vssd1 vccd1 vccd1 _01611_ sky130_fd_sc_hd__mux2_1
XANTENNA__11046__A net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14650_ clknet_leaf_148_wb_clk_i _02414_ _01015_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1004\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_24_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11862_ _06499_ net2190 net377 vssd1 vssd1 vccd1 vccd1 _01678_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13601_ net1307 vssd1 vssd1 vccd1 vccd1 _01365_ sky130_fd_sc_hd__inv_2
XANTENNA__08058__C net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10813_ _05866_ net316 _06404_ team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[27\]
+ vssd1 vssd1 vccd1 vccd1 _06419_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_0_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14581_ clknet_leaf_107_wb_clk_i _02345_ _00946_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[935\]
+ sky130_fd_sc_hd__dfstp_1
X_11793_ net2201 _06623_ net328 vssd1 vssd1 vccd1 vccd1 _01745_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_2451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13532_ net1307 vssd1 vssd1 vccd1 vccd1 _01296_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_60_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10744_ team_03_WB.instance_to_wrap.core.pc.current_pc\[9\] net604 vssd1 vssd1 vccd1
+ vccd1 _06364_ sky130_fd_sc_hd__or2_1
XANTENNA__10804__A2 _05563_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_446 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13463_ net1328 vssd1 vssd1 vccd1 vccd1 _01227_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_11_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07681__A1 net1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10675_ team_03_WB.instance_to_wrap.core.pc.current_pc\[28\] _06316_ vssd1 vssd1
+ vccd1 vccd1 _06317_ sky130_fd_sc_hd__or2_1
XANTENNA__09958__A0 net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12414_ net1386 vssd1 vssd1 vccd1 vccd1 _00178_ sky130_fd_sc_hd__inv_2
XANTENNA__08505__D _04444_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13394_ net1431 vssd1 vssd1 vccd1 vccd1 _01158_ sky130_fd_sc_hd__inv_2
XFILLER_0_35_395 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11765__B1 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12345_ net1355 vssd1 vssd1 vccd1 vccd1 _00109_ sky130_fd_sc_hd__inv_2
XFILLER_0_50_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15064_ net1450 vssd1 vssd1 vccd1 vccd1 la_data_out[0] sky130_fd_sc_hd__buf_2
XFILLER_0_26_1039 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12276_ net1308 vssd1 vssd1 vccd1 vccd1 _00040_ sky130_fd_sc_hd__inv_2
X_14015_ clknet_leaf_169_wb_clk_i _01779_ _00380_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[369\]
+ sky130_fd_sc_hd__dfrtp_1
X_11227_ _06527_ net2238 net488 vssd1 vssd1 vccd1 vccd1 _02184_ sky130_fd_sc_hd__mux2_1
XANTENNA__10125__A _04532_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08394__C1 net1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09914__A _05659_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_156_wb_clk_i clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_156_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_11158_ net513 net656 _06656_ net415 net1931 vssd1 vssd1 vccd1 vccd1 _02226_ sky130_fd_sc_hd__a32o_1
XANTENNA__10740__A1 _05676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_147_3388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_147_3399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11655__S net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10109_ _04770_ net676 _05949_ _03060_ vssd1 vssd1 vccd1 vccd1 _05953_ sky130_fd_sc_hd__o211ai_2
X_11089_ _06621_ net2628 net416 vssd1 vssd1 vccd1 vccd1 _02260_ sky130_fd_sc_hd__mux2_1
XANTENNA__08146__C1 net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07434__A net1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14917_ clknet_leaf_50_wb_clk_i _02672_ _01282_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_O\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_125_2941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_125_2952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11296__A2 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_159_Right_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14848_ clknet_leaf_83_wb_clk_i _02612_ _01213_ vssd1 vssd1 vccd1 vccd1 net134 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_19_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11048__A2 net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14779_ clknet_leaf_100_wb_clk_i _02543_ _01144_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_I\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_07320_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[29\] net768
+ net743 _03261_ vssd1 vssd1 vccd1 vccd1 _03262_ sky130_fd_sc_hd__a211o_1
XANTENNA__13171__A net1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_173_3927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07251_ _03190_ _03192_ net815 vssd1 vssd1 vccd1 vccd1 _03193_ sky130_fd_sc_hd__a21o_1
XANTENNA__07672__A1 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10008__A0 _02921_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07182_ net1175 team_03_WB.instance_to_wrap.core.register_file.registers_state\[723\]
+ net762 team_03_WB.instance_to_wrap.core.register_file.registers_state\[755\] net741
+ vssd1 vssd1 vccd1 vccd1 _03124_ sky130_fd_sc_hd__o221a_1
XFILLER_0_14_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11122__C net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_15_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11756__B1 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_490 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_30_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07424__A1 net1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10734__S _06295_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11771__A3 net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout404 _06717_ vssd1 vssd1 vccd1 vccd1 net404 sky130_fd_sc_hd__buf_8
Xfanout415 _06635_ vssd1 vssd1 vccd1 vccd1 net415 sky130_fd_sc_hd__clkbuf_4
Xfanout426 _04079_ vssd1 vssd1 vccd1 vccd1 net426 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08924__A1 net1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout437 net438 vssd1 vssd1 vccd1 vccd1 net437 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09824__A _05073_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09823_ _05265_ _05267_ vssd1 vssd1 vccd1 vccd1 _05765_ sky130_fd_sc_hd__xnor2_1
Xfanout448 _06801_ vssd1 vssd1 vccd1 vccd1 net448 sky130_fd_sc_hd__clkbuf_4
Xfanout459 net460 vssd1 vssd1 vccd1 vccd1 net459 sky130_fd_sc_hd__clkbuf_2
X_09754_ net351 _05569_ _05690_ _05691_ _05695_ vssd1 vssd1 vccd1 vccd1 _05696_ sky130_fd_sc_hd__a221o_1
X_06966_ net1113 team_03_WB.instance_to_wrap.core.register_file.registers_state\[965\]
+ net802 team_03_WB.instance_to_wrap.core.register_file.registers_state\[997\] net1137
+ vssd1 vssd1 vccd1 vccd1 _02908_ sky130_fd_sc_hd__a221o_1
XFILLER_0_20_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09035__S net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08705_ _04646_ vssd1 vssd1 vccd1 vccd1 _04647_ sky130_fd_sc_hd__inv_2
XFILLER_0_146_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09685_ net664 _05626_ _03988_ _04178_ vssd1 vssd1 vccd1 vccd1 _05627_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_69_708 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout554_A _03064_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06897_ _02815_ _02828_ _02832_ _02794_ vssd1 vssd1 vccd1 vccd1 _02839_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_154_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10495__B1 net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_169_Left_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_126_Right_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_1115 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08636_ net1065 _04576_ _04577_ vssd1 vssd1 vccd1 vccd1 _04578_ sky130_fd_sc_hd__a21o_1
XFILLER_0_68_218 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_538 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07360__B1 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_81_2034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11039__A2 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_2045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08567_ net1235 team_03_WB.instance_to_wrap.core.register_file.registers_state\[93\]
+ net966 team_03_WB.instance_to_wrap.core.register_file.registers_state\[125\] net922
+ vssd1 vssd1 vccd1 vccd1 _04509_ sky130_fd_sc_hd__o221a_1
XANTENNA__10909__S net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout721_A _02863_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout342_X net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_54_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout1084_X net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout819_A net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07518_ team_03_WB.instance_to_wrap.core.decoder.inst\[26\] net826 vssd1 vssd1 vccd1
+ vccd1 _03460_ sky130_fd_sc_hd__and2_2
XFILLER_0_92_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10798__A1 net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08498_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[443\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[411\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[315\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[283\]
+ net987 net1079 vssd1 vssd1 vccd1 vccd1 _04440_ sky130_fd_sc_hd__mux4_1
XANTENNA__07112__B1 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_153_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09652__A2 _05545_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11995__B1 net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07663__A1 net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07449_ _03389_ _03390_ net610 vssd1 vssd1 vccd1 vccd1 _03391_ sky130_fd_sc_hd__mux2_4
XFILLER_0_134_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout607_X net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08860__B1 net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_788 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10460_ net304 _05945_ _06043_ _06050_ vssd1 vssd1 vccd1 vccd1 _06274_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_134_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08903__A net1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11747__B1 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09119_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[686\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[654\]
+ net976 vssd1 vssd1 vccd1 vccd1 _05061_ sky130_fd_sc_hd__mux2_1
XANTENNA__07415__A1 net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10391_ net284 _06144_ _06215_ net680 vssd1 vssd1 vccd1 vccd1 _06219_ sky130_fd_sc_hd__o31a_1
XANTENNA__10644__S net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08612__B1 net992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_1__f_wb_clk_i_X clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_12130_ net1549 vssd1 vssd1 vccd1 vccd1 _02423_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_130_551 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout976_X net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12061_ _06505_ net2615 net357 vssd1 vssd1 vccd1 vccd1 _01485_ sky130_fd_sc_hd__mux2_1
Xhold480 team_03_WB.instance_to_wrap.core.ru.state\[3\] vssd1 vssd1 vccd1 vccd1 net1973
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_129_3030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold491 team_03_WB.instance_to_wrap.core.register_file.registers_state\[443\] vssd1
+ vssd1 vccd1 vccd1 net1984 sky130_fd_sc_hd__dlygate4sd3_1
X_11012_ net500 net652 _06579_ net421 net1919 vssd1 vssd1 vccd1 vccd1 _02295_ sky130_fd_sc_hd__a32o_1
XFILLER_0_25_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_53_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout960 net962 vssd1 vssd1 vccd1 vccd1 net960 sky130_fd_sc_hd__clkbuf_4
Xfanout971 net973 vssd1 vssd1 vccd1 vccd1 net971 sky130_fd_sc_hd__clkbuf_2
Xfanout982 net983 vssd1 vssd1 vccd1 vccd1 net982 sky130_fd_sc_hd__clkbuf_4
Xfanout993 net994 vssd1 vssd1 vccd1 vccd1 net993 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_5_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_93_wb_clk_i_A clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__07254__A net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12963_ net1374 vssd1 vssd1 vccd1 vccd1 _00727_ sky130_fd_sc_hd__inv_2
XANTENNA__11278__A2 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_142_3285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1180 team_03_WB.instance_to_wrap.core.register_file.registers_state\[870\] vssd1
+ vssd1 vccd1 vccd1 net2673 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_87_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14702_ clknet_leaf_56_wb_clk_i _02466_ _01067_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.SEL_I\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1191 team_03_WB.instance_to_wrap.core.register_file.registers_state\[128\] vssd1
+ vssd1 vccd1 vccd1 net2684 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10486__B1 net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_142_3296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11914_ _06615_ net2744 net368 vssd1 vssd1 vccd1 vccd1 _01628_ sky130_fd_sc_hd__mux2_1
XFILLER_0_158_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12894_ net1409 vssd1 vssd1 vccd1 vccd1 _00658_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_16_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14633_ clknet_leaf_78_wb_clk_i _02397_ _00998_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[987\]
+ sky130_fd_sc_hd__dfstp_1
X_11845_ _06413_ net2018 net376 vssd1 vssd1 vccd1 vccd1 _01695_ sky130_fd_sc_hd__mux2_1
XFILLER_0_169_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_796 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14564_ clknet_leaf_15_wb_clk_i _02328_ _00929_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[918\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_83_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11776_ net1042 _06462_ net382 vssd1 vssd1 vccd1 vccd1 _06810_ sky130_fd_sc_hd__and3_4
XFILLER_0_126_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11986__A0 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08300__C1 net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13515_ net1307 vssd1 vssd1 vccd1 vccd1 _01279_ sky130_fd_sc_hd__inv_2
XFILLER_0_82_232 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10727_ net1742 net527 net522 _06355_ vssd1 vssd1 vccd1 vccd1 _02452_ sky130_fd_sc_hd__a22o_1
XFILLER_0_126_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14495_ clknet_leaf_167_wb_clk_i _02259_ _00860_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[849\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08851__B1 net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_479 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13446_ net1406 vssd1 vssd1 vccd1 vccd1 _01210_ sky130_fd_sc_hd__inv_2
XFILLER_0_125_356 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10658_ team_03_WB.instance_to_wrap.core.control_logic.instruction\[3\] team_03_WB.instance_to_wrap.CPU_DAT_O\[3\]
+ net846 vssd1 vssd1 vccd1 vccd1 _02470_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload14 clknet_leaf_189_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload14/Y sky130_fd_sc_hd__clkinv_4
XANTENNA__11738__B1 _06808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07406__A1 net1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload25 clknet_leaf_16_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload25/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_24_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkload36 clknet_leaf_182_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload36/Y sky130_fd_sc_hd__inv_6
X_13377_ net1431 vssd1 vssd1 vccd1 vccd1 _01141_ sky130_fd_sc_hd__inv_2
Xclkload47 clknet_leaf_167_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload47/Y sky130_fd_sc_hd__clkinv_4
X_10589_ net1142 team_03_WB.instance_to_wrap.WRITE_I net1145 _06292_ vssd1 vssd1 vccd1
+ vccd1 _02534_ sky130_fd_sc_hd__a22o_1
XFILLER_0_11_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload58 clknet_leaf_37_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload58/Y sky130_fd_sc_hd__clkinv_1
Xclkload69 clknet_leaf_49_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload69/Y sky130_fd_sc_hd__clkinvlp_4
XTAP_TAPCELL_ROW_77_1958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15116_ net912 vssd1 vssd1 vccd1 vccd1 net249 sky130_fd_sc_hd__clkbuf_1
X_12328_ net1290 vssd1 vssd1 vccd1 vccd1 _00092_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_149_3428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_149_3439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09159__A1 net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15047_ net171 vssd1 vssd1 vccd1 vccd1 net170 sky130_fd_sc_hd__clkbuf_1
X_12259_ net1372 vssd1 vssd1 vccd1 vccd1 _00023_ sky130_fd_sc_hd__inv_2
XANTENNA__08906__A1 net1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_166_3775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_166_3786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06917__B1 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13166__A net1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08119__C1 net1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10477__B1 net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09470_ net569 _05407_ _05411_ net321 vssd1 vssd1 vccd1 vccd1 _05412_ sky130_fd_sc_hd__o211a_1
XFILLER_0_78_538 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07342__B1 net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08421_ net1228 team_03_WB.instance_to_wrap.core.register_file.registers_state\[346\]
+ net954 team_03_WB.instance_to_wrap.core.register_file.registers_state\[378\] net1072
+ vssd1 vssd1 vccd1 vccd1 _04363_ sky130_fd_sc_hd__o221a_1
XANTENNA__14993__Q team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[12\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_83 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07893__A1 net1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_53_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_53_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_08352_ _04280_ _04293_ net849 vssd1 vssd1 vccd1 vccd1 _04294_ sky130_fd_sc_hd__mux2_4
XFILLER_0_50_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11977__A0 _06413_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07303_ net1185 team_03_WB.instance_to_wrap.core.register_file.registers_state\[701\]
+ net879 vssd1 vssd1 vccd1 vccd1 _03245_ sky130_fd_sc_hd__and3_1
XANTENNA__07645__A1 net1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11441__A2 net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08842__B1 net1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08283_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[759\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[727\]
+ net963 vssd1 vssd1 vccd1 vccd1 _04225_ sky130_fd_sc_hd__mux2_1
XFILLER_0_144_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_138_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xclkload8 clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload8/Y sky130_fd_sc_hd__clkinv_2
XFILLER_0_74_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07234_ net1096 team_03_WB.instance_to_wrap.core.register_file.registers_state\[680\]
+ net896 vssd1 vssd1 vccd1 vccd1 _03176_ sky130_fd_sc_hd__or3_1
XFILLER_0_116_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08723__A net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07165_ _02808_ net1016 team_03_WB.instance_to_wrap.core.decoder.inst\[31\] vssd1
+ vssd1 vccd1 vccd1 _03107_ sky130_fd_sc_hd__o21a_4
XFILLER_0_131_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout302_A _06422_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08442__B net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08070__A1 net1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07096_ net1196 team_03_WB.instance_to_wrap.core.register_file.registers_state\[865\]
+ net884 _03037_ net1155 vssd1 vssd1 vccd1 vccd1 _03038_ sky130_fd_sc_hd__a311o_1
XFILLER_0_30_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1211_A net1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1309_A net1330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08358__C1 net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09554__A net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout671_A _06563_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout292_X net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11901__B1 net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout769_A net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09570__A1 net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09806_ _05268_ _05747_ vssd1 vssd1 vccd1 vccd1 _05748_ sky130_fd_sc_hd__nor2_1
XANTENNA__07030__C1 net1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout267 _06550_ vssd1 vssd1 vccd1 vccd1 net267 sky130_fd_sc_hd__buf_2
XFILLER_0_157_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout278 _06426_ vssd1 vssd1 vccd1 vccd1 net278 sky130_fd_sc_hd__buf_2
Xfanout289 net290 vssd1 vssd1 vccd1 vccd1 net289 sky130_fd_sc_hd__clkbuf_4
X_07998_ _03935_ _03936_ net814 vssd1 vssd1 vccd1 vccd1 _03940_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07581__B1 net1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09737_ _03790_ _04953_ vssd1 vssd1 vccd1 vccd1 _05679_ sky130_fd_sc_hd__or2_1
X_06949_ net612 _02888_ _02890_ vssd1 vssd1 vccd1 vccd1 _02891_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_2_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout936_A net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09668_ net321 _05533_ _05603_ net352 _05608_ vssd1 vssd1 vccd1 vccd1 _05610_ sky130_fd_sc_hd__a221oi_4
XANTENNA__11027__C net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_177_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_16_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08619_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[421\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[389\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[293\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[261\]
+ net992 net1078 vssd1 vssd1 vccd1 vccd1 _04561_ sky130_fd_sc_hd__mux4_1
XANTENNA__10639__S net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09599_ net594 _05519_ _05540_ vssd1 vssd1 vccd1 vccd1 _05541_ sky130_fd_sc_hd__o21a_2
XANTENNA_fanout724_X net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11680__A2 net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_155_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11630_ _06704_ net384 net348 net2290 vssd1 vssd1 vccd1 vccd1 _01902_ sky130_fd_sc_hd__a22o_1
XFILLER_0_37_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09086__B1 net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_166_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11968__B1 net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11043__B _06517_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07097__C1 net1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_370 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_917 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11432__A2 net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11561_ net657 _06671_ vssd1 vssd1 vccd1 vccd1 _06795_ sky130_fd_sc_hd__nor2_1
XFILLER_0_135_632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13300_ net1327 vssd1 vssd1 vccd1 vccd1 _01064_ sky130_fd_sc_hd__inv_2
XANTENNA__10640__A0 net1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10512_ net1967 net1031 net1024 net1925 vssd1 vssd1 vccd1 vccd1 _02598_ sky130_fd_sc_hd__a22o_1
XFILLER_0_107_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_682 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14280_ clknet_leaf_9_wb_clk_i _02044_ _00645_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[634\]
+ sky130_fd_sc_hd__dfrtp_1
X_11492_ _06613_ net2728 net388 vssd1 vssd1 vccd1 vccd1 _02014_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_2383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_2394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13231_ net1339 vssd1 vssd1 vccd1 vccd1 _00995_ sky130_fd_sc_hd__inv_2
X_10443_ team_03_WB.instance_to_wrap.core.pc.current_pc\[6\] _06135_ team_03_WB.instance_to_wrap.core.pc.current_pc\[7\]
+ vssd1 vssd1 vccd1 vccd1 _06261_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_27_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08597__C1 net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_1097 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07249__A net1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input65_A gpio_in[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13162_ net1284 vssd1 vssd1 vccd1 vccd1 _00926_ sky130_fd_sc_hd__inv_2
XANTENNA__08061__A1 net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10374_ net282 _06204_ net677 vssd1 vssd1 vccd1 vccd1 _06205_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_27_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08071__C net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12113_ net1143 net1845 _06282_ team_03_WB.instance_to_wrap.core.ru.state\[5\] vssd1
+ vssd1 vccd1 vccd1 _00005_ sky130_fd_sc_hd__a22o_1
XFILLER_0_23_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13093_ net1348 vssd1 vssd1 vccd1 vccd1 _00857_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_72_1855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12044_ _06613_ net2692 net355 vssd1 vssd1 vccd1 vccd1 _01502_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_72_1866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_3325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_3336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_49 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout790 _02851_ vssd1 vssd1 vccd1 vccd1 net790 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_161_3672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13995_ clknet_leaf_40_wb_clk_i _01759_ _00360_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[349\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_161_3683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10459__A0 team_03_WB.instance_to_wrap.core.pc.current_pc\[4\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11933__S net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12946_ net1338 vssd1 vssd1 vccd1 vccd1 _00710_ sky130_fd_sc_hd__inv_2
XANTENNA__07324__B1 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08521__C1 net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_37 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_158_735 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12877_ net1293 vssd1 vssd1 vccd1 vccd1 _00641_ sky130_fd_sc_hd__inv_2
XFILLER_0_34_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14616_ clknet_leaf_3_wb_clk_i _02380_ _00981_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[970\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_157_256 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09077__B1 net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11828_ _06661_ net469 net325 net2077 vssd1 vssd1 vccd1 vccd1 _01711_ sky130_fd_sc_hd__a22o_1
XFILLER_0_55_210 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_530 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11959__B1 net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14547_ clknet_leaf_100_wb_clk_i _02311_ _00912_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[901\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08824__B1 net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11759_ net657 _06585_ net477 net334 net2164 vssd1 vssd1 vccd1 vccd1 _01778_ sky130_fd_sc_hd__a32o_1
XANTENNA__10631__A0 team_03_WB.instance_to_wrap.core.decoder.inst\[30\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11521__X _06779_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14478_ clknet_leaf_130_wb_clk_i _02242_ _00843_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[832\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10792__B net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload103 clknet_leaf_150_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload103/Y sky130_fd_sc_hd__inv_4
XTAP_TAPCELL_ROW_116_2748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload114 clknet_leaf_122_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload114/Y sky130_fd_sc_hd__inv_8
X_13429_ net1428 vssd1 vssd1 vccd1 vccd1 _01193_ sky130_fd_sc_hd__inv_2
XFILLER_0_113_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkload125 clknet_leaf_138_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload125/Y sky130_fd_sc_hd__bufinv_16
XTAP_TAPCELL_ROW_116_2759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload136 clknet_leaf_131_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload136/Y sky130_fd_sc_hd__clkinvlp_4
XANTENNA__11187__A1 net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload147 clknet_leaf_112_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload147/Y sky130_fd_sc_hd__bufinv_16
Xclkload158 clknet_leaf_101_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload158/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_3_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_168_3815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload169 clknet_leaf_130_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload169/Y sky130_fd_sc_hd__inv_6
XTAP_TAPCELL_ROW_168_3826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_171_wb_clk_i clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_171_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_11_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_100_wb_clk_i clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_100_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_08970_ net1059 team_03_WB.instance_to_wrap.core.register_file.registers_state\[649\]
+ net1013 team_03_WB.instance_to_wrap.core.register_file.registers_state\[681\] net929
+ vssd1 vssd1 vccd1 vccd1 _04912_ sky130_fd_sc_hd__a221o_1
XFILLER_0_11_379 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10016__C net69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14988__Q team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[7\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07921_ net1138 _03852_ _03862_ vssd1 vssd1 vccd1 vccd1 _03863_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10698__B1 net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07852_ net1200 team_03_WB.instance_to_wrap.core.register_file.registers_state\[603\]
+ net784 team_03_WB.instance_to_wrap.core.register_file.registers_state\[635\] net737
+ vssd1 vssd1 vccd1 vccd1 _03794_ sky130_fd_sc_hd__o221a_1
Xinput1 ACK_I vssd1 vssd1 vccd1 vccd1 net1 sky130_fd_sc_hd__buf_4
X_07783_ net616 _03724_ vssd1 vssd1 vccd1 vccd1 _03725_ sky130_fd_sc_hd__nor2_1
XFILLER_0_36_60 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11843__S net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09522_ _05351_ _05373_ net562 vssd1 vssd1 vccd1 vccd1 _05464_ sky130_fd_sc_hd__mux2_1
XANTENNA__06937__S net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07315__B1 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10967__B net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07622__A team_03_WB.instance_to_wrap.core.decoder.inst\[25\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09453_ _05109_ _05112_ vssd1 vssd1 vccd1 vccd1 _05395_ sky130_fd_sc_hd__nor2_1
XFILLER_0_78_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08404_ net947 _04345_ _04344_ net1068 vssd1 vssd1 vccd1 vccd1 _04346_ sky130_fd_sc_hd__o211a_1
XANTENNA__11144__A net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09384_ _03529_ _05157_ vssd1 vssd1 vccd1 vccd1 _05326_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_19_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08335_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[885\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[853\]
+ net968 vssd1 vssd1 vccd1 vccd1 _04277_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_1069 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08815__B1 net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11414__A2 net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1161_A net1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_574 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1259_A net1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08266_ net433 net427 _04207_ vssd1 vssd1 vccd1 vccd1 _04208_ sky130_fd_sc_hd__nor3_1
XFILLER_0_144_451 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11965__A3 net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08830__A3 _04770_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07217_ net1160 _03158_ _03155_ vssd1 vssd1 vccd1 vccd1 _03159_ sky130_fd_sc_hd__o21a_1
XFILLER_0_116_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08197_ net1045 team_03_WB.instance_to_wrap.core.register_file.registers_state\[659\]
+ net995 team_03_WB.instance_to_wrap.core.register_file.registers_state\[691\] net918
+ vssd1 vssd1 vccd1 vccd1 _04139_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout1426_A net1436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09983__S net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1047_X net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08043__A1 net1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07148_ net752 _03088_ net814 vssd1 vssd1 vccd1 vccd1 _03090_ sky130_fd_sc_hd__o21a_1
XFILLER_0_14_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout886_A net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_2280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_2291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07079_ _03016_ _03020_ _03019_ net1119 vssd1 vssd1 vccd1 vccd1 _03021_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA_fanout1214_X net1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_7_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09284__A _04922_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10090_ _05623_ _05632_ _05659_ vssd1 vssd1 vccd1 vccd1 _05934_ sky130_fd_sc_hd__nor3_1
Xfanout1007 net1008 vssd1 vssd1 vccd1 vccd1 net1007 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_100_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1018 _02809_ vssd1 vssd1 vccd1 vccd1 net1018 sky130_fd_sc_hd__clkbuf_4
Xfanout1029 net1035 vssd1 vssd1 vccd1 vccd1 net1029 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout674_X net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11350__A1 net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07554__B1 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11038__B net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout841_X net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout939_X net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12800_ net1402 vssd1 vssd1 vccd1 vccd1 _00564_ sky130_fd_sc_hd__inv_2
X_13780_ clknet_leaf_124_wb_clk_i _01544_ _00145_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[134\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07306__B1 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10992_ net627 _06567_ vssd1 vssd1 vccd1 vccd1 _06568_ sky130_fd_sc_hd__nor2_1
XANTENNA__07532__A net1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12731_ net1361 vssd1 vssd1 vccd1 vccd1 _00495_ sky130_fd_sc_hd__inv_2
XANTENNA__07857__A1 net1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12662_ net1262 vssd1 vssd1 vccd1 vccd1 _00426_ sky130_fd_sc_hd__inv_2
XFILLER_0_32_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09059__B1 net1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14401_ clknet_leaf_180_wb_clk_i _02165_ _00766_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[755\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08066__C net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11613_ _06687_ net381 net346 net1968 vssd1 vssd1 vccd1 vccd1 _01919_ sky130_fd_sc_hd__a22o_1
XANTENNA__08806__B1 net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12593_ net1266 vssd1 vssd1 vccd1 vccd1 _00357_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_137_3184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14332_ clknet_leaf_157_wb_clk_i _02096_ _00697_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[686\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_3195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07085__A2 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11956__A3 net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11544_ net651 _06654_ vssd1 vssd1 vccd1 vccd1 _06788_ sky130_fd_sc_hd__nor2_1
XFILLER_0_53_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_150_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07490__C1 net1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14263_ clknet_leaf_115_wb_clk_i _02027_ _00628_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[617\]
+ sky130_fd_sc_hd__dfrtp_1
X_11475_ net657 _06600_ vssd1 vssd1 vccd1 vccd1 _06773_ sky130_fd_sc_hd__nor2_1
XFILLER_0_34_983 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11169__B2 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13214_ net1413 vssd1 vssd1 vccd1 vccd1 _00978_ sky130_fd_sc_hd__inv_2
X_10426_ _06021_ _06062_ _06017_ vssd1 vssd1 vccd1 vccd1 _06247_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_122_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08034__A1 net1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_1906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14194_ clknet_leaf_163_wb_clk_i _01958_ _00559_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[548\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10916__A1 net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09782__A1 net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11928__S net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13145_ net1359 vssd1 vssd1 vccd1 vccd1 _00909_ sky130_fd_sc_hd__inv_2
X_10357_ net283 _06190_ vssd1 vssd1 vccd1 vccd1 _06191_ sky130_fd_sc_hd__nand2_1
XANTENNA__09906__B _05833_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10832__S net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_2656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07793__B1 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08990__C1 net1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07707__A net1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_163_3712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13076_ net1313 vssd1 vssd1 vccd1 vccd1 _00840_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_163_3723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10288_ _05363_ _06129_ vssd1 vssd1 vccd1 vccd1 _06130_ sky130_fd_sc_hd__xnor2_1
X_12027_ _06769_ net468 net361 net2326 vssd1 vssd1 vccd1 vccd1 _01518_ sky130_fd_sc_hd__a22o_1
XANTENNA__07545__B1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07640__S0 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11663__S net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13978_ clknet_leaf_145_wb_clk_i _01742_ _00343_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[332\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10787__B net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_666 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07848__A1 _03789_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12929_ net1272 vssd1 vssd1 vccd1 vccd1 _00693_ sky130_fd_sc_hd__inv_2
XFILLER_0_38_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_124_Left_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_390 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_31 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_930 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_928 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08120_ _04059_ _04061_ net1160 vssd1 vssd1 vccd1 vccd1 _04062_ sky130_fd_sc_hd__o21a_1
XFILLER_0_142_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11947__A3 net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08273__A1 net1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08051_ net1186 team_03_WB.instance_to_wrap.core.register_file.registers_state\[182\]
+ vssd1 vssd1 vccd1 vccd1 _03993_ sky130_fd_sc_hd__and2_1
XFILLER_0_43_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07002_ net608 _02940_ _02943_ vssd1 vssd1 vccd1 vccd1 _02944_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_4_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08025__A1 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10742__S net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08953_ _04863_ _04894_ net550 vssd1 vssd1 vccd1 vccd1 _04895_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07904_ net1090 team_03_WB.instance_to_wrap.core.register_file.registers_state\[719\]
+ net794 team_03_WB.instance_to_wrap.core.register_file.registers_state\[751\] net729
+ vssd1 vssd1 vccd1 vccd1 _03846_ sky130_fd_sc_hd__a221o_1
XANTENNA__07336__B net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08884_ net544 _04825_ _04772_ vssd1 vssd1 vccd1 vccd1 _04826_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_138_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07536__B1 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1007_A net1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08733__C1 net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07835_ net1082 team_03_WB.instance_to_wrap.core.register_file.registers_state\[842\]
+ net791 team_03_WB.instance_to_wrap.core.register_file.registers_state\[874\] net1149
+ vssd1 vssd1 vccd1 vccd1 _03777_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout467_A net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_168_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07766_ net1098 team_03_WB.instance_to_wrap.core.register_file.registers_state\[620\]
+ net897 vssd1 vssd1 vccd1 vccd1 _03708_ sky130_fd_sc_hd__or3_1
XFILLER_0_155_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11096__A0 _06624_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09505_ _04416_ _04446_ _04505_ _04533_ net547 net559 vssd1 vssd1 vccd1 vccd1 _05447_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__07352__A net1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11635__A2 net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_603 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07697_ team_03_WB.instance_to_wrap.core.decoder.inst\[30\] net1020 vssd1 vssd1 vccd1
+ vccd1 _03639_ sky130_fd_sc_hd__nand2_1
XFILLER_0_52_1024 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout634_A net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1376_A net1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09436_ _05374_ _05377_ net567 vssd1 vssd1 vccd1 vccd1 _05378_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09978__S net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07814__A1_N net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09367_ _05183_ _05190_ _05308_ vssd1 vssd1 vccd1 vccd1 _05309_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_23_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout801_A net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout422_X net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11024__D net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1164_X net1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07498__S net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09279__A _04893_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08318_ net1073 _04258_ _04259_ net875 vssd1 vssd1 vccd1 vccd1 _04260_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_43_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08264__A1 net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_298 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_224 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09298_ _05239_ vssd1 vssd1 vccd1 vccd1 _05240_ sky130_fd_sc_hd__inv_2
XFILLER_0_105_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_95_2320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_566 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_2331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07472__C1 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08249_ net1062 _04188_ _04189_ vssd1 vssd1 vccd1 vccd1 _04191_ sky130_fd_sc_hd__or3_1
XFILLER_0_104_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10218__A _06057_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11260_ net494 net623 _06697_ net408 net2297 vssd1 vssd1 vccd1 vccd1 _02165_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_132_3081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout791_X net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_3092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_91_2239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout889_X net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10211_ _06051_ _06052_ _06040_ vssd1 vssd1 vccd1 vccd1 _06053_ sky130_fd_sc_hd__a21o_1
XANTENNA__09764__A1 net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10652__S net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11191_ net2313 net414 _06676_ net507 vssd1 vssd1 vccd1 vccd1 _02213_ sky130_fd_sc_hd__a22o_1
X_15109__1484 vssd1 vssd1 vccd1 vccd1 _15109__1484/HI net1484 sky130_fd_sc_hd__conb_1
XFILLER_0_31_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08972__C1 net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11571__B2 net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10142_ team_03_WB.instance_to_wrap.core.pc.current_pc\[19\] net672 vssd1 vssd1 vccd1
+ vccd1 _05984_ sky130_fd_sc_hd__nand2_1
Xoutput190 net190 vssd1 vssd1 vccd1 vccd1 gpio_oeb[25] sky130_fd_sc_hd__buf_2
XANTENNA__11049__A net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10073_ _02814_ _05916_ vssd1 vssd1 vccd1 vccd1 _05917_ sky130_fd_sc_hd__or2_1
X_14950_ clknet_leaf_101_wb_clk_i _02702_ _01315_ vssd1 vssd1 vccd1 vccd1 net233 sky130_fd_sc_hd__dfrtp_1
XANTENNA__07814__X _03756_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13901_ clknet_leaf_188_wb_clk_i _01665_ _00266_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[255\]
+ sky130_fd_sc_hd__dfrtp_1
X_14881_ clknet_leaf_82_wb_clk_i _02644_ _01246_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.pc.current_pc\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input28_A DAT_I[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13264__A net1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13832_ clknet_leaf_6_wb_clk_i _01596_ _00197_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[186\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09819__A2 _04679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13763_ clknet_leaf_34_wb_clk_i _01527_ _00128_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[117\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_67_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10975_ _02829_ net692 _06552_ _06553_ vssd1 vssd1 vccd1 vccd1 _06554_ sky130_fd_sc_hd__and4b_1
XFILLER_0_43_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11626__A2 net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09295__A3 _05144_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_139_3224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12714_ net1284 vssd1 vssd1 vccd1 vccd1 _00478_ sky130_fd_sc_hd__inv_2
XFILLER_0_84_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_139_3235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13694_ clknet_leaf_118_wb_clk_i _01458_ _00059_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[48\]
+ sky130_fd_sc_hd__dfrtp_1
X_12645_ net1355 vssd1 vssd1 vccd1 vccd1 _00409_ sky130_fd_sc_hd__inv_2
XFILLER_0_155_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10827__S net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_156_3571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_156_3582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08093__A net1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12576_ net1399 vssd1 vssd1 vccd1 vccd1 _00340_ sky130_fd_sc_hd__inv_2
XFILLER_0_80_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10062__A1 net13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14315_ clknet_leaf_46_wb_clk_i _02079_ _00680_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[669\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10062__B2 team_03_WB.instance_to_wrap.CPU_DAT_O\[1\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_11527_ net2236 net482 _06782_ net499 vssd1 vssd1 vccd1 vccd1 _01983_ sky130_fd_sc_hd__a22o_1
XFILLER_0_135_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_966 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09917__A _05082_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold309 team_03_WB.instance_to_wrap.core.register_file.registers_state\[316\] vssd1
+ vssd1 vccd1 vccd1 net1802 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08007__A1 net1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14246_ clknet_leaf_27_wb_clk_i _02010_ _00611_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[600\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_151_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11458_ net648 _06583_ vssd1 vssd1 vccd1 vccd1 _06766_ sky130_fd_sc_hd__nor2_1
XFILLER_0_151_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09755__A1 net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11658__S net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10409_ team_03_WB.instance_to_wrap.core.pc.current_pc\[13\] _06140_ vssd1 vssd1
+ vccd1 vccd1 _06233_ sky130_fd_sc_hd__nor2_1
XANTENNA__08102__S1 net1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14177_ clknet_leaf_183_wb_clk_i _01941_ _00542_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[531\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_3_4_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_4_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_68_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11389_ net712 net268 net697 vssd1 vssd1 vccd1 vccd1 _06747_ sky130_fd_sc_hd__and3_1
XFILLER_0_21_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11562__B2 net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13128_ net1296 vssd1 vssd1 vccd1 vccd1 _00892_ sky130_fd_sc_hd__inv_2
Xclkbuf_4_12__f_wb_clk_i clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_12__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
X_13059_ net1354 vssd1 vssd1 vccd1 vccd1 _00823_ sky130_fd_sc_hd__inv_2
XFILLER_0_139_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1009 team_03_WB.instance_to_wrap.core.register_file.registers_state\[157\] vssd1
+ vssd1 vccd1 vccd1 net2502 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_108_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1360 net1364 vssd1 vssd1 vccd1 vccd1 net1360 sky130_fd_sc_hd__buf_4
Xfanout1371 net1373 vssd1 vssd1 vccd1 vccd1 net1371 sky130_fd_sc_hd__buf_4
XFILLER_0_75_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1382 net1384 vssd1 vssd1 vccd1 vccd1 net1382 sky130_fd_sc_hd__buf_4
XFILLER_0_84_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1393 net1437 vssd1 vssd1 vccd1 vccd1 net1393 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_128_2994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07620_ net819 _03560_ _03561_ _03553_ _03556_ vssd1 vssd1 vccd1 vccd1 _03562_ sky130_fd_sc_hd__a32o_1
XFILLER_0_89_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_132_Left_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07551_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[24\] net783
+ net750 _03492_ vssd1 vssd1 vccd1 vccd1 _03493_ sky130_fd_sc_hd__a211o_1
XFILLER_0_159_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11617__A2 net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_496 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07482_ net1147 _03419_ _03421_ _03423_ net717 vssd1 vssd1 vccd1 vccd1 _03424_ sky130_fd_sc_hd__a41o_1
XFILLER_0_174_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09221_ _03641_ _05162_ vssd1 vssd1 vccd1 vccd1 _05163_ sky130_fd_sc_hd__xor2_1
XFILLER_0_146_535 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_173_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12518__A net1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire592_X net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09152_ net431 net425 _04444_ net541 vssd1 vssd1 vccd1 vccd1 _05094_ sky130_fd_sc_hd__o31a_1
XANTENNA__09443__A0 _05378_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08246__A1 net1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08103_ net1161 _04044_ vssd1 vssd1 vccd1 vccd1 _04045_ sky130_fd_sc_hd__or2_1
XFILLER_0_86_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10053__B2 team_03_WB.instance_to_wrap.CPU_DAT_O\[10\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11250__B1 net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09083_ net1069 _05022_ _05023_ vssd1 vssd1 vccd1 vccd1 _05025_ sky130_fd_sc_hd__or3_1
XPHY_EDGE_ROW_141_Left_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09181__A2_N _04807_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08034_ net1085 team_03_WB.instance_to_wrap.core.register_file.registers_state\[497\]
+ net890 _03975_ net1150 vssd1 vssd1 vccd1 vccd1 _03976_ sky130_fd_sc_hd__o311a_1
XANTENNA__09827__A _05768_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput70 wbs_adr_i[12] vssd1 vssd1 vccd1 vccd1 net70 sky130_fd_sc_hd__buf_1
XFILLER_0_31_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput81 wbs_adr_i[22] vssd1 vssd1 vccd1 vccd1 net81 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold810 team_03_WB.instance_to_wrap.core.register_file.registers_state\[778\] vssd1
+ vssd1 vccd1 vccd1 net2303 sky130_fd_sc_hd__dlygate4sd3_1
Xhold821 team_03_WB.instance_to_wrap.core.register_file.registers_state\[886\] vssd1
+ vssd1 vccd1 vccd1 net2314 sky130_fd_sc_hd__dlygate4sd3_1
Xhold832 team_03_WB.instance_to_wrap.core.register_file.registers_state\[550\] vssd1
+ vssd1 vccd1 vccd1 net2325 sky130_fd_sc_hd__dlygate4sd3_1
Xinput92 wbs_adr_i[3] vssd1 vssd1 vccd1 vccd1 net92 sky130_fd_sc_hd__clkbuf_1
XANTENNA__13349__A net1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07206__C1 net1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold843 team_03_WB.instance_to_wrap.core.register_file.registers_state\[360\] vssd1
+ vssd1 vccd1 vccd1 net2336 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold854 team_03_WB.instance_to_wrap.core.register_file.registers_state\[672\] vssd1
+ vssd1 vccd1 vccd1 net2347 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1124_A net1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold865 team_03_WB.instance_to_wrap.core.register_file.registers_state\[504\] vssd1
+ vssd1 vccd1 vccd1 net2358 sky130_fd_sc_hd__dlygate4sd3_1
Xhold876 team_03_WB.instance_to_wrap.core.register_file.registers_state\[760\] vssd1
+ vssd1 vccd1 vccd1 net2369 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11553__B2 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold887 team_03_WB.instance_to_wrap.core.register_file.registers_state\[784\] vssd1
+ vssd1 vccd1 vccd1 net2380 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09038__S net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold898 team_03_WB.instance_to_wrap.CPU_DAT_O\[28\] vssd1 vssd1 vccd1 vccd1 net2391
+ sky130_fd_sc_hd__dlygate4sd3_1
X_09985_ _05870_ net1885 net289 vssd1 vssd1 vccd1 vccd1 _02729_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08936_ net1046 team_03_WB.instance_to_wrap.core.register_file.registers_state\[971\]
+ net997 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1003\] net1061
+ vssd1 vssd1 vccd1 vccd1 _04878_ sky130_fd_sc_hd__a221o_1
XANTENNA__10108__A2 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07509__B1 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08867_ _02937_ net556 net544 vssd1 vssd1 vccd1 vccd1 _04809_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout372_X net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout751_A net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_150_Left_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11019__D net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout849_A _04097_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07818_ net1085 team_03_WB.instance_to_wrap.core.register_file.registers_state\[42\]
+ net890 vssd1 vssd1 vccd1 vccd1 _03760_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_88_2190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08798_ net434 net429 net592 net544 vssd1 vssd1 vccd1 vccd1 _04740_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_28_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_8_wb_clk_i clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_8_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_07749_ net748 _03689_ _03690_ net809 vssd1 vssd1 vccd1 vccd1 _03691_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_28_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout637_X net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10760_ _05784_ net604 vssd1 vssd1 vccd1 vccd1 _06374_ sky130_fd_sc_hd__nand2_1
XANTENNA__11035__C net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_811 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09419_ _04820_ _05341_ vssd1 vssd1 vccd1 vccd1 _05361_ sky130_fd_sc_hd__nand2_1
X_10691_ net606 _06318_ _06330_ vssd1 vssd1 vccd1 vccd1 _06331_ sky130_fd_sc_hd__and3_1
XANTENNA__10647__S net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout804_X net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08625__B net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_522 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12430_ net1274 vssd1 vssd1 vccd1 vccd1 _00194_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_134_3121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_134_3132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12033__A2 net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10044__A1 net12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11051__B net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_145_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08332__S1 net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12361_ net1253 vssd1 vssd1 vccd1 vccd1 _00125_ sky130_fd_sc_hd__inv_2
XFILLER_0_63_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_739 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14100_ clknet_leaf_132_wb_clk_i _01864_ _00465_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[454\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07996__B1 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11312_ _06469_ net2551 net404 vssd1 vssd1 vccd1 vccd1 _02133_ sky130_fd_sc_hd__mux2_1
X_15080_ net1466 vssd1 vssd1 vccd1 vccd1 la_data_out[16] sky130_fd_sc_hd__buf_2
XFILLER_0_133_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12292_ net1356 vssd1 vssd1 vccd1 vccd1 _00056_ sky130_fd_sc_hd__inv_2
XFILLER_0_160_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14031_ clknet_leaf_144_wb_clk_i _01795_ _00396_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[385\]
+ sky130_fd_sc_hd__dfrtp_1
X_11243_ net302 net714 net830 vssd1 vssd1 vccd1 vccd1 _06689_ sky130_fd_sc_hd__and3_1
XFILLER_0_28_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07257__A net1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11174_ net491 net647 _06666_ net412 net1895 vssd1 vssd1 vccd1 vccd1 _02220_ sky130_fd_sc_hd__a32o_1
X_10125_ _04532_ net672 vssd1 vssd1 vccd1 vccd1 _05967_ sky130_fd_sc_hd__or2_1
XANTENNA__06971__A1 net1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14933_ clknet_leaf_51_wb_clk_i _02688_ _01298_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_O\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_10056_ net31 net1036 net909 team_03_WB.instance_to_wrap.CPU_DAT_O\[7\] vssd1 vssd1
+ vccd1 vccd1 _02675_ sky130_fd_sc_hd__o22a_1
XANTENNA__09903__C _05429_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08173__B1 net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14864_ clknet_leaf_64_wb_clk_i _02628_ _01229_ vssd1 vssd1 vccd1 vccd1 net120 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_106_2544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07920__B1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13815_ clknet_leaf_112_wb_clk_i _01579_ _00180_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[169\]
+ sky130_fd_sc_hd__dfrtp_1
X_14795_ clknet_leaf_94_wb_clk_i _02559_ _01160_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_I\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_158_3611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_158_3622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10807__A0 _06413_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13746_ clknet_leaf_164_wb_clk_i _01510_ _00111_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[100\]
+ sky130_fd_sc_hd__dfrtp_1
X_10958_ net688 _05784_ vssd1 vssd1 vccd1 vccd1 _06540_ sky130_fd_sc_hd__nand2_1
XFILLER_0_70_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08816__A net1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09411__S net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11480__B1 net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13677_ clknet_leaf_181_wb_clk_i _01441_ _00042_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10889_ net272 net2364 net521 vssd1 vssd1 vccd1 vccd1 _02322_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_14_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12628_ net1305 vssd1 vssd1 vccd1 vccd1 _00392_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_14_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12024__A2 net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11232__A0 net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_171_3877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_171_3888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12559_ net1337 vssd1 vssd1 vccd1 vccd1 _00323_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_514 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10586__A2 net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11783__A1 _06616_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_171 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold106 team_03_WB.instance_to_wrap.ADR_I\[0\] vssd1 vssd1 vccd1 vccd1 net1599 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold117 team_03_WB.instance_to_wrap.core.register_file.registers_state\[24\] vssd1
+ vssd1 vccd1 vccd1 net1610 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_9_Right_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold128 net173 vssd1 vssd1 vccd1 vccd1 net1621 sky130_fd_sc_hd__dlygate4sd3_1
Xhold139 team_03_WB.instance_to_wrap.core.register_file.registers_state\[988\] vssd1
+ vssd1 vccd1 vccd1 net1632 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13169__A net1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14229_ clknet_leaf_105_wb_clk_i _01993_ _00594_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[583\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_78_wb_clk_i clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_78_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_145_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1050 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07739__B1 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08936__C1 net1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11535__B2 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout608 net609 vssd1 vssd1 vccd1 vccd1 net608 sky130_fd_sc_hd__buf_2
XFILLER_0_0_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08400__A1 net1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout619 net620 vssd1 vssd1 vccd1 vccd1 net619 sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_107_Right_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09653__Y _05595_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09770_ net584 _05710_ _05711_ net352 vssd1 vssd1 vccd1 vccd1 _05712_ sky130_fd_sc_hd__o22a_1
XANTENNA__07754__A3 net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06982_ _02807_ _02811_ vssd1 vssd1 vccd1 vccd1 _02924_ sky130_fd_sc_hd__nor2_1
XFILLER_0_77_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09382__A _04354_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08721_ _04657_ _04662_ net874 vssd1 vssd1 vccd1 vccd1 _04663_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11838__A2 net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1190 net1206 vssd1 vssd1 vccd1 vccd1 net1190 sky130_fd_sc_hd__clkbuf_4
X_08652_ _04566_ _04593_ net557 vssd1 vssd1 vccd1 vccd1 _04594_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07911__B1 net1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_1011 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07603_ net1167 _03543_ _03544_ vssd1 vssd1 vccd1 vccd1 _03545_ sky130_fd_sc_hd__o21ai_1
XANTENNA__11136__B net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08583_ net1207 _04521_ _04524_ vssd1 vssd1 vccd1 vccd1 _04525_ sky130_fd_sc_hd__or3_1
XANTENNA__11851__S net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_44_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_113_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07534_ _03473_ _03475_ net809 vssd1 vssd1 vccd1 vccd1 _03476_ sky130_fd_sc_hd__o21a_1
XFILLER_0_77_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_1028 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08467__A1 net1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08011__S0 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06945__S net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09664__B1 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10467__S net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07465_ _03405_ _03406_ net817 vssd1 vssd1 vccd1 vccd1 _03407_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_76_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout332_A _06809_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1074_A _02789_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_499 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09204_ net526 _03491_ _05144_ vssd1 vssd1 vccd1 vccd1 _05146_ sky130_fd_sc_hd__nand3_2
XANTENNA__11152__A net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12015__A2 net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07396_ _03336_ _03337_ net740 vssd1 vssd1 vccd1 vccd1 _03338_ sky130_fd_sc_hd__mux2_1
XFILLER_0_146_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11223__A0 _06513_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09135_ net584 _05076_ vssd1 vssd1 vccd1 vccd1 _05077_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10991__A net1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1241_A net1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10577__A2 net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1339_A net1346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09066_ net1219 _05006_ _05007_ vssd1 vssd1 vccd1 vccd1 _05008_ sky130_fd_sc_hd__and3_1
XFILLER_0_170_880 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_994 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_744 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout799_A net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08017_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[657\] net792
+ net745 _03958_ vssd1 vssd1 vccd1 vccd1 _03959_ sky130_fd_sc_hd__o211a_1
Xhold640 team_03_WB.instance_to_wrap.core.register_file.registers_state\[673\] vssd1
+ vssd1 vccd1 vccd1 net2133 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_766 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold651 team_03_WB.instance_to_wrap.core.register_file.registers_state\[224\] vssd1
+ vssd1 vccd1 vccd1 net2144 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09991__S net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1127_X net1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_794 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold662 team_03_WB.instance_to_wrap.core.register_file.registers_state\[433\] vssd1
+ vssd1 vccd1 vccd1 net2155 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_38_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08927__C1 net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold673 team_03_WB.instance_to_wrap.core.register_file.registers_state\[160\] vssd1
+ vssd1 vccd1 vccd1 net2166 sky130_fd_sc_hd__dlygate4sd3_1
Xhold684 team_03_WB.instance_to_wrap.core.register_file.registers_state\[450\] vssd1
+ vssd1 vccd1 vccd1 net2177 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold695 team_03_WB.instance_to_wrap.core.register_file.registers_state\[749\] vssd1
+ vssd1 vccd1 vccd1 net2188 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout966_A net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09968_ _05888_ net1693 net294 vssd1 vssd1 vccd1 vccd1 _02743_ sky130_fd_sc_hd__mux2_1
XANTENNA__12711__A net1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08919_ net848 _04847_ _04860_ vssd1 vssd1 vccd1 vccd1 _04861_ sky130_fd_sc_hd__a21oi_2
XANTENNA__07805__A net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_83_wb_clk_i_A clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09899_ net352 _05735_ _05839_ _05840_ vssd1 vssd1 vccd1 vccd1 _05841_ sky130_fd_sc_hd__a211oi_4
XANTENNA_fanout754_X net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11930_ _06627_ net2548 net367 vssd1 vssd1 vccd1 vccd1 _01612_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_86_2149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10231__A _03864_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11861_ net298 net2474 net377 vssd1 vssd1 vccd1 vccd1 _01679_ sky130_fd_sc_hd__mux2_1
XANTENNA__11046__B net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout921_X net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_64_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13600_ net1268 vssd1 vssd1 vccd1 vccd1 _01364_ sky130_fd_sc_hd__inv_2
XFILLER_0_39_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10812_ _06418_ net2529 net518 vssd1 vssd1 vccd1 vccd1 _02334_ sky130_fd_sc_hd__mux2_1
XFILLER_0_170_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_0_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08458__A1 net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14580_ clknet_leaf_133_wb_clk_i _02344_ _00945_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[934\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_0_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11792_ net2197 _06622_ net330 vssd1 vssd1 vccd1 vccd1 _01746_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_101_2441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13531_ net1316 vssd1 vssd1 vccd1 vccd1 _01295_ sky130_fd_sc_hd__inv_2
XANTENNA__07540__A net1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_2452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10743_ net1654 net529 net524 _06363_ vssd1 vssd1 vccd1 vccd1 _02444_ sky130_fd_sc_hd__a22o_1
XANTENNA__07666__C1 net1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07130__A1 net1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_354 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13462_ net1328 vssd1 vssd1 vccd1 vccd1 _01226_ sky130_fd_sc_hd__inv_2
X_10674_ team_03_WB.instance_to_wrap.core.pc.current_pc\[25\] team_03_WB.instance_to_wrap.core.pc.current_pc\[24\]
+ team_03_WB.instance_to_wrap.core.pc.current_pc\[27\] team_03_WB.instance_to_wrap.core.pc.current_pc\[26\]
+ vssd1 vssd1 vccd1 vccd1 _06316_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_11_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input95_A wbs_adr_i[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_11_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_184 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12413_ net1383 vssd1 vssd1 vccd1 vccd1 _00177_ sky130_fd_sc_hd__inv_2
XANTENNA__07418__C1 net1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13393_ net1428 vssd1 vssd1 vccd1 vccd1 _01157_ sky130_fd_sc_hd__inv_2
XFILLER_0_106_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10568__A2 net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_508 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11765__A1 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1023 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12344_ net1379 vssd1 vssd1 vccd1 vccd1 _00108_ sky130_fd_sc_hd__inv_2
XFILLER_0_161_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07433__A2 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08630__A1 net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15063_ net1449 vssd1 vssd1 vccd1 vccd1 irq[2] sky130_fd_sc_hd__buf_2
XFILLER_0_50_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12275_ net1256 vssd1 vssd1 vccd1 vccd1 _00039_ sky130_fd_sc_hd__inv_2
XFILLER_0_65_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08918__C1 net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14014_ clknet_leaf_120_wb_clk_i _01778_ _00379_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[368\]
+ sky130_fd_sc_hd__dfrtp_1
X_11226_ net295 net2124 net489 vssd1 vssd1 vccd1 vccd1 _02185_ sky130_fd_sc_hd__mux2_1
XANTENNA__11936__S net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08394__B1 net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11157_ net707 net272 net699 vssd1 vssd1 vccd1 vccd1 _06656_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_147_3389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10108_ _04770_ net660 _05951_ _03060_ vssd1 vssd1 vccd1 vccd1 _05952_ sky130_fd_sc_hd__a211o_1
XANTENNA__07715__A net1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11088_ net832 net273 vssd1 vssd1 vccd1 vccd1 _06621_ sky130_fd_sc_hd__and2_2
XANTENNA__11237__A net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10039_ net18 net1040 _05906_ team_03_WB.instance_to_wrap.CPU_DAT_O\[24\] vssd1 vssd1
+ vccd1 vccd1 _02692_ sky130_fd_sc_hd__a22o_1
X_14916_ clknet_leaf_43_wb_clk_i _02671_ _01281_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_O\[3\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_125_2942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08697__A1 net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09894__B1 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14847_ clknet_leaf_83_wb_clk_i net1613 _01212_ vssd1 vssd1 vccd1 vccd1 net133 sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_125_wb_clk_i clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_125_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_19_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11671__S net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08449__A1 net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14778_ clknet_leaf_96_wb_clk_i _02542_ _01143_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_I\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_105_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_173_3917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_173_3928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10287__S net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13729_ clknet_leaf_179_wb_clk_i _01493_ _00094_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[83\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_129_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_156_663 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07250_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[136\] net774
+ net730 _03191_ vssd1 vssd1 vccd1 vccd1 _03192_ sky130_fd_sc_hd__a211o_1
XANTENNA_clkbuf_leaf_128_wb_clk_i_A clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_144_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_110 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11205__A0 _06430_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07181_ net1175 team_03_WB.instance_to_wrap.core.register_file.registers_state\[595\]
+ net762 team_03_WB.instance_to_wrap.core.register_file.registers_state\[627\] net726
+ vssd1 vssd1 vccd1 vccd1 _03123_ sky130_fd_sc_hd__o221a_1
XFILLER_0_82_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_171_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11122__D net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10559__A2 net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11756__A1 net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_30_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07449__X _03391_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08621__A1 net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_777 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08909__C1 net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout405 _06717_ vssd1 vssd1 vccd1 vccd1 net405 sky130_fd_sc_hd__buf_4
Xfanout416 _06610_ vssd1 vssd1 vccd1 vccd1 net416 sky130_fd_sc_hd__buf_8
XFILLER_0_39_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout427 _04079_ vssd1 vssd1 vccd1 vccd1 net427 sky130_fd_sc_hd__buf_2
X_09822_ _04777_ _05762_ _05763_ _05761_ vssd1 vssd1 vccd1 vccd1 _05764_ sky130_fd_sc_hd__a31o_1
XANTENNA__11846__S net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout438 _04075_ vssd1 vssd1 vccd1 vccd1 net438 sky130_fd_sc_hd__clkbuf_2
Xfanout449 _06801_ vssd1 vssd1 vccd1 vccd1 net449 sky130_fd_sc_hd__clkbuf_8
XANTENNA__10731__A2 net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09753_ net1020 _03724_ _04820_ _05692_ _05694_ vssd1 vssd1 vccd1 vccd1 _05695_ sky130_fd_sc_hd__a221o_1
X_06965_ net1113 team_03_WB.instance_to_wrap.core.register_file.registers_state\[837\]
+ net802 team_03_WB.instance_to_wrap.core.register_file.registers_state\[869\] net1159
+ vssd1 vssd1 vccd1 vccd1 _02907_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout282_A net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08704_ _04632_ _04645_ net849 vssd1 vssd1 vccd1 vccd1 _04646_ sky130_fd_sc_hd__mux2_8
X_09684_ _03988_ _04178_ _04816_ vssd1 vssd1 vccd1 vccd1 _05626_ sky130_fd_sc_hd__a21o_1
XANTENNA__08232__S0 net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06896_ _02794_ _02815_ vssd1 vssd1 vccd1 vccd1 _02838_ sky130_fd_sc_hd__nor2_1
XANTENNA_clkbuf_leaf_0_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_08635_ net1224 _04574_ _04575_ vssd1 vssd1 vccd1 vccd1 _04577_ sky130_fd_sc_hd__and3_1
XANTENNA_clkbuf_leaf_167_wb_clk_i_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11692__B1 net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10986__A _06463_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1191_A net1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07360__A1 net1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11581__S net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1289_A net1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_2035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08566_ net938 _04506_ _04507_ vssd1 vssd1 vccd1 vccd1 _04508_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_81_2046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07517_ _03430_ _03458_ net615 vssd1 vssd1 vccd1 vccd1 _03459_ sky130_fd_sc_hd__mux2_4
XFILLER_0_37_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08497_ net1243 team_03_WB.instance_to_wrap.core.register_file.registers_state\[475\]
+ net987 team_03_WB.instance_to_wrap.core.register_file.registers_state\[507\] net1216
+ vssd1 vssd1 vccd1 vccd1 _04439_ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout714_A net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout335_X net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10798__A2 net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1077_X net1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09986__S net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07448_ net1190 net1019 net684 vssd1 vssd1 vccd1 vccd1 _03390_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_135_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07663__A2 net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout502_X net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07379_ net1082 team_03_WB.instance_to_wrap.core.register_file.registers_state\[255\]
+ net888 vssd1 vssd1 vccd1 vccd1 _03321_ sky130_fd_sc_hd__or3_1
XANTENNA_fanout1244_X net1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11747__A1 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09118_ net1066 _05056_ _05059_ vssd1 vssd1 vccd1 vccd1 _05060_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08073__C1 net1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10390_ net304 net303 _06216_ _06217_ vssd1 vssd1 vccd1 vccd1 _06218_ sky130_fd_sc_hd__a211o_1
XANTENNA__08612__A1 net1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07415__A2 net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09049_ net1047 team_03_WB.instance_to_wrap.core.register_file.registers_state\[207\]
+ net998 team_03_WB.instance_to_wrap.core.register_file.registers_state\[239\] net921
+ vssd1 vssd1 vccd1 vccd1 _04991_ sky130_fd_sc_hd__a221o_1
XFILLER_0_102_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09574__X _05516_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12060_ _06626_ net2737 net357 vssd1 vssd1 vccd1 vccd1 _01486_ sky130_fd_sc_hd__mux2_1
Xhold470 team_03_WB.instance_to_wrap.core.register_file.registers_state\[236\] vssd1
+ vssd1 vccd1 vccd1 net1963 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_3020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold481 team_03_WB.instance_to_wrap.core.register_file.registers_state\[750\] vssd1
+ vssd1 vccd1 vccd1 net1974 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07179__A1 net1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout871_X net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_287 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_129_3031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout969_X net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold492 team_03_WB.instance_to_wrap.ADR_I\[17\] vssd1 vssd1 vccd1 vccd1 net1985 sky130_fd_sc_hd__dlygate4sd3_1
X_11011_ net275 net704 net828 vssd1 vssd1 vccd1 vccd1 _06579_ sky130_fd_sc_hd__and3_1
XANTENNA__10183__A0 _04619_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10660__S net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_53_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06926__A1 net1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10722__A2 net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout950 net952 vssd1 vssd1 vccd1 vccd1 net950 sky130_fd_sc_hd__clkbuf_4
Xfanout961 net962 vssd1 vssd1 vccd1 vccd1 net961 sky130_fd_sc_hd__clkbuf_4
Xfanout972 net973 vssd1 vssd1 vccd1 vccd1 net972 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08128__B1 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout983 net994 vssd1 vssd1 vccd1 vccd1 net983 sky130_fd_sc_hd__clkbuf_4
Xfanout994 _04086_ vssd1 vssd1 vccd1 vccd1 net994 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_5_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11057__A net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12962_ net1350 vssd1 vssd1 vccd1 vccd1 _00726_ sky130_fd_sc_hd__inv_2
Xhold1170 team_03_WB.instance_to_wrap.core.register_file.registers_state\[451\] vssd1
+ vssd1 vccd1 vccd1 net2663 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_input10_A DAT_I[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14701_ clknet_leaf_57_wb_clk_i _02465_ _01066_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.ADR_I\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_142_3286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1181 team_03_WB.instance_to_wrap.core.register_file.registers_state\[454\] vssd1
+ vssd1 vccd1 vccd1 net2674 sky130_fd_sc_hd__dlygate4sd3_1
X_11913_ _06614_ net2719 net369 vssd1 vssd1 vccd1 vccd1 _01629_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_142_3297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11683__B1 net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1192 team_03_WB.instance_to_wrap.core.register_file.registers_state\[221\] vssd1
+ vssd1 vccd1 vccd1 net2685 sky130_fd_sc_hd__dlygate4sd3_1
X_12893_ net1384 vssd1 vssd1 vccd1 vccd1 _00657_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_539 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11491__S net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_16_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11844_ _06409_ net2382 net376 vssd1 vssd1 vccd1 vccd1 _01696_ sky130_fd_sc_hd__mux2_1
X_14632_ clknet_leaf_10_wb_clk_i _02396_ _00997_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[986\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__09628__B1 net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_120_2850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14563_ clknet_leaf_47_wb_clk_i _02327_ _00928_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[917\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_28_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_166_950 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07701__C net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11775_ _06608_ net477 net333 net2247 vssd1 vssd1 vccd1 vccd1 _01762_ sky130_fd_sc_hd__a22o_1
XANTENNA__08300__B1 net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10726_ team_03_WB.instance_to_wrap.core.pc.current_pc\[18\] net315 net602 vssd1
+ vssd1 vccd1 vccd1 _06355_ sky130_fd_sc_hd__mux2_1
X_13514_ net1306 vssd1 vssd1 vccd1 vccd1 _01278_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14494_ clknet_leaf_119_wb_clk_i _02258_ _00859_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[848\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_153_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13445_ net1424 vssd1 vssd1 vccd1 vccd1 _01209_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10657_ team_03_WB.instance_to_wrap.core.control_logic.instruction\[4\] team_03_WB.instance_to_wrap.CPU_DAT_O\[4\]
+ net846 vssd1 vssd1 vccd1 vccd1 _02471_ sky130_fd_sc_hd__mux2_1
XANTENNA__09909__B _05563_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11738__A1 net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_828 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload15 clknet_leaf_191_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload15/Y sky130_fd_sc_hd__clkinv_4
Xclkload26 clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload26/Y sky130_fd_sc_hd__inv_8
X_13376_ net1427 vssd1 vssd1 vccd1 vccd1 _01140_ sky130_fd_sc_hd__inv_2
Xclkload37 clknet_leaf_183_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload37/X sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_118_2790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10588_ net1818 net534 net601 _03103_ vssd1 vssd1 vccd1 vccd1 _02535_ sky130_fd_sc_hd__a22o_1
Xclkload48 clknet_leaf_168_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload48/X sky130_fd_sc_hd__clkbuf_8
Xclkload59 clknet_leaf_38_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload59/Y sky130_fd_sc_hd__inv_4
X_15115_ net1486 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[20] sky130_fd_sc_hd__buf_2
XFILLER_0_23_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12327_ net1368 vssd1 vssd1 vccd1 vccd1 _00091_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_77_1959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_149_3429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15046_ net171 vssd1 vssd1 vccd1 vccd1 net169 sky130_fd_sc_hd__clkbuf_1
XANTENNA__09925__A _05646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09159__A2 net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12258_ net1360 vssd1 vssd1 vccd1 vccd1 _00022_ sky130_fd_sc_hd__inv_2
XFILLER_0_103_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11666__S net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11209_ net275 net2379 net487 vssd1 vssd1 vccd1 vccd1 _02199_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_166_3776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12189_ net1687 vssd1 vssd1 vccd1 vccd1 _02364_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_166_3787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06917__A1 net1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07445__A net1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09931__Y _05870_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07164__B _03104_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08975__S net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08828__X _04770_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_46 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07342__A1 net1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08420_ net860 _04358_ _04361_ vssd1 vssd1 vccd1 vccd1 _04362_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_25_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_164_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08351_ _04287_ _04292_ net872 vssd1 vssd1 vccd1 vccd1 _04293_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07302_ _03208_ _03243_ vssd1 vssd1 vccd1 vccd1 _03244_ sky130_fd_sc_hd__and2b_1
XFILLER_0_11_1106 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_611 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08282_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[695\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[663\]
+ net965 vssd1 vssd1 vccd1 vccd1 _04224_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkload9 clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload9/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_116_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07233_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[520\] net796
+ net730 _03174_ vssd1 vssd1 vccd1 vccd1 _03175_ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_93_wb_clk_i clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_93_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_171_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11729__A1 net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11908__D_N net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07164_ _03066_ _03104_ vssd1 vssd1 vccd1 vccd1 _03106_ sky130_fd_sc_hd__nand2_2
Xclkbuf_leaf_22_wb_clk_i clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_22_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08055__C1 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08442__C _04382_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07095_ net1100 team_03_WB.instance_to_wrap.core.register_file.registers_state\[833\]
+ vssd1 vssd1 vccd1 vccd1 _03037_ sky130_fd_sc_hd__and2_1
XANTENNA__08070__A2 net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1037_A net1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11576__S net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08358__B1 net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout497_A net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1204_A net1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11901__A1 net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09570__A2 _05378_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09805_ _05249_ _05250_ vssd1 vssd1 vccd1 vccd1 _05747_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_31_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input2_A DAT_I[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout268 _06541_ vssd1 vssd1 vccd1 vccd1 net268 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_31_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout279 _06418_ vssd1 vssd1 vccd1 vccd1 net279 sky130_fd_sc_hd__buf_2
X_07997_ net750 _03937_ _03938_ vssd1 vssd1 vccd1 vccd1 _03939_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout285_X net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout664_A net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06948_ net615 _02889_ vssd1 vssd1 vccd1 vccd1 _02890_ sky130_fd_sc_hd__or2_1
X_09736_ _05662_ _05677_ net582 vssd1 vssd1 vccd1 vccd1 _05678_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_2_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09667_ net575 _05532_ _05602_ vssd1 vssd1 vccd1 vccd1 _05609_ sky130_fd_sc_hd__o21a_1
X_06879_ _02799_ _02801_ _02810_ _02812_ vssd1 vssd1 vccd1 vccd1 _02821_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout452_X net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout831_A _06558_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07333__A1 net1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout929_A net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_19_Left_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08618_ net1058 team_03_WB.instance_to_wrap.core.register_file.registers_state\[453\]
+ net1011 team_03_WB.instance_to_wrap.core.register_file.registers_state\[485\] net1079
+ vssd1 vssd1 vccd1 vccd1 _04560_ sky130_fd_sc_hd__a221o_1
X_09598_ _05539_ vssd1 vssd1 vccd1 vccd1 _05540_ sky130_fd_sc_hd__inv_2
XANTENNA__11417__A0 _06491_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08549_ net1207 _04483_ _04490_ net849 vssd1 vssd1 vccd1 vccd1 _04491_ sky130_fd_sc_hd__a211o_1
XANTENNA__09086__A1 net1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout717_X net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_211 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11968__A1 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07097__B1 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11560_ net2156 net484 _06794_ net503 vssd1 vssd1 vccd1 vccd1 _01962_ sky130_fd_sc_hd__a22o_1
XANTENNA__12090__B1 net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11043__C net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08473__X _04415_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11432__A3 _06756_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07192__S0 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10511_ net156 net1031 net1023 net1876 vssd1 vssd1 vccd1 vccd1 _02599_ sky130_fd_sc_hd__a22o_1
XFILLER_0_163_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_644 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10655__S net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11491_ _06612_ net2639 net388 vssd1 vssd1 vccd1 vccd1 _02015_ sky130_fd_sc_hd__mux2_1
XFILLER_0_162_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_98_2384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13230_ net1303 vssd1 vssd1 vccd1 vccd1 _00994_ sky130_fd_sc_hd__inv_2
X_10442_ _05925_ _05945_ _06259_ vssd1 vssd1 vccd1 vccd1 _06260_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_123_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_2395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08597__B1 net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13161_ net1256 vssd1 vssd1 vccd1 vccd1 _00925_ sky130_fd_sc_hd__inv_2
X_10373_ team_03_WB.instance_to_wrap.core.pc.current_pc\[20\] _06145_ vssd1 vssd1
+ vccd1 vccd1 _06204_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_33_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12112_ net1143 net1624 net1784 _06282_ vssd1 vssd1 vccd1 vccd1 _00004_ sky130_fd_sc_hd__a22o_1
XFILLER_0_27_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input58_A gpio_in[33] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13092_ net1385 vssd1 vssd1 vccd1 vccd1 _00856_ sky130_fd_sc_hd__inv_2
X_12043_ _06612_ net2709 net355 vssd1 vssd1 vccd1 vccd1 _01503_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_72_1856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_3326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07265__A net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07021__B1 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_144_3337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07572__A1 net1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout780 _02851_ vssd1 vssd1 vccd1 vccd1 net780 sky130_fd_sc_hd__buf_4
XFILLER_0_102_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout791 net792 vssd1 vssd1 vccd1 vccd1 net791 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_137_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_14__f_wb_clk_i_A clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_161_3673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13994_ clknet_leaf_0_wb_clk_i _01758_ _00359_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[348\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_161_3684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input13_X net13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12945_ net1274 vssd1 vssd1 vccd1 vccd1 _00709_ sky130_fd_sc_hd__inv_2
XANTENNA__07324__A1 net1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_49 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12876_ net1313 vssd1 vssd1 vccd1 vccd1 _00640_ sky130_fd_sc_hd__inv_2
XFILLER_0_158_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11408__A0 net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14615_ clknet_leaf_110_wb_clk_i _02379_ _00980_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[969\]
+ sky130_fd_sc_hd__dfstp_1
X_11827_ net653 _06659_ net465 net325 net1770 vssd1 vssd1 vccd1 vccd1 _01712_ sky130_fd_sc_hd__a32o_1
XFILLER_0_8_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09077__A1 net1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_157_268 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11959__A1 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_380 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_419 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07088__B1 net1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07627__A2 net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_907 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08824__A1 net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11758_ _06584_ net456 net331 net2193 vssd1 vssd1 vccd1 vccd1 _01779_ sky130_fd_sc_hd__a22o_1
XFILLER_0_55_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14546_ clknet_leaf_164_wb_clk_i _02310_ _00911_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[900\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12081__B1 net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_255 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10709_ _05500_ _05932_ net606 vssd1 vssd1 vccd1 vccd1 _06345_ sky130_fd_sc_hd__or3_1
XFILLER_0_37_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14477_ clknet_leaf_187_wb_clk_i _02241_ _00842_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[831\]
+ sky130_fd_sc_hd__dfrtp_1
X_11689_ _06731_ net380 net338 net2168 vssd1 vssd1 vccd1 vccd1 _01845_ sky130_fd_sc_hd__a22o_1
XANTENNA__12346__A net1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_463 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkload104 clknet_leaf_152_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload104/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_10_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_141_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13428_ net1433 vssd1 vssd1 vccd1 vccd1 _01192_ sky130_fd_sc_hd__inv_2
XFILLER_0_144_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_116_2749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload115 clknet_leaf_159_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload115/Y sky130_fd_sc_hd__inv_8
Xclkload126 clknet_leaf_139_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload126/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_3_525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload137 clknet_leaf_132_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload137/Y sky130_fd_sc_hd__bufinv_16
XANTENNA__11187__A2 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload148 clknet_leaf_114_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload148/Y sky130_fd_sc_hd__clkinv_2
Xclkload159 clknet_leaf_102_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload159/Y sky130_fd_sc_hd__clkinv_2
XTAP_TAPCELL_ROW_168_3816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13359_ net1319 vssd1 vssd1 vccd1 vccd1 _01123_ sky130_fd_sc_hd__inv_2
XFILLER_0_140_157 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08052__A2 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_168_3827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10934__A2 _05730_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07874__S net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07260__B1 net1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07920_ net1147 _03857_ _03859_ _03861_ net720 vssd1 vssd1 vccd1 vccd1 _03862_ sky130_fd_sc_hd__a41o_1
X_15029_ clknet_leaf_101_wb_clk_i _02749_ _01394_ vssd1 vssd1 vccd1 vccd1 net185 sky130_fd_sc_hd__dfrtp_1
XANTENNA__09001__A1 net1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07851_ net1201 team_03_WB.instance_to_wrap.core.register_file.registers_state\[731\]
+ net784 team_03_WB.instance_to_wrap.core.register_file.registers_state\[763\] net751
+ vssd1 vssd1 vccd1 vccd1 _03793_ sky130_fd_sc_hd__o221a_1
XANTENNA__11895__B1 net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_140_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_140_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__07606__C net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07563__A1 net1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07782_ team_03_WB.instance_to_wrap.core.decoder.inst\[12\] _02821_ _03107_ vssd1
+ vssd1 vccd1 vccd1 _03724_ sky130_fd_sc_hd__a21o_2
Xinput2 DAT_I[0] vssd1 vssd1 vccd1 vccd1 net2 sky130_fd_sc_hd__buf_1
XFILLER_0_127_74 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09521_ _04829_ _05462_ net577 vssd1 vssd1 vccd1 vccd1 _05463_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07315__A1 net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08512__B1 net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09452_ _05111_ _05128_ vssd1 vssd1 vccd1 vccd1 _05394_ sky130_fd_sc_hd__nor2_1
XFILLER_0_149_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07622__B net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_818 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_758 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08403_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[569\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[537\]
+ net992 vssd1 vssd1 vccd1 vccd1 _04345_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09383_ _05323_ _05324_ vssd1 vssd1 vccd1 vccd1 _05325_ sky130_fd_sc_hd__and2b_1
XANTENNA__09068__A1 net1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08334_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[821\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[789\]
+ net969 vssd1 vssd1 vccd1 vccd1 _04276_ sky130_fd_sc_hd__mux2_1
XANTENNA__08276__C1 net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06953__S net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08815__A1 net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08293__X _04235_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10983__B net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10083__C1 _05082_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10622__A1 team_03_WB.instance_to_wrap.CPU_DAT_O\[7\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_74_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08265_ _04193_ _04206_ net850 vssd1 vssd1 vccd1 vccd1 _04207_ sky130_fd_sc_hd__mux2_8
XFILLER_0_28_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_288 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout412_A _06635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1154_A net1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11160__A net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07216_ _03156_ _03157_ net740 vssd1 vssd1 vccd1 vccd1 _03158_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08196_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[563\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[531\]
+ net959 vssd1 vssd1 vccd1 vccd1 _04138_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08579__B1 net1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_770 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07147_ net1103 team_03_WB.instance_to_wrap.core.register_file.registers_state\[192\]
+ net800 team_03_WB.instance_to_wrap.core.register_file.registers_state\[224\] net735
+ vssd1 vssd1 vccd1 vccd1 _03089_ sky130_fd_sc_hd__a221o_1
XFILLER_0_160_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08237__C_N _04178_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10925__A2 _06511_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1419_A net1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07251__B1 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_2281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07078_ net1131 _03018_ net1164 vssd1 vssd1 vccd1 vccd1 _03020_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_93_2292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout781_A net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout879_A net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10138__A0 _04119_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13087__A net1347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1008 _04085_ vssd1 vssd1 vccd1 vccd1 net1008 sky130_fd_sc_hd__clkbuf_4
Xfanout1019 net1022 vssd1 vssd1 vccd1 vccd1 net1019 sky130_fd_sc_hd__buf_4
XANTENNA_fanout1207_X net1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11886__B1 net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout667_X net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11350__A2 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07372__X _03314_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_27_Left_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09719_ _05239_ _05271_ _05273_ _05231_ vssd1 vssd1 vccd1 vccd1 _05661_ sky130_fd_sc_hd__a31o_1
XANTENNA__11638__B1 net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout834_X net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10991_ net1247 net832 _06414_ net668 vssd1 vssd1 vccd1 vccd1 _06567_ sky130_fd_sc_hd__or4_1
XANTENNA__07306__A1 net1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11335__A net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12730_ net1380 vssd1 vssd1 vccd1 vccd1 _00494_ sky130_fd_sc_hd__inv_2
XFILLER_0_85_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_48_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10861__A1 net1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12661_ net1275 vssd1 vssd1 vccd1 vccd1 _00425_ sky130_fd_sc_hd__inv_2
X_14400_ clknet_leaf_192_wb_clk_i _02164_ _00765_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[754\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_65_531 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11612_ _06686_ net381 net346 net2339 vssd1 vssd1 vccd1 vccd1 _01920_ sky130_fd_sc_hd__a22o_1
XANTENNA__12063__A0 _06628_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12592_ net1400 vssd1 vssd1 vccd1 vccd1 _00356_ sky130_fd_sc_hd__inv_2
XFILLER_0_136_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10613__A1 team_03_WB.instance_to_wrap.CPU_DAT_O\[16\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_11543_ net490 net618 _06653_ net482 net1834 vssd1 vssd1 vccd1 vccd1 _01972_ sky130_fd_sc_hd__a32o_1
X_14331_ clknet_leaf_122_wb_clk_i _02095_ _00696_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[685\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_93_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_3185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11810__B1 net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_3196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11070__A net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_36_Left_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14262_ clknet_leaf_178_wb_clk_i _02026_ _00627_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[616\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08019__C1 net1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_102 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11474_ net2680 net393 _06772_ net503 vssd1 vssd1 vccd1 vccd1 _02026_ sky130_fd_sc_hd__a22o_1
XANTENNA__07490__B1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_647 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11169__A2 net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13213_ net1388 vssd1 vssd1 vccd1 vccd1 _00977_ sky130_fd_sc_hd__inv_2
X_10425_ team_03_WB.instance_to_wrap.core.pc.current_pc\[10\] _06138_ vssd1 vssd1
+ vccd1 vccd1 _06246_ sky130_fd_sc_hd__nor2_1
XFILLER_0_34_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14193_ clknet_leaf_143_wb_clk_i _01957_ _00558_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[547\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_74_1907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10916__A2 net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07547__X _03489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13144_ net1375 vssd1 vssd1 vccd1 vccd1 _00908_ sky130_fd_sc_hd__inv_2
X_10356_ _06098_ _06189_ vssd1 vssd1 vccd1 vccd1 _06190_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09782__A2 _05638_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_2646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_111_2657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07793__A1 net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_11__f_wb_clk_i clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_11__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_103_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08990__B1 net995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13075_ net1267 vssd1 vssd1 vccd1 vccd1 _00839_ sky130_fd_sc_hd__inv_2
X_10287_ _04475_ _02766_ net673 vssd1 vssd1 vccd1 vccd1 _06129_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_163_3713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_163_3724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12026_ _06768_ net469 net361 net2720 vssd1 vssd1 vccd1 vccd1 _01519_ sky130_fd_sc_hd__a22o_1
XANTENNA__09534__A2 _04777_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11877__B1 net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07426__C net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07545__A1 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08742__B1 net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_45_Left_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09922__B _05541_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07640__S1 net1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11892__A3 net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11629__B1 net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13977_ clknet_leaf_154_wb_clk_i _01741_ _00342_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[331\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10787__C net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11245__A net1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12928_ net1402 vssd1 vssd1 vccd1 vccd1 _00692_ sky130_fd_sc_hd__inv_2
XFILLER_0_88_678 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10852__A1 team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[20\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12859_ net1360 vssd1 vssd1 vccd1 vccd1 _00623_ sky130_fd_sc_hd__inv_2
XFILLER_0_173_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_43 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_154_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14529_ clknet_leaf_180_wb_clk_i _02293_ _00894_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[883\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09470__A1 net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07076__A3 net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_154_772 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08050_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[22\] net771
+ net755 _03991_ vssd1 vssd1 vccd1 vccd1 _03992_ sky130_fd_sc_hd__a211o_1
XFILLER_0_113_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07001_ _02939_ _02941_ _02942_ vssd1 vssd1 vccd1 vccd1 _02943_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_98_56 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_308 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09385__A _04267_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07233__B1 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14999__Q team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[18\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08430__C1 net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08952_ net436 net428 _04893_ vssd1 vssd1 vccd1 vccd1 _04894_ sky130_fd_sc_hd__nor3_1
XANTENNA__11868__A0 _06527_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07903_ net1090 team_03_WB.instance_to_wrap.core.register_file.registers_state\[591\]
+ net794 team_03_WB.instance_to_wrap.core.register_file.registers_state\[623\] net755
+ vssd1 vssd1 vccd1 vccd1 _03845_ sky130_fd_sc_hd__a221o_1
X_08883_ net434 net429 _04807_ vssd1 vssd1 vccd1 vccd1 _04825_ sky130_fd_sc_hd__or3_1
XANTENNA__11854__S net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08733__B1 net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07834_ net821 _03775_ net721 vssd1 vssd1 vccd1 vccd1 _03776_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10540__B1 net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11883__A3 net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07765_ net1098 team_03_WB.instance_to_wrap.core.register_file.registers_state\[748\]
+ net883 _03706_ net1155 vssd1 vssd1 vccd1 vccd1 _03707_ sky130_fd_sc_hd__o2111a_1
XANTENNA_fanout362_A _06817_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11155__A net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09504_ _03823_ _04444_ net665 _05445_ vssd1 vssd1 vccd1 vccd1 _05446_ sky130_fd_sc_hd__a22o_1
XFILLER_0_155_1086 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_154_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07696_ _03620_ _03621_ _03629_ _03637_ vssd1 vssd1 vccd1 vccd1 _03638_ sky130_fd_sc_hd__o22a_4
XANTENNA__08497__C1 net1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_13__f_wb_clk_i_X clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_116_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09435_ _05375_ _05376_ net558 vssd1 vssd1 vccd1 vccd1 _05377_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10994__A net1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1271_A net1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout627_A net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1369_A net1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09366_ _05185_ _05191_ vssd1 vssd1 vccd1 vccd1 _05308_ sky130_fd_sc_hd__and2_1
XFILLER_0_118_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_23_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08317_ net1237 team_03_WB.instance_to_wrap.core.register_file.registers_state\[984\]
+ net973 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1016\] net1220
+ vssd1 vssd1 vccd1 vccd1 _04259_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_43_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_586 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_43_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09297_ _04619_ _05238_ vssd1 vssd1 vccd1 vccd1 _05239_ sky130_fd_sc_hd__or2_2
XFILLER_0_151_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout415_X net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1157_X net1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09994__S net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_400 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_2321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08248_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[434\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[402\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[306\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[274\]
+ net951 net1070 vssd1 vssd1 vccd1 vccd1 _04190_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_95_2332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout996_A net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_162_1024 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08179_ net548 _04120_ vssd1 vssd1 vccd1 vccd1 _04121_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_132_3082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_3093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10210_ _02889_ _06039_ vssd1 vssd1 vccd1 vccd1 _06052_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07224__B1 net1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07808__A net1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08403__S net992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11190_ net655 net705 net268 net697 vssd1 vssd1 vccd1 vccd1 _06676_ sky130_fd_sc_hd__and4_1
XANTENNA__08421__C1 net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_1127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout784_X net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11571__A2 net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10141_ _05981_ _05982_ vssd1 vssd1 vccd1 vccd1 _05983_ sky130_fd_sc_hd__and2_1
XFILLER_0_24_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput180 net180 vssd1 vssd1 vccd1 vccd1 gpio_oeb[15] sky130_fd_sc_hd__buf_2
Xoutput191 net191 vssd1 vssd1 vccd1 vccd1 gpio_oeb[26] sky130_fd_sc_hd__clkbuf_4
XANTENNA__07019__S net1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11859__A0 _06487_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10072_ _02811_ _02830_ _02833_ vssd1 vssd1 vccd1 vccd1 _05916_ sky130_fd_sc_hd__nor3_1
XANTENNA__11049__B net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13900_ clknet_leaf_19_wb_clk_i _01664_ _00265_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[254\]
+ sky130_fd_sc_hd__dfrtp_1
X_14880_ clknet_leaf_83_wb_clk_i _02643_ _01245_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.pc.current_pc\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10531__B1 net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13831_ clknet_leaf_109_wb_clk_i _01595_ _00196_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[185\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09819__A3 net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10974_ net312 _05845_ net318 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[0\]
+ vssd1 vssd1 vccd1 vccd1 _06553_ sky130_fd_sc_hd__a31o_1
X_13762_ clknet_leaf_174_wb_clk_i _01526_ _00127_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[116\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_67_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10834__A1 net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_139_3225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12713_ net1253 vssd1 vssd1 vccd1 vccd1 _00477_ sky130_fd_sc_hd__inv_2
XFILLER_0_70_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_139_3236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_339 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13693_ clknet_leaf_27_wb_clk_i _01457_ _00058_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[47\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_155_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12036__B1 net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12644_ net1366 vssd1 vssd1 vccd1 vccd1 _00408_ sky130_fd_sc_hd__inv_2
XFILLER_0_84_158 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_156_3572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_156_3583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12575_ net1285 vssd1 vssd1 vccd1 vccd1 _00339_ sky130_fd_sc_hd__inv_2
XFILLER_0_53_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_142_219 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14314_ clknet_leaf_5_wb_clk_i _02078_ _00679_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[668\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11526_ net649 _06638_ vssd1 vssd1 vccd1 vccd1 _06782_ sky130_fd_sc_hd__nor2_1
XFILLER_0_108_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08660__C1 team_03_WB.instance_to_wrap.core.decoder.inst\[17\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xwire274 _06453_ vssd1 vssd1 vccd1 vccd1 net274 sky130_fd_sc_hd__buf_4
XANTENNA__11939__S net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11457_ net490 net618 _06582_ net392 net2059 vssd1 vssd1 vccd1 vccd1 _02036_ sky130_fd_sc_hd__a32o_1
X_14245_ clknet_leaf_40_wb_clk_i _02009_ _00610_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[599\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09917__B _05852_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12624__A net1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10408_ team_03_WB.instance_to_wrap.core.pc.current_pc\[14\] net681 _06230_ _06232_
+ vssd1 vssd1 vccd1 vccd1 _02648_ sky130_fd_sc_hd__o22a_1
XFILLER_0_141_1108 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_639 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14176_ clknet_leaf_190_wb_clk_i _01940_ _00541_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[530\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08313__S net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11388_ net511 net639 _06746_ net402 net2208 vssd1 vssd1 vccd1 vccd1 _02086_ sky130_fd_sc_hd__a32o_1
XFILLER_0_110_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11562__A2 net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10339_ _06112_ _06115_ vssd1 vssd1 vccd1 vccd1 _06176_ sky130_fd_sc_hd__xnor2_1
X_13127_ net1400 vssd1 vssd1 vccd1 vccd1 _00891_ sky130_fd_sc_hd__inv_2
XANTENNA__10144__A _03109_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06974__C1 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09933__A _03821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13058_ net1289 vssd1 vssd1 vccd1 vccd1 _00822_ sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_4_9__f_wb_clk_i_X clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11674__S net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1350 net1352 vssd1 vssd1 vccd1 vccd1 net1350 sky130_fd_sc_hd__buf_4
X_12009_ _06759_ net453 net359 net2590 vssd1 vssd1 vccd1 vccd1 _01536_ sky130_fd_sc_hd__a22o_1
Xfanout1361 net1363 vssd1 vssd1 vccd1 vccd1 net1361 sky130_fd_sc_hd__buf_4
XANTENNA__10522__B1 net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1372 net1373 vssd1 vssd1 vccd1 vccd1 net1372 sky130_fd_sc_hd__buf_4
XANTENNA__08191__A1 net1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1383 net1384 vssd1 vssd1 vccd1 vccd1 net1383 sky130_fd_sc_hd__buf_4
XFILLER_0_75_1025 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1394 net1396 vssd1 vssd1 vccd1 vccd1 net1394 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_128_2995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07550_ net1200 team_03_WB.instance_to_wrap.core.register_file.registers_state\[56\]
+ net886 vssd1 vssd1 vccd1 vccd1 _03492_ sky130_fd_sc_hd__and3_1
XANTENNA_clkbuf_leaf_34_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__08479__C1 net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10825__A1 team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[25\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07481_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[917\] net793
+ _03422_ vssd1 vssd1 vccd1 vccd1 _03423_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_5_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_159_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09220_ _03280_ _03314_ _05160_ net607 vssd1 vssd1 vccd1 vccd1 _05162_ sky130_fd_sc_hd__a31o_1
XANTENNA__13190__A net1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12027__B1 net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_106 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09151_ net575 _05092_ vssd1 vssd1 vccd1 vccd1 _05093_ sky130_fd_sc_hd__nand2_1
XFILLER_0_57_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09443__A1 _05384_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08102_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[442\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[410\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[314\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[282\]
+ net759 net1124 vssd1 vssd1 vccd1 vccd1 _04044_ sky130_fd_sc_hd__mux4_1
XFILLER_0_173_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09082_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[429\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[397\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[301\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[269\]
+ net982 net1076 vssd1 vssd1 vccd1 vccd1 _05024_ sky130_fd_sc_hd__mux4_1
XANTENNA__11250__A1 net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11849__S net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08033_ net1178 team_03_WB.instance_to_wrap.core.register_file.registers_state\[465\]
+ vssd1 vssd1 vccd1 vccd1 _03975_ sky130_fd_sc_hd__or2_1
Xinput60 gpio_in[35] vssd1 vssd1 vccd1 vccd1 net60 sky130_fd_sc_hd__clkbuf_1
Xhold800 team_03_WB.instance_to_wrap.core.register_file.registers_state\[373\] vssd1
+ vssd1 vccd1 vccd1 net2293 sky130_fd_sc_hd__dlygate4sd3_1
Xinput71 wbs_adr_i[13] vssd1 vssd1 vccd1 vccd1 net71 sky130_fd_sc_hd__buf_1
XFILLER_0_114_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold811 team_03_WB.instance_to_wrap.core.register_file.registers_state\[375\] vssd1
+ vssd1 vccd1 vccd1 net2304 sky130_fd_sc_hd__dlygate4sd3_1
Xinput82 wbs_adr_i[23] vssd1 vssd1 vccd1 vccd1 net82 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold822 team_03_WB.instance_to_wrap.core.register_file.registers_state\[322\] vssd1
+ vssd1 vccd1 vccd1 net2315 sky130_fd_sc_hd__dlygate4sd3_1
Xinput93 wbs_adr_i[4] vssd1 vssd1 vccd1 vccd1 net93 sky130_fd_sc_hd__clkbuf_1
XANTENNA__11002__B2 net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold833 team_03_WB.instance_to_wrap.core.register_file.registers_state\[108\] vssd1
+ vssd1 vccd1 vccd1 net2326 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07628__A net1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold844 team_03_WB.instance_to_wrap.core.register_file.registers_state\[331\] vssd1
+ vssd1 vccd1 vccd1 net2337 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08223__S net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold855 team_03_WB.instance_to_wrap.core.register_file.registers_state\[378\] vssd1
+ vssd1 vccd1 vccd1 net2348 sky130_fd_sc_hd__dlygate4sd3_1
Xhold866 team_03_WB.instance_to_wrap.core.register_file.registers_state\[127\] vssd1
+ vssd1 vccd1 vccd1 net2359 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07757__A1 net1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11553__A2 net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold877 team_03_WB.instance_to_wrap.core.register_file.registers_state\[350\] vssd1
+ vssd1 vccd1 vccd1 net2370 sky130_fd_sc_hd__dlygate4sd3_1
Xhold888 team_03_WB.instance_to_wrap.core.register_file.registers_state\[339\] vssd1
+ vssd1 vccd1 vccd1 net2381 sky130_fd_sc_hd__dlygate4sd3_1
X_09984_ _05869_ net1862 net289 vssd1 vssd1 vccd1 vccd1 _02730_ sky130_fd_sc_hd__mux2_1
Xhold899 team_03_WB.instance_to_wrap.core.register_file.registers_state\[530\] vssd1
+ vssd1 vccd1 vccd1 net2392 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10761__B1 net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06965__C1 net1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1117_A _02786_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08935_ _04875_ _04876_ net868 vssd1 vssd1 vccd1 vccd1 _04877_ sky130_fd_sc_hd__a21o_1
XANTENNA__10989__A net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_73_wb_clk_i_A clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout577_A _02993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11584__S net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13365__A net1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10513__B1 net1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08866_ net545 _04807_ vssd1 vssd1 vccd1 vccd1 _04808_ sky130_fd_sc_hd__nand2_1
XANTENNA__08182__A1 net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08459__A net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07817_ _03756_ _03758_ net611 vssd1 vssd1 vccd1 vccd1 _03759_ sky130_fd_sc_hd__mux2_1
X_08797_ net848 _04738_ _04727_ vssd1 vssd1 vccd1 vccd1 _04739_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_88_2180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07390__C1 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout365_X net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_2191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout744_A net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09989__S net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07748_ net1195 team_03_WB.instance_to_wrap.core.register_file.registers_state\[204\]
+ vssd1 vssd1 vccd1 vccd1 _03690_ sky130_fd_sc_hd__or2_1
XANTENNA__08893__S net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_45_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout532_X net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07679_ net821 _03614_ net717 vssd1 vssd1 vccd1 vccd1 _03621_ sky130_fd_sc_hd__o21ai_1
XANTENNA__12709__A net1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_823 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09418_ _04268_ _04355_ vssd1 vssd1 vccd1 vccd1 _05360_ sky130_fd_sc_hd__nor2_1
XANTENNA__12018__B1 net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10690_ team_03_WB.instance_to_wrap.core.pc.current_pc\[29\] _06317_ vssd1 vssd1
+ vccd1 vccd1 _06330_ sky130_fd_sc_hd__nand2_1
XFILLER_0_54_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07693__B1 net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09349_ _05285_ _05290_ vssd1 vssd1 vccd1 vccd1 _05291_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_134_3122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_134_3133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07586__A_N net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_934 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12360_ net1291 vssd1 vssd1 vccd1 vccd1 _00124_ sky130_fd_sc_hd__inv_2
XANTENNA__11051__C net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout999_X net999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11311_ _06454_ net2531 net404 vssd1 vssd1 vccd1 vccd1 _02134_ sky130_fd_sc_hd__mux2_1
XANTENNA__07996__A1 net1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_151_3480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09737__B _04953_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12291_ net1371 vssd1 vssd1 vccd1 vccd1 _00055_ sky130_fd_sc_hd__inv_2
XFILLER_0_62_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14030_ clknet_leaf_127_wb_clk_i _01794_ _00395_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[384\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_121_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11242_ net491 net619 _06688_ net408 net2125 vssd1 vssd1 vccd1 vccd1 _02174_ sky130_fd_sc_hd__a32o_1
XFILLER_0_30_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11173_ net1044 net836 net270 net668 vssd1 vssd1 vccd1 vccd1 _06666_ sky130_fd_sc_hd__and4_1
XFILLER_0_38_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06956__C1 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input40_A gpio_in[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10124_ team_03_WB.instance_to_wrap.core.pc.current_pc\[29\] net672 vssd1 vssd1 vccd1
+ vccd1 _05966_ sky130_fd_sc_hd__nand2_1
XFILLER_0_100_182 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11494__S net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14932_ clknet_leaf_44_wb_clk_i _02687_ _01297_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_O\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_10055_ net32 net1039 net911 team_03_WB.instance_to_wrap.CPU_DAT_O\[8\] vssd1 vssd1
+ vccd1 vccd1 _02676_ sky130_fd_sc_hd__a22o_1
XANTENNA__10504__B1 net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08173__A1 net1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14863_ clknet_leaf_64_wb_clk_i net1766 _01228_ vssd1 vssd1 vccd1 vccd1 net119 sky130_fd_sc_hd__dfrtp_1
XANTENNA__07920__A1 net1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_2545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13814_ clknet_leaf_154_wb_clk_i _01578_ _00179_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[168\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_159_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14794_ clknet_leaf_84_wb_clk_i _02558_ _01159_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_I\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_158_3612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_626 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_158_3623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13745_ clknet_leaf_140_wb_clk_i _01509_ _00110_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[99\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_74_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_423 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10957_ team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[3\] net308 net688 vssd1
+ vssd1 vccd1 vccd1 _06539_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_123_2892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11082__X _06619_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12009__B1 net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07684__B1 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11480__A1 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13676_ clknet_leaf_5_wb_clk_i _01440_ _00041_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_118_wb_clk_i_A clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_167_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10888_ _06480_ _06481_ _06482_ net586 vssd1 vssd1 vccd1 vccd1 _06483_ sky130_fd_sc_hd__o211a_2
XFILLER_0_94_990 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12627_ net1255 vssd1 vssd1 vccd1 vccd1 _00391_ sky130_fd_sc_hd__inv_2
XANTENNA__09425__A1 net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10139__A _03390_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08859__S0 net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09487__X _05429_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07436__B1 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_171_3878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_720 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08633__C1 net1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12558_ net1310 vssd1 vssd1 vccd1 vccd1 _00322_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_171_3889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07987__A1 net1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_526 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11669__S net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11509_ _06505_ net2501 net390 vssd1 vssd1 vccd1 vccd1 _01997_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_151_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_1041 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12489_ net1254 vssd1 vssd1 vccd1 vccd1 _00253_ sky130_fd_sc_hd__inv_2
XFILLER_0_79_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold107 team_03_WB.instance_to_wrap.CPU_DAT_I\[3\] vssd1 vssd1 vccd1 vccd1 net1600
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold118 team_03_WB.instance_to_wrap.ADR_I\[9\] vssd1 vssd1 vccd1 vccd1 net1611 sky130_fd_sc_hd__dlygate4sd3_1
Xhold129 team_03_WB.instance_to_wrap.CPU_DAT_I\[6\] vssd1 vssd1 vccd1 vccd1 net1622
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11941__D_N net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14228_ clknet_leaf_132_wb_clk_i _01992_ _00593_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[582\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_88 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08936__B1 net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11535__A2 net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_283 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14159_ clknet_leaf_134_wb_clk_i _01923_ _00524_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[513\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10743__B1 net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout609 _02938_ vssd1 vssd1 vccd1 vccd1 net609 sky130_fd_sc_hd__buf_4
XFILLER_0_120_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09663__A net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06981_ net615 _02921_ _02922_ vssd1 vssd1 vccd1 vccd1 _02923_ sky130_fd_sc_hd__a21oi_2
X_08720_ net1067 _04660_ _04661_ vssd1 vssd1 vccd1 vccd1 _04662_ sky130_fd_sc_hd__a21o_1
Xclkbuf_leaf_47_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_47_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_119_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08279__A net1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1180 net1206 vssd1 vssd1 vccd1 vccd1 net1180 sky130_fd_sc_hd__clkbuf_4
X_08651_ net435 net430 _04592_ net545 vssd1 vssd1 vccd1 vccd1 _04593_ sky130_fd_sc_hd__o31a_1
Xfanout1191 net1193 vssd1 vssd1 vccd1 vccd1 net1191 sky130_fd_sc_hd__clkbuf_4
XANTENNA_clkbuf_leaf_157_wb_clk_i_A clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_07602_ net1135 _03539_ _03540_ _03542_ net1121 vssd1 vssd1 vccd1 vccd1 _03544_ sky130_fd_sc_hd__a311o_1
XFILLER_0_117_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08582_ net937 _04523_ _04522_ net1064 vssd1 vssd1 vccd1 vccd1 _04524_ sky130_fd_sc_hd__o211a_1
XFILLER_0_152_1023 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11136__C net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_1131 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07533_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[166\] net779
+ net747 _03474_ vssd1 vssd1 vccd1 vccd1 _03475_ sky130_fd_sc_hd__o211a_1
XANTENNA__08011__S1 net1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_171 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07464_ net1116 _03402_ _03403_ vssd1 vssd1 vccd1 vccd1 _03406_ sky130_fd_sc_hd__or3_1
XFILLER_0_36_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09203_ net526 _03491_ _05144_ vssd1 vssd1 vccd1 vccd1 _05145_ sky130_fd_sc_hd__and3_1
XFILLER_0_146_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07395_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[703\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[671\]
+ net763 vssd1 vssd1 vccd1 vccd1 _03337_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_40_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_180 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout325_A _06811_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09134_ net526 _02948_ _05075_ vssd1 vssd1 vccd1 vccd1 _05076_ sky130_fd_sc_hd__and3_1
XFILLER_0_8_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1067_A net1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09838__A net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07427__B1 net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10991__B net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07522__S0 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11774__A2 net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11579__S net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09065_ net1048 team_03_WB.instance_to_wrap.core.register_file.registers_state\[975\]
+ net999 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1007\] net921
+ vssd1 vssd1 vccd1 vccd1 _05007_ sky130_fd_sc_hd__a221o_1
XFILLER_0_130_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1234_A net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08016_ net1085 team_03_WB.instance_to_wrap.core.register_file.registers_state\[689\]
+ net890 vssd1 vssd1 vccd1 vccd1 _03958_ sky130_fd_sc_hd__or3_1
XFILLER_0_114_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold630 team_03_WB.instance_to_wrap.core.register_file.registers_state\[56\] vssd1
+ vssd1 vccd1 vccd1 net2123 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold641 team_03_WB.instance_to_wrap.core.register_file.registers_state\[754\] vssd1
+ vssd1 vccd1 vccd1 net2134 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout694_A _06562_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08927__B1 net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold652 team_03_WB.instance_to_wrap.core.register_file.registers_state\[740\] vssd1
+ vssd1 vccd1 vccd1 net2145 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold663 team_03_WB.instance_to_wrap.core.register_file.registers_state\[552\] vssd1
+ vssd1 vccd1 vccd1 net2156 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold674 team_03_WB.instance_to_wrap.core.register_file.registers_state\[738\] vssd1
+ vssd1 vccd1 vccd1 net2167 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1022_X net1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold685 team_03_WB.instance_to_wrap.core.register_file.registers_state\[779\] vssd1
+ vssd1 vccd1 vccd1 net2178 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1401_A net1408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold696 team_03_WB.instance_to_wrap.core.register_file.registers_state\[390\] vssd1
+ vssd1 vccd1 vccd1 net2189 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07792__S net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09967_ _03788_ net663 vssd1 vssd1 vccd1 vccd1 _05888_ sky130_fd_sc_hd__nor2_2
XANTENNA_fanout861_A net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout482_X net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout959_A net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11608__A net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10071__X _05915_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08918_ net868 _04859_ _04854_ net852 vssd1 vssd1 vccd1 vccd1 _04860_ sky130_fd_sc_hd__o211a_1
X_09898_ _05355_ _05397_ _05403_ _05513_ vssd1 vssd1 vccd1 vccd1 _05840_ sky130_fd_sc_hd__a22o_1
XFILLER_0_99_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_86_2139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08849_ net1068 _04790_ vssd1 vssd1 vccd1 vccd1 _04791_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout747_X net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07902__A1 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11860_ net271 net2118 net377 vssd1 vssd1 vccd1 vccd1 _01680_ sky130_fd_sc_hd__mux2_1
XFILLER_0_170_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09104__B1 net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10811_ _06415_ _06416_ _06417_ vssd1 vssd1 vccd1 vccd1 _06418_ sky130_fd_sc_hd__a21oi_4
XTAP_TAPCELL_ROW_0_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10658__S net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11791_ net2237 _06479_ net328 vssd1 vssd1 vccd1 vccd1 _01747_ sky130_fd_sc_hd__mux2_1
XANTENNA__09655__A1 _05278_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11343__A net1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13530_ net1306 vssd1 vssd1 vccd1 vccd1 _01294_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07666__B1 net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_2442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10742_ team_03_WB.instance_to_wrap.core.pc.current_pc\[10\] _05686_ net605 vssd1
+ vssd1 vccd1 vccd1 _06363_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_101_2453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11462__B2 net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13461_ net1323 vssd1 vssd1 vccd1 vccd1 _01225_ sky130_fd_sc_hd__inv_2
X_10673_ team_03_WB.instance_to_wrap.core.pc.current_pc\[25\] team_03_WB.instance_to_wrap.core.pc.current_pc\[24\]
+ vssd1 vssd1 vccd1 vccd1 _06315_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_153_3520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_11_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_173_Right_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_168_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12412_ net1411 vssd1 vssd1 vccd1 vccd1 _00176_ sky130_fd_sc_hd__inv_2
XANTENNA__07418__B1 net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08615__C1 net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11214__B2 net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13392_ net1433 vssd1 vssd1 vccd1 vccd1 _01156_ sky130_fd_sc_hd__inv_2
XANTENNA_input88_A wbs_adr_i[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_591 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_347 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_168_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11489__S net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12343_ net1390 vssd1 vssd1 vccd1 vccd1 _00107_ sky130_fd_sc_hd__inv_2
XFILLER_0_65_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07268__A net1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15062_ net1448 vssd1 vssd1 vccd1 vccd1 irq[1] sky130_fd_sc_hd__buf_2
X_12274_ net1397 vssd1 vssd1 vccd1 vccd1 _00038_ sky130_fd_sc_hd__inv_2
XFILLER_0_49_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_79_1990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11225_ net2771 net486 _06683_ net494 vssd1 vssd1 vccd1 vccd1 _02186_ sky130_fd_sc_hd__a22o_1
X_14013_ clknet_leaf_25_wb_clk_i _01777_ _00378_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[367\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10725__B1 net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12902__A net1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08394__A1 net1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11156_ net2175 net412 _06655_ net501 vssd1 vssd1 vccd1 vccd1 _02227_ sky130_fd_sc_hd__a22o_1
XANTENNA__06900__A net1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10107_ team_03_WB.instance_to_wrap.core.pc.current_pc\[1\] net660 vssd1 vssd1 vccd1
+ vccd1 _05951_ sky130_fd_sc_hd__nor2_1
X_11087_ _06469_ net2547 net416 vssd1 vssd1 vccd1 vccd1 _02261_ sky130_fd_sc_hd__mux2_1
XFILLER_0_171_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10038_ net19 net1038 net910 net1785 vssd1 vssd1 vccd1 vccd1 _02693_ sky130_fd_sc_hd__o22a_1
XFILLER_0_136_1007 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14915_ clknet_leaf_43_wb_clk_i _02670_ _01280_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_O\[2\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__11237__B net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14846_ clknet_leaf_85_wb_clk_i _02610_ _01211_ vssd1 vssd1 vccd1 vccd1 net132 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_19_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14777_ clknet_leaf_93_wb_clk_i _02541_ _01142_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_I\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_11989_ _06753_ net462 net443 net2365 vssd1 vssd1 vccd1 vccd1 _01555_ sky130_fd_sc_hd__a22o_1
XFILLER_0_85_231 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11253__A _06442_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_173_3918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13728_ clknet_leaf_191_wb_clk_i _01492_ _00093_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[82\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_173_3929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11453__B2 net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_165_wb_clk_i clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_165_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_105_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07121__A2 _03059_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_156_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13659_ clknet_leaf_145_wb_clk_i _01423_ _00024_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_140_Right_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07409__B1 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07180_ _03116_ _03121_ net821 vssd1 vssd1 vccd1 vccd1 _03122_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_170_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08562__A _04503_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11399__S net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08082__B1 net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07424__A3 net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_200 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07178__A net1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08909__B1 net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout406 _06717_ vssd1 vssd1 vccd1 vccd1 net406 sky130_fd_sc_hd__buf_6
X_09821_ net570 _05114_ vssd1 vssd1 vccd1 vccd1 _05763_ sky130_fd_sc_hd__or2_1
Xfanout417 _06610_ vssd1 vssd1 vccd1 vccd1 net417 sky130_fd_sc_hd__buf_4
Xfanout428 net430 vssd1 vssd1 vccd1 vccd1 net428 sky130_fd_sc_hd__buf_2
XANTENNA__08501__S net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout439 _06819_ vssd1 vssd1 vccd1 vccd1 net439 sky130_fd_sc_hd__buf_6
XANTENNA__07593__C1 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09752_ _03727_ net591 _05693_ vssd1 vssd1 vccd1 vccd1 _05694_ sky130_fd_sc_hd__a21oi_1
X_06964_ _02900_ _02905_ net825 vssd1 vssd1 vccd1 vccd1 _02906_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_33_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09680__X _05622_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08703_ _04639_ _04644_ net873 vssd1 vssd1 vccd1 vccd1 _04645_ sky130_fd_sc_hd__mux2_1
X_09683_ _05298_ _05597_ _05296_ vssd1 vssd1 vccd1 vccd1 _05625_ sky130_fd_sc_hd__a21o_1
X_06895_ team_03_WB.instance_to_wrap.core.control_logic.instruction\[6\] net1018 _02836_
+ vssd1 vssd1 vccd1 vccd1 _02837_ sky130_fd_sc_hd__or3_4
XANTENNA__08232__S1 net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout275_A _06446_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11862__S net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10495__A2 net1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08634_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[422\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[390\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[294\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[262\]
+ net983 net1077 vssd1 vssd1 vccd1 vccd1 _04576_ sky130_fd_sc_hd__mux4_1
XANTENNA__07896__B1 net1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10986__B _06562_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08565_ net1235 team_03_WB.instance_to_wrap.core.register_file.registers_state\[189\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[157\] net966 net922
+ vssd1 vssd1 vccd1 vccd1 _04507_ sky130_fd_sc_hd__a221o_1
XANTENNA__09098__C1 net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_2036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout442_A _06819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_81_2047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1184_A net1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07516_ net719 _03441_ _03450_ _03457_ vssd1 vssd1 vccd1 vccd1 _03458_ sky130_fd_sc_hd__o22a_4
X_08496_ net1243 team_03_WB.instance_to_wrap.core.register_file.registers_state\[347\]
+ net987 team_03_WB.instance_to_wrap.core.register_file.registers_state\[379\] net1079
+ vssd1 vssd1 vccd1 vccd1 _04438_ sky130_fd_sc_hd__o221a_1
XANTENNA__11444__B2 net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07112__A2 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10798__A3 net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07447_ net721 _03382_ _03388_ _03373_ vssd1 vssd1 vccd1 vccd1 _03389_ sky130_fd_sc_hd__o31a_4
XANTENNA__11995__A2 net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout707_A net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout328_X net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07378_ net1180 team_03_WB.instance_to_wrap.core.register_file.registers_state\[95\]
+ net758 team_03_WB.instance_to_wrap.core.register_file.registers_state\[127\] net725
+ vssd1 vssd1 vccd1 vccd1 _03320_ sky130_fd_sc_hd__o221a_1
XFILLER_0_33_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09117_ net1222 _05057_ _05058_ vssd1 vssd1 vccd1 vccd1 _05059_ sky130_fd_sc_hd__and3_1
XANTENNA__11610__B net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08073__B1 net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1237_X net1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10955__B1 net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09048_ net1047 team_03_WB.instance_to_wrap.core.register_file.registers_state\[79\]
+ net998 team_03_WB.instance_to_wrap.core.register_file.registers_state\[111\] net939
+ vssd1 vssd1 vccd1 vccd1 _04990_ sky130_fd_sc_hd__a221o_1
XFILLER_0_32_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout697_X net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_57_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold460 team_03_WB.instance_to_wrap.core.register_file.registers_state\[821\] vssd1
+ vssd1 vccd1 vccd1 net1953 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1030 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12722__A net1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10707__B1 net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold471 team_03_WB.instance_to_wrap.CPU_DAT_O\[20\] vssd1 vssd1 vccd1 vccd1 net1964
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_3021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold482 team_03_WB.instance_to_wrap.core.register_file.registers_state\[915\] vssd1
+ vssd1 vccd1 vccd1 net1975 sky130_fd_sc_hd__dlygate4sd3_1
X_11010_ net2314 net421 _06578_ net501 vssd1 vssd1 vccd1 vccd1 _02296_ sky130_fd_sc_hd__a22o_1
XANTENNA__09573__B1 _05384_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_3032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold493 team_03_WB.instance_to_wrap.core.register_file.registers_state\[808\] vssd1
+ vssd1 vccd1 vccd1 net1986 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_53_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout864_X net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11380__B1 net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout940 net943 vssd1 vssd1 vccd1 vccd1 net940 sky130_fd_sc_hd__buf_4
Xfanout951 net952 vssd1 vssd1 vccd1 vccd1 net951 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_95_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout962 net974 vssd1 vssd1 vccd1 vccd1 net962 sky130_fd_sc_hd__buf_2
XFILLER_0_95_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08128__A1 team_03_WB.instance_to_wrap.core.decoder.inst\[26\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout973 net974 vssd1 vssd1 vccd1 vccd1 net973 sky130_fd_sc_hd__buf_2
Xfanout984 net988 vssd1 vssd1 vccd1 vccd1 net984 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_5_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout995 net997 vssd1 vssd1 vccd1 vccd1 net995 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11057__B net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12961_ net1262 vssd1 vssd1 vccd1 vccd1 _00725_ sky130_fd_sc_hd__inv_2
XANTENNA__09876__A1 net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1160 team_03_WB.instance_to_wrap.core.register_file.registers_state\[589\] vssd1
+ vssd1 vccd1 vccd1 net2653 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14700_ clknet_leaf_57_wb_clk_i _02464_ _01065_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.ADR_I\[30\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1171 team_03_WB.instance_to_wrap.core.register_file.registers_state\[607\] vssd1
+ vssd1 vccd1 vccd1 net2664 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09750__B net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11912_ _06613_ net2701 net367 vssd1 vssd1 vccd1 vccd1 _01630_ sky130_fd_sc_hd__mux2_1
Xhold1182 team_03_WB.instance_to_wrap.core.register_file.registers_state\[621\] vssd1
+ vssd1 vccd1 vccd1 net2675 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_142_3287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_142_3298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12892_ net1411 vssd1 vssd1 vccd1 vccd1 _00656_ sky130_fd_sc_hd__inv_2
Xhold1193 team_03_WB.instance_to_wrap.core.register_file.registers_state\[711\] vssd1
+ vssd1 vccd1 vccd1 net2686 sky130_fd_sc_hd__dlygate4sd3_1
X_14631_ clknet_leaf_97_wb_clk_i _02395_ _00996_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[985\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_16_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11843_ net281 net2130 net375 vssd1 vssd1 vccd1 vccd1 _01697_ sky130_fd_sc_hd__mux2_1
XANTENNA__09089__C1 net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_2840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14562_ clknet_leaf_175_wb_clk_i _02326_ _00927_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[916\]
+ sky130_fd_sc_hd__dfrtp_1
X_11774_ _06607_ net471 net333 net2299 vssd1 vssd1 vccd1 vccd1 _01763_ sky130_fd_sc_hd__a22o_1
XANTENNA__08300__A1 net1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_962 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13513_ net1321 vssd1 vssd1 vccd1 vccd1 _01277_ sky130_fd_sc_hd__inv_2
X_10725_ net522 _06353_ _06354_ net527 net1642 vssd1 vssd1 vccd1 vccd1 _02453_ sky130_fd_sc_hd__a32o_1
X_14493_ clknet_leaf_166_wb_clk_i _02257_ _00858_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[847\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_36_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_908 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13444_ net1404 vssd1 vssd1 vccd1 vccd1 _01208_ sky130_fd_sc_hd__inv_2
XFILLER_0_67_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08382__A _04323_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10656_ team_03_WB.instance_to_wrap.core.control_logic.instruction\[5\] team_03_WB.instance_to_wrap.CPU_DAT_O\[5\]
+ net846 vssd1 vssd1 vccd1 vccd1 _02472_ sky130_fd_sc_hd__mux2_1
XANTENNA__11199__A0 net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11738__A2 net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_153_689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkload16 clknet_leaf_192_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload16/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_140_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10587_ net1614 net534 net601 _03059_ vssd1 vssd1 vccd1 vccd1 _02536_ sky130_fd_sc_hd__a22o_1
Xclkload27 clknet_leaf_18_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload27/Y sky130_fd_sc_hd__inv_6
X_13375_ net1416 vssd1 vssd1 vccd1 vccd1 _01139_ sky130_fd_sc_hd__inv_2
XFILLER_0_134_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload38 clknet_leaf_184_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload38/Y sky130_fd_sc_hd__inv_6
XTAP_TAPCELL_ROW_118_2791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload49 clknet_leaf_169_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload49/X sky130_fd_sc_hd__clkbuf_4
X_15114_ net913 vssd1 vssd1 vccd1 vccd1 net247 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_77_1949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07811__B1 net1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12326_ net1332 vssd1 vssd1 vccd1 vccd1 _00090_ sky130_fd_sc_hd__inv_2
X_15045_ net171 vssd1 vssd1 vccd1 vccd1 net168 sky130_fd_sc_hd__clkbuf_1
XANTENNA__09159__A3 _04503_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_17 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09925__B _05676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12257_ net1290 vssd1 vssd1 vccd1 vccd1 _00021_ sky130_fd_sc_hd__inv_2
XANTENNA__12632__A net1376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11208_ net300 net2327 net487 vssd1 vssd1 vccd1 vccd1 _02200_ sky130_fd_sc_hd__mux2_1
X_12188_ net1515 vssd1 vssd1 vccd1 vccd1 _02365_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_166_3777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_166_3788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10152__A _03985_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11139_ net2084 net413 _06645_ net502 vssd1 vssd1 vccd1 vccd1 _02234_ sky130_fd_sc_hd__a22o_1
XANTENNA__08119__A1 net1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09941__A _03900_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09867__A1 net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09867__B2 net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13463__A net1328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07878__B1 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_710 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14829_ clknet_leaf_92_wb_clk_i net1736 _01194_ vssd1 vssd1 vccd1 vccd1 net150 sky130_fd_sc_hd__dfrtp_1
XANTENNA__09619__A1 net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09619__B2 net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07893__A3 net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08350_ net1220 _04290_ _04291_ vssd1 vssd1 vccd1 vccd1 _04292_ sky130_fd_sc_hd__o21a_1
XFILLER_0_58_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07301_ _03241_ _03242_ net612 vssd1 vssd1 vccd1 vccd1 _03243_ sky130_fd_sc_hd__mux2_2
XFILLER_0_129_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08281_ _04217_ _04222_ net872 vssd1 vssd1 vccd1 vccd1 _04223_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07232_ net1096 team_03_WB.instance_to_wrap.core.register_file.registers_state\[552\]
+ net896 vssd1 vssd1 vccd1 vccd1 _03174_ sky130_fd_sc_hd__or3_1
XFILLER_0_143_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_678 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07163_ _03066_ _03104_ vssd1 vssd1 vccd1 vccd1 _03105_ sky130_fd_sc_hd__and2_1
XANTENNA__08055__B1 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07094_ _03027_ _03030_ _03035_ net1118 net1139 vssd1 vssd1 vccd1 vccd1 _03036_ sky130_fd_sc_hd__o221a_1
XANTENNA__07802__B1 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_62_wb_clk_i clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_62_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__09004__C1 net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12542__A net1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08358__A1 net1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11362__B1 net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout392_A net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07566__C1 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09804_ _02954_ _05735_ _05745_ _05733_ vssd1 vssd1 vccd1 vccd1 _05746_ sky130_fd_sc_hd__a211oi_2
XANTENNA__07030__B2 net1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout269 _06532_ vssd1 vssd1 vccd1 vccd1 net269 sky130_fd_sc_hd__buf_2
X_07996_ net1106 team_03_WB.instance_to_wrap.core.register_file.registers_state\[656\]
+ net804 team_03_WB.instance_to_wrap.core.register_file.registers_state\[688\] net734
+ vssd1 vssd1 vccd1 vccd1 _03938_ sky130_fd_sc_hd__a221o_1
XANTENNA__07581__A2 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09735_ _05227_ _05660_ _05217_ vssd1 vssd1 vccd1 vccd1 _05677_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_2_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06947_ team_03_WB.instance_to_wrap.core.decoder.inst\[11\] _02808_ _02818_ team_03_WB.instance_to_wrap.core.decoder.inst\[24\]
+ vssd1 vssd1 vccd1 vccd1 _02889_ sky130_fd_sc_hd__a22o_4
XTAP_TAPCELL_ROW_2_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10997__A net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout657_A net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout278_X net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11592__S net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1399_A net1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09666_ _05513_ _05521_ _05522_ net320 _05607_ vssd1 vssd1 vccd1 vccd1 _05608_ sky130_fd_sc_hd__a221o_1
X_06878_ _02800_ _02802_ _02811_ _02813_ vssd1 vssd1 vccd1 vccd1 _02820_ sky130_fd_sc_hd__o22a_4
X_08617_ net1058 team_03_WB.instance_to_wrap.core.register_file.registers_state\[325\]
+ net1011 team_03_WB.instance_to_wrap.core.register_file.registers_state\[357\] net1216
+ vssd1 vssd1 vccd1 vccd1 _04559_ sky130_fd_sc_hd__a221o_1
XFILLER_0_173_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09597_ _05371_ _05523_ _05538_ vssd1 vssd1 vccd1 vccd1 _05539_ sky130_fd_sc_hd__a21bo_1
XANTENNA_fanout445_X net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout824_A net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1187_X net1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10001__S net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08818__C1 net1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08548_ _04486_ _04489_ net1207 vssd1 vssd1 vccd1 vccd1 _04490_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_148_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07097__A1 net1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout612_X net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08479_ net1243 team_03_WB.instance_to_wrap.core.register_file.registers_state\[603\]
+ net986 team_03_WB.instance_to_wrap.core.register_file.registers_state\[635\] net929
+ vssd1 vssd1 vccd1 vccd1 _04421_ sky130_fd_sc_hd__o221a_1
XFILLER_0_135_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1354_X net1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10510_ net157 net1033 net1025 net1855 vssd1 vssd1 vccd1 vccd1 _02600_ sky130_fd_sc_hd__a22o_1
XANTENNA__07192__S1 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11490_ _06611_ net2636 net389 vssd1 vssd1 vccd1 vccd1 _02016_ sky130_fd_sc_hd__mux2_1
XFILLER_0_163_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08406__S net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10441_ _06028_ _06056_ vssd1 vssd1 vccd1 vccd1 _06259_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_98_2385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_98_2396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08597__A1 net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10372_ net282 _06089_ _06202_ vssd1 vssd1 vccd1 vccd1 _06203_ sky130_fd_sc_hd__and3_1
XFILLER_0_150_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13160_ net1298 vssd1 vssd1 vccd1 vccd1 _00924_ sky130_fd_sc_hd__inv_2
XFILLER_0_103_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout981_X net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08061__A3 net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12111_ net1143 net1578 net1973 _06302_ vssd1 vssd1 vccd1 vccd1 _00003_ sky130_fd_sc_hd__a22o_1
X_13091_ net1371 vssd1 vssd1 vccd1 vccd1 _00855_ sky130_fd_sc_hd__inv_2
XFILLER_0_32_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_4_10__f_wb_clk_i clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_10__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_131_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12452__A net1376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09546__B1 net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12042_ _06611_ net2599 net355 vssd1 vssd1 vccd1 vccd1 _01504_ sky130_fd_sc_hd__mux2_1
Xhold290 _02581_ vssd1 vssd1 vccd1 vccd1 net1783 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10156__A1 net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_1846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11068__A net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_144_3327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07265__B _03206_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_144_3338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout770 net773 vssd1 vssd1 vccd1 vccd1 net770 sky130_fd_sc_hd__buf_2
Xfanout781 net790 vssd1 vssd1 vccd1 vccd1 net781 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11105__A0 _06628_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout792 net795 vssd1 vssd1 vccd1 vccd1 net792 sky130_fd_sc_hd__buf_4
XANTENNA__07309__C1 net1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13993_ clknet_leaf_75_wb_clk_i _01757_ _00358_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[347\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_161_3674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_161_3685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12944_ net1412 vssd1 vssd1 vccd1 vccd1 _00708_ sky130_fd_sc_hd__inv_2
XFILLER_0_172_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08521__A1 net1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08521__B2 net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12875_ net1283 vssd1 vssd1 vccd1 vccd1 _00639_ sky130_fd_sc_hd__inv_2
XFILLER_0_157_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14614_ clknet_leaf_151_wb_clk_i _02378_ _00979_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[968\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_139_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11826_ _06658_ net462 net324 net2258 vssd1 vssd1 vccd1 vccd1 _01713_ sky130_fd_sc_hd__a22o_1
XANTENNA__11234__C net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09904__C_N _05429_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07088__A1 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14545_ clknet_leaf_141_wb_clk_i _02309_ _00910_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[899\]
+ sky130_fd_sc_hd__dfrtp_1
X_11757_ net646 _06582_ net451 net331 net2212 vssd1 vssd1 vccd1 vccd1 _01780_ sky130_fd_sc_hd__a32o_1
XFILLER_0_166_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10708_ _06149_ net603 _06315_ vssd1 vssd1 vccd1 vccd1 _06344_ sky130_fd_sc_hd__or3_1
XFILLER_0_55_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14476_ clknet_leaf_17_wb_clk_i _02240_ _00841_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[830\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_83_587 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11688_ _06730_ net380 net338 net1946 vssd1 vssd1 vccd1 vccd1 _01846_ sky130_fd_sc_hd__a22o_1
XFILLER_0_36_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_475 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkload105 clknet_leaf_153_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload105/Y sky130_fd_sc_hd__bufinv_16
X_13427_ net1415 vssd1 vssd1 vccd1 vccd1 _01191_ sky130_fd_sc_hd__inv_2
X_10639_ net1152 net1806 net844 vssd1 vssd1 vccd1 vccd1 _02489_ sky130_fd_sc_hd__mux2_1
Xclkload116 clknet_leaf_160_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload116/Y sky130_fd_sc_hd__inv_8
Xclkload127 clknet_leaf_140_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload127/Y sky130_fd_sc_hd__clkinv_2
XFILLER_0_144_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkload138 clknet_leaf_133_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload138/Y sky130_fd_sc_hd__clkinv_4
Xclkload149 clknet_leaf_115_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload149/X sky130_fd_sc_hd__clkbuf_4
X_13358_ net1319 vssd1 vssd1 vccd1 vccd1 _01122_ sky130_fd_sc_hd__inv_2
XFILLER_0_80_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_168_3817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10395__A1 net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11592__A0 net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_168_3828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07260__A1 net1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12309_ net1271 vssd1 vssd1 vccd1 vccd1 _00073_ sky130_fd_sc_hd__inv_2
XFILLER_0_122_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13289_ net1322 vssd1 vssd1 vccd1 vccd1 _01053_ sky130_fd_sc_hd__inv_2
X_15028_ clknet_leaf_101_wb_clk_i _02748_ _01393_ vssd1 vssd1 vccd1 vccd1 net184 sky130_fd_sc_hd__dfrtp_1
XANTENNA__07456__A net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_871 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_18_Right_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11344__B1 net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10698__A2 net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07850_ net1108 team_03_WB.instance_to_wrap.core.register_file.registers_state\[827\]
+ net903 vssd1 vssd1 vccd1 vccd1 _03792_ sky130_fd_sc_hd__or3_1
XANTENNA__11895__A1 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07781_ _03700_ _03701_ _03722_ vssd1 vssd1 vccd1 vccd1 _03723_ sky130_fd_sc_hd__o21a_2
XFILLER_0_78_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput3 DAT_I[10] vssd1 vssd1 vccd1 vccd1 net3 sky130_fd_sc_hd__clkbuf_1
X_09520_ net566 _05459_ _05461_ vssd1 vssd1 vccd1 vccd1 _05462_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_127_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_180_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_180_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_09451_ _05391_ _05392_ net555 vssd1 vssd1 vccd1 vccd1 _05393_ sky130_fd_sc_hd__mux2_1
XFILLER_0_149_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07720__C1 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08402_ net1059 team_03_WB.instance_to_wrap.core.register_file.registers_state\[665\]
+ net1012 team_03_WB.instance_to_wrap.core.register_file.registers_state\[697\] net930
+ vssd1 vssd1 vccd1 vccd1 _04344_ sky130_fd_sc_hd__a221o_1
X_09382_ _04354_ _05322_ vssd1 vssd1 vccd1 vccd1 _05324_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_27_Right_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_163_206 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08333_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[949\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[917\]
+ net968 vssd1 vssd1 vccd1 vccd1 _04275_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07079__B2 net1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08276__B1 net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08264_ net867 _04204_ _04205_ vssd1 vssd1 vccd1 vccd1 _04206_ sky130_fd_sc_hd__o21ai_1
X_07215_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[690\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[658\]
+ net756 vssd1 vssd1 vccd1 vccd1 _03157_ sky130_fd_sc_hd__mux2_1
X_08195_ _04135_ _04136_ net860 vssd1 vssd1 vccd1 vccd1 _04137_ sky130_fd_sc_hd__o21a_1
XFILLER_0_104_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout405_A _06717_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1147_A net1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09846__A net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07146_ net1198 team_03_WB.instance_to_wrap.core.register_file.registers_state\[96\]
+ net885 _03087_ vssd1 vssd1 vccd1 vccd1 _03088_ sky130_fd_sc_hd__a31o_1
XFILLER_0_30_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_160_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11583__A0 net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11587__S net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07787__C1 net1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07077_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[418\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[386\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[290\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[258\]
+ net776 net1132 vssd1 vssd1 vccd1 vccd1 _03019_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_93_2282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1314_A net1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_36_Right_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_93_2293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_7_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout774_A net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07539__C1 net1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1009 net1010 vssd1 vssd1 vccd1 vccd1 net1009 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout395_X net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1102_X net1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11886__A1 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout562_X net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout941_A net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07979_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[400\] net804
+ _02869_ _03920_ vssd1 vssd1 vccd1 vccd1 _03921_ sky130_fd_sc_hd__o211a_1
XANTENNA__11038__D net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09718_ _05239_ _05271_ _05273_ _05232_ vssd1 vssd1 vccd1 vccd1 _05660_ sky130_fd_sc_hd__a31o_1
X_10990_ net2672 net420 _06566_ net501 vssd1 vssd1 vccd1 vccd1 _02304_ sky130_fd_sc_hd__a22o_1
XANTENNA__07937__S0 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10846__C1 net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11335__B net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09649_ _03428_ _04295_ net665 _05590_ vssd1 vssd1 vccd1 vccd1 _05591_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_45_Right_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07711__C1 net1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout827_X net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_48_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12660_ net1312 vssd1 vssd1 vccd1 vccd1 _00424_ sky130_fd_sc_hd__inv_2
X_11611_ _06685_ net379 net346 net2312 vssd1 vssd1 vccd1 vccd1 _01921_ sky130_fd_sc_hd__a22o_1
XANTENNA__08267__B1 net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_852 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12591_ net1337 vssd1 vssd1 vccd1 vccd1 _00355_ sky130_fd_sc_hd__inv_2
XFILLER_0_167_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11351__A net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14330_ clknet_leaf_145_wb_clk_i _02094_ _00695_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[684\]
+ sky130_fd_sc_hd__dfrtp_1
X_11542_ net493 net622 _06652_ net482 net1900 vssd1 vssd1 vccd1 vccd1 _01973_ sky130_fd_sc_hd__a32o_1
XFILLER_0_37_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_3186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_3197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11070__B net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14261_ clknet_leaf_105_wb_clk_i _02025_ _00626_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[615\]
+ sky130_fd_sc_hd__dfrtp_1
X_11473_ net653 _06598_ vssd1 vssd1 vccd1 vccd1 _06772_ sky130_fd_sc_hd__nor2_1
XANTENNA_input70_A wbs_adr_i[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13212_ net1419 vssd1 vssd1 vccd1 vccd1 _00976_ sky130_fd_sc_hd__inv_2
X_10424_ team_03_WB.instance_to_wrap.core.pc.current_pc\[11\] _06245_ net682 vssd1
+ vssd1 vccd1 vccd1 _02645_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14192_ clknet_leaf_161_wb_clk_i _01956_ _00557_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[546\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08034__A3 net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07778__C1 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_54_Right_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11497__S net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10916__A3 _06505_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13143_ net1385 vssd1 vssd1 vccd1 vccd1 _00907_ sky130_fd_sc_hd__inv_2
X_10355_ _06100_ _06188_ vssd1 vssd1 vccd1 vccd1 _06189_ sky130_fd_sc_hd__or2_1
XFILLER_0_131_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_111_2647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_2658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08990__A1 net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10286_ _05971_ _05973_ _06126_ _05968_ _05965_ vssd1 vssd1 vccd1 vccd1 _06128_ sky130_fd_sc_hd__a311o_1
XFILLER_0_130_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13074_ net1397 vssd1 vssd1 vccd1 vccd1 _00838_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_163_3714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_163_3725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12025_ net632 _06588_ net464 net361 net1978 vssd1 vssd1 vccd1 vccd1 _01520_ sky130_fd_sc_hd__a32o_1
XANTENNA__11877__A1 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09922__C _05563_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11526__A net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13976_ clknet_leaf_185_wb_clk_i _01740_ _00341_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[330\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_63_Right_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_24_wb_clk_i_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_12927_ net1347 vssd1 vssd1 vccd1 vccd1 _00691_ sky130_fd_sc_hd__inv_2
XANTENNA__11245__B net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10852__A2 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12858_ net1378 vssd1 vssd1 vccd1 vccd1 _00622_ sky130_fd_sc_hd__inv_2
XANTENNA__08835__A net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_212 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11809_ _06634_ _06803_ vssd1 vssd1 vccd1 vccd1 _06811_ sky130_fd_sc_hd__or2_4
XFILLER_0_28_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12789_ net1272 vssd1 vssd1 vccd1 vccd1 _00553_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_1_Left_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_173_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11261__A net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14528_ clknet_leaf_192_wb_clk_i _02292_ _00893_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[882\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_113_77 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10148__Y _05990_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_160_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_784 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14459_ clknet_leaf_121_wb_clk_i _02223_ _00824_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[813\]
+ sky130_fd_sc_hd__dfrtp_1
X_07000_ team_03_WB.instance_to_wrap.core.decoder.inst\[14\] _02928_ _02933_ _02941_
+ vssd1 vssd1 vccd1 vccd1 _02942_ sky130_fd_sc_hd__nand4_1
XPHY_EDGE_ROW_72_Right_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_136 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_68 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10368__A1 net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11565__B1 net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07769__C1 net1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13188__A net1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08430__B1 net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11200__S net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_180 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08951_ net849 _04871_ _04877_ _04892_ vssd1 vssd1 vccd1 vccd1 _04893_ sky130_fd_sc_hd__a31o_4
XANTENNA__11317__A0 _06624_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_63_wb_clk_i_A clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_138_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07902_ net817 _03833_ _03843_ vssd1 vssd1 vccd1 vccd1 _03844_ sky130_fd_sc_hd__a21oi_1
X_08882_ _04080_ _04807_ vssd1 vssd1 vccd1 vccd1 _04824_ sky130_fd_sc_hd__nor2_1
XANTENNA__08194__C1 net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08733__A1 net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07833_ _03773_ _03774_ net1114 vssd1 vssd1 vccd1 vccd1 _03775_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_81_Right_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11436__A _06405_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07764_ net1194 team_03_WB.instance_to_wrap.core.register_file.registers_state\[716\]
+ vssd1 vssd1 vccd1 vccd1 _03706_ sky130_fd_sc_hd__or2_1
XFILLER_0_2_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_168_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09503_ net538 _05443_ vssd1 vssd1 vccd1 vccd1 _05445_ sky130_fd_sc_hd__nand2_1
XFILLER_0_116_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08497__B1 net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07695_ net1146 _03632_ _03634_ _03636_ net717 vssd1 vssd1 vccd1 vccd1 _03637_ sky130_fd_sc_hd__a41o_1
XFILLER_0_91_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_155_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout355_A _06818_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11870__S net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1097_A net1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09434_ net546 _04894_ _04955_ vssd1 vssd1 vccd1 vccd1 _05376_ sky130_fd_sc_hd__o21ba_1
XANTENNA__06964__S net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10994__B net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09365_ _05193_ _05305_ vssd1 vssd1 vccd1 vccd1 _05307_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout522_A _06322_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12267__A net1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_228 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1264_A net1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09997__A0 _05882_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10056__B1 net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11171__A net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08316_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[920\] net999
+ _04252_ net1064 vssd1 vssd1 vccd1 vccd1 _04258_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_23_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09296_ _03459_ _05237_ vssd1 vssd1 vccd1 vccd1 _05238_ sky130_fd_sc_hd__xor2_1
XFILLER_0_117_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_43_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_598 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_90_Right_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout310_X net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07472__A1 net1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08247_ net1226 team_03_WB.instance_to_wrap.core.register_file.registers_state\[466\]
+ net950 team_03_WB.instance_to_wrap.core.register_file.registers_state\[498\] net1210
+ vssd1 vssd1 vccd1 vccd1 _04189_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_95_2322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1431_A net1435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07472__B2 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_95_2333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1052_X net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout408_X net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_160_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08178_ net433 net427 _04119_ vssd1 vssd1 vccd1 vccd1 _04120_ sky130_fd_sc_hd__nor3_1
XANTENNA__10359__B2 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11556__B1 net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout891_A net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_3083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_3094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout989_A net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07129_ net1109 team_03_WB.instance_to_wrap.core.register_file.registers_state\[576\]
+ vssd1 vssd1 vccd1 vccd1 _03071_ sky130_fd_sc_hd__and2_1
XFILLER_0_30_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10140_ _03390_ _05980_ vssd1 vssd1 vccd1 vccd1 _05982_ sky130_fd_sc_hd__nand2_1
XANTENNA__08972__A1 net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput170 net170 vssd1 vssd1 vccd1 vccd1 SEL_O[2] sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout777_X net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput181 net181 vssd1 vssd1 vccd1 vccd1 gpio_oeb[16] sky130_fd_sc_hd__buf_2
Xoutput192 net192 vssd1 vssd1 vccd1 vccd1 gpio_oeb[27] sky130_fd_sc_hd__clkbuf_4
X_10071_ team_03_WB.instance_to_wrap.core.i_hit _05914_ vssd1 vssd1 vccd1 vccd1 _05915_
+ sky130_fd_sc_hd__and2_4
XANTENNA__12730__A net1380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11049__C _06527_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout944_X net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13830_ clknet_leaf_73_wb_clk_i _01594_ _00195_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[184\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_98_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13761_ clknet_leaf_179_wb_clk_i _01525_ _00126_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[115\]
+ sky130_fd_sc_hd__dfrtp_1
X_10973_ team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[0\] net314 net309 _05928_
+ vssd1 vssd1 vccd1 vccd1 _06552_ sky130_fd_sc_hd__or4_1
XFILLER_0_134_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_67_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11780__S net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12712_ net1297 vssd1 vssd1 vccd1 vccd1 _00476_ sky130_fd_sc_hd__inv_2
XANTENNA__10834__A2 net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_139_3226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13692_ clknet_leaf_149_wb_clk_i _01456_ _00057_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[46\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_139_3237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_108_wb_clk_i_A clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_128_718 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12643_ net1356 vssd1 vssd1 vccd1 vccd1 _00407_ sky130_fd_sc_hd__inv_2
XFILLER_0_155_526 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10047__B1 net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_156_3573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_156_3584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12574_ net1391 vssd1 vssd1 vccd1 vccd1 _00338_ sky130_fd_sc_hd__inv_2
XANTENNA__07999__C1 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14313_ clknet_leaf_70_wb_clk_i _02077_ _00678_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[667\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11525_ net2300 net482 _06781_ net492 vssd1 vssd1 vccd1 vccd1 _01984_ sky130_fd_sc_hd__a22o_1
XFILLER_0_136_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08660__B1 net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14244_ clknet_leaf_24_wb_clk_i _02008_ _00609_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[598\]
+ sky130_fd_sc_hd__dfrtp_1
X_11456_ net494 net623 _06581_ net392 net2332 vssd1 vssd1 vccd1 vccd1 _02037_ sky130_fd_sc_hd__a32o_1
XANTENNA__08007__A3 net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1099 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10407_ net284 _06231_ net681 vssd1 vssd1 vccd1 vccd1 _06232_ sky130_fd_sc_hd__o21ai_1
X_14175_ clknet_leaf_20_wb_clk_i _01939_ _00540_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[529\]
+ sky130_fd_sc_hd__dfrtp_1
X_11387_ net1249 net839 _06536_ net669 vssd1 vssd1 vccd1 vccd1 _06746_ sky130_fd_sc_hd__and4_1
XFILLER_0_0_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13126_ net1299 vssd1 vssd1 vccd1 vccd1 _00890_ sky130_fd_sc_hd__inv_2
X_10338_ _06150_ _06174_ vssd1 vssd1 vccd1 vccd1 _06175_ sky130_fd_sc_hd__and2b_1
XANTENNA__06974__B1 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_119_wb_clk_i clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_119_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__09933__B net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13057_ net1271 vssd1 vssd1 vccd1 vccd1 _00821_ sky130_fd_sc_hd__inv_2
X_10269_ _06107_ _06109_ _05976_ _05979_ vssd1 vssd1 vccd1 vccd1 _06111_ sky130_fd_sc_hd__a211o_1
XANTENNA__12640__A net1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08176__C1 net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1340 net1341 vssd1 vssd1 vccd1 vccd1 net1340 sky130_fd_sc_hd__buf_4
XANTENNA__08715__A1 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_1016 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12008_ _06758_ net453 net359 net2359 vssd1 vssd1 vccd1 vccd1 _01537_ sky130_fd_sc_hd__a22o_1
Xfanout1351 net1352 vssd1 vssd1 vccd1 vccd1 net1351 sky130_fd_sc_hd__buf_4
Xfanout1362 net1363 vssd1 vssd1 vccd1 vccd1 net1362 sky130_fd_sc_hd__buf_4
Xfanout1373 net1381 vssd1 vssd1 vccd1 vccd1 net1373 sky130_fd_sc_hd__clkbuf_2
XANTENNA_clkbuf_leaf_147_wb_clk_i_A clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout1384 net1393 vssd1 vssd1 vccd1 vccd1 net1384 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_108_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1395 net1396 vssd1 vssd1 vccd1 vccd1 net1395 sky130_fd_sc_hd__buf_4
XANTENNA__10160__A _03679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_2996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13959_ clknet_leaf_111_wb_clk_i _01723_ _00324_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[313\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08479__B1 net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08836__Y _04778_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_10 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07480_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[949\] net770
+ net1014 vssd1 vssd1 vccd1 vccd1 _03422_ sky130_fd_sc_hd__o21a_1
XFILLER_0_159_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10038__B1 net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09979__A0 _03059_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09150_ _05084_ _05086_ _05089_ _05091_ net554 net567 vssd1 vssd1 vccd1 vccd1 _05092_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_90_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_140_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08100__C1 net1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08101_ net1172 team_03_WB.instance_to_wrap.core.register_file.registers_state\[474\]
+ net759 team_03_WB.instance_to_wrap.core.register_file.registers_state\[506\] net1151
+ vssd1 vssd1 vccd1 vccd1 _04043_ sky130_fd_sc_hd__o221a_1
XFILLER_0_71_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07454__A1 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09081_ net1240 team_03_WB.instance_to_wrap.core.register_file.registers_state\[461\]
+ net982 team_03_WB.instance_to_wrap.core.register_file.registers_state\[493\] net1215
+ vssd1 vssd1 vccd1 vccd1 _05023_ sky130_fd_sc_hd__o221a_1
XANTENNA__11250__A2 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_900 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08032_ net1085 team_03_WB.instance_to_wrap.core.register_file.registers_state\[369\]
+ net890 _03973_ net1126 vssd1 vssd1 vccd1 vccd1 _03974_ sky130_fd_sc_hd__o311a_1
Xinput50 gpio_in[25] vssd1 vssd1 vccd1 vccd1 net50 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput61 gpio_in[5] vssd1 vssd1 vccd1 vccd1 net61 sky130_fd_sc_hd__clkbuf_1
Xinput72 wbs_adr_i[14] vssd1 vssd1 vccd1 vccd1 net72 sky130_fd_sc_hd__buf_1
Xhold801 team_03_WB.instance_to_wrap.core.register_file.registers_state\[926\] vssd1
+ vssd1 vccd1 vccd1 net2294 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold812 team_03_WB.instance_to_wrap.core.register_file.registers_state\[630\] vssd1
+ vssd1 vccd1 vccd1 net2305 sky130_fd_sc_hd__dlygate4sd3_1
Xinput83 wbs_adr_i[24] vssd1 vssd1 vccd1 vccd1 net83 sky130_fd_sc_hd__clkbuf_1
Xhold823 team_03_WB.instance_to_wrap.core.register_file.registers_state\[494\] vssd1
+ vssd1 vccd1 vccd1 net2316 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07206__A1 net1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput94 wbs_adr_i[5] vssd1 vssd1 vccd1 vccd1 net94 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__11002__A2 net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold834 team_03_WB.instance_to_wrap.core.register_file.registers_state\[790\] vssd1
+ vssd1 vccd1 vccd1 net2327 sky130_fd_sc_hd__dlygate4sd3_1
Xhold845 team_03_WB.instance_to_wrap.core.register_file.registers_state\[773\] vssd1
+ vssd1 vccd1 vccd1 net2338 sky130_fd_sc_hd__dlygate4sd3_1
Xhold856 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[1\] vssd1 vssd1 vccd1
+ vccd1 net2349 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_2230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08954__A1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[9\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_186_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold867 team_03_WB.instance_to_wrap.core.register_file.registers_state\[374\] vssd1
+ vssd1 vccd1 vccd1 net2360 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold878 team_03_WB.instance_to_wrap.core.register_file.registers_state\[502\] vssd1
+ vssd1 vccd1 vccd1 net2371 sky130_fd_sc_hd__dlygate4sd3_1
X_09983_ _05868_ net1912 net289 vssd1 vssd1 vccd1 vccd1 _02731_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold889 team_03_WB.instance_to_wrap.core.register_file.registers_state\[286\] vssd1
+ vssd1 vccd1 vccd1 net2382 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10761__A1 net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06965__B1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11865__S net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08934_ net1222 _04872_ _04873_ vssd1 vssd1 vccd1 vccd1 _04876_ sky130_fd_sc_hd__nand3_1
XANTENNA__12550__A net1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1012_A net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1097 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08167__C1 net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10989__B net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08865_ net848 _04787_ _04793_ _04806_ vssd1 vssd1 vccd1 vccd1 _04807_ sky130_fd_sc_hd__a31o_4
XANTENNA_fanout472_A net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07914__C1 net1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07816_ net1189 _02814_ _02924_ net1252 _03757_ vssd1 vssd1 vccd1 vccd1 _03758_ sky130_fd_sc_hd__a221oi_4
X_08796_ _04730_ _04731_ _04737_ _04734_ net1066 net1081 vssd1 vssd1 vccd1 vccd1 _04738_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_88_2181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_2192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08178__C _04119_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07747_ net1098 team_03_WB.instance_to_wrap.core.register_file.registers_state\[236\]
+ net898 vssd1 vssd1 vccd1 vccd1 _03689_ sky130_fd_sc_hd__or3_1
XPHY_EDGE_ROW_154_Right_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1381_A net1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout737_A net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout358_X net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_64_Left_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_487 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08475__A net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_342 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07678_ _03618_ _03619_ net820 vssd1 vssd1 vccd1 vccd1 _03620_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_0_Right_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09417_ net553 _05357_ _05358_ net568 vssd1 vssd1 vccd1 vccd1 _05359_ sky130_fd_sc_hd__o211a_1
XANTENNA__12018__A1 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_149_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout525_X net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11105__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1267_X net1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09348_ _05288_ _05289_ vssd1 vssd1 vccd1 vccd1 _05290_ sky130_fd_sc_hd__and2_1
XANTENNA__11332__C net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_134_3123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_902 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10229__B net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_134_3134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09279_ _04893_ _05219_ vssd1 vssd1 vccd1 vccd1 _05221_ sky130_fd_sc_hd__xor2_1
XFILLER_0_117_283 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_946 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08922__B net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11310_ _06620_ net2436 net405 vssd1 vssd1 vccd1 vccd1 _02135_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_151_3470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12290_ net1296 vssd1 vssd1 vccd1 vccd1 _00054_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_151_3481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout894_X net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14713__Q team_03_WB.instance_to_wrap.core.decoder.inst\[10\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11241_ net1247 net836 net279 net670 vssd1 vssd1 vccd1 vccd1 _06688_ sky130_fd_sc_hd__and4_1
XPHY_EDGE_ROW_73_Left_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11172_ net2267 net412 _06665_ net495 vssd1 vssd1 vccd1 vccd1 _02221_ sky130_fd_sc_hd__a22o_1
XFILLER_0_30_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06956__B1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10123_ _05964_ vssd1 vssd1 vccd1 vccd1 _05965_ sky130_fd_sc_hd__inv_2
XFILLER_0_98_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14931_ clknet_leaf_43_wb_clk_i _02686_ _01296_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_O\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_10054_ net33 net1036 net909 net2777 vssd1 vssd1 vccd1 vccd1 _02677_ sky130_fd_sc_hd__o22a_1
XANTENNA_input33_A DAT_I[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10504__A1 net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11701__B1 net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11076__A net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14862_ clknet_leaf_59_wb_clk_i net1629 _01227_ vssd1 vssd1 vccd1 vccd1 net118 sky130_fd_sc_hd__dfrtp_1
XANTENNA__09502__A1_N team_03_WB.instance_to_wrap.core.decoder.inst\[27\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07381__B1 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13813_ clknet_leaf_127_wb_clk_i _01577_ _00178_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[167\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_106_2546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_82_Left_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14793_ clknet_leaf_92_wb_clk_i _02557_ _01158_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_I\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_240 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_121_Right_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_158_3613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_158_3624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13744_ clknet_leaf_157_wb_clk_i _01508_ _00109_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[98\]
+ sky130_fd_sc_hd__dfrtp_1
X_10956_ team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[3\] net306 vssd1 vssd1
+ vccd1 vccd1 _06538_ sky130_fd_sc_hd__and2_1
XFILLER_0_58_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_123_2893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07133__B1 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_156_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13675_ clknet_leaf_42_wb_clk_i _01439_ _00040_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11480__A2 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10887_ net688 _05811_ vssd1 vssd1 vccd1 vccd1 _06482_ sky130_fd_sc_hd__nand2_1
XFILLER_0_128_548 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12626_ net1395 vssd1 vssd1 vccd1 vccd1 _00390_ sky130_fd_sc_hd__inv_2
XFILLER_0_155_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08859__S1 net1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11768__B1 net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08633__B1 net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12557_ net1311 vssd1 vssd1 vccd1 vccd1 _00321_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_171_3879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11508_ _06626_ net2746 net390 vssd1 vssd1 vccd1 vccd1 _01998_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_696 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_91_Left_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_151_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_34 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12488_ net1290 vssd1 vssd1 vccd1 vccd1 _00252_ sky130_fd_sc_hd__inv_2
Xhold108 _02574_ vssd1 vssd1 vccd1 vccd1 net1601 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_151_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold119 team_03_WB.instance_to_wrap.ADR_I\[8\] vssd1 vssd1 vccd1 vccd1 net1612 sky130_fd_sc_hd__dlygate4sd3_1
X_14227_ clknet_leaf_99_wb_clk_i _01991_ _00592_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[581\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_151_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11439_ net2676 net392 _06759_ net492 vssd1 vssd1 vccd1 vccd1 _02048_ sky130_fd_sc_hd__a22o_1
XFILLER_0_46_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08936__A1 net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07295__S0 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14158_ clknet_leaf_128_wb_clk_i _01922_ _00523_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[512\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13109_ net1275 vssd1 vssd1 vccd1 vccd1 _00873_ sky130_fd_sc_hd__inv_2
X_06980_ net615 _02893_ vssd1 vssd1 vccd1 vccd1 _02922_ sky130_fd_sc_hd__nor2_1
X_14089_ clknet_leaf_75_wb_clk_i _01853_ _00454_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[443\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_28_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07464__A net1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1170 net1171 vssd1 vssd1 vccd1 vccd1 net1170 sky130_fd_sc_hd__clkbuf_4
X_08650_ _04591_ vssd1 vssd1 vccd1 vccd1 _04592_ sky130_fd_sc_hd__inv_2
XANTENNA__07183__B net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1181 net1183 vssd1 vssd1 vccd1 vccd1 net1181 sky130_fd_sc_hd__buf_2
XANTENNA__07372__A0 _03312_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1192 net1193 vssd1 vssd1 vccd1 vccd1 net1192 sky130_fd_sc_hd__clkbuf_2
X_07601_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[441\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[409\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[313\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[281\]
+ net788 net1137 vssd1 vssd1 vccd1 vccd1 _03543_ sky130_fd_sc_hd__mux4_1
XFILLER_0_117_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08581_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[573\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[541\]
+ net967 vssd1 vssd1 vccd1 vccd1 _04523_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_87_wb_clk_i clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_87_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__11136__D net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07532_ net1198 team_03_WB.instance_to_wrap.core.register_file.registers_state\[134\]
+ vssd1 vssd1 vccd1 vccd1 _03474_ sky130_fd_sc_hd__or2_1
XFILLER_0_48_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_1143 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_16_wb_clk_i clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_16_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__09664__A2 _04207_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07463_ net1163 _03404_ vssd1 vssd1 vccd1 vccd1 _03405_ sky130_fd_sc_hd__or2_1
XANTENNA__08872__B1 net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09202_ net583 net579 net572 _05124_ vssd1 vssd1 vccd1 vccd1 _05144_ sky130_fd_sc_hd__and4_2
XANTENNA__11152__C net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_524 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07394_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[575\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[543\]
+ net763 vssd1 vssd1 vccd1 vccd1 _03336_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_40_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11759__B1 net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09133_ _02804_ _02944_ net594 vssd1 vssd1 vccd1 vccd1 _05075_ sky130_fd_sc_hd__and3_1
XFILLER_0_115_710 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_173_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_161_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout318_A _05927_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10991__C _06414_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07522__S1 net1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09064_ net1047 team_03_WB.instance_to_wrap.core.register_file.registers_state\[847\]
+ net998 team_03_WB.instance_to_wrap.core.register_file.registers_state\[879\] net949
+ vssd1 vssd1 vccd1 vccd1 _05006_ sky130_fd_sc_hd__a221o_1
XFILLER_0_142_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_163_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08015_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[561\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[529\]
+ net765 vssd1 vssd1 vccd1 vccd1 _03957_ sky130_fd_sc_hd__mux2_1
XANTENNA__10065__A team_03_WB.instance_to_wrap.core.decoder.inst\[24\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold620 team_03_WB.instance_to_wrap.core.register_file.registers_state\[182\] vssd1
+ vssd1 vccd1 vccd1 net2113 sky130_fd_sc_hd__dlygate4sd3_1
Xhold631 team_03_WB.instance_to_wrap.core.register_file.registers_state\[775\] vssd1
+ vssd1 vccd1 vccd1 net2124 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap350 _04863_ vssd1 vssd1 vccd1 vccd1 net350 sky130_fd_sc_hd__buf_1
Xhold642 team_03_WB.instance_to_wrap.core.register_file.registers_state\[115\] vssd1
+ vssd1 vccd1 vccd1 net2135 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1227_A net1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08927__A1 net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold653 team_03_WB.instance_to_wrap.core.register_file.registers_state\[768\] vssd1
+ vssd1 vccd1 vccd1 net2146 sky130_fd_sc_hd__dlygate4sd3_1
Xhold664 team_03_WB.instance_to_wrap.core.register_file.registers_state\[545\] vssd1
+ vssd1 vccd1 vccd1 net2157 sky130_fd_sc_hd__dlygate4sd3_1
Xhold675 team_03_WB.instance_to_wrap.core.register_file.registers_state\[435\] vssd1
+ vssd1 vccd1 vccd1 net2168 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11931__A0 _06628_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11595__S net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold686 team_03_WB.instance_to_wrap.core.register_file.registers_state\[295\] vssd1
+ vssd1 vccd1 vccd1 net2179 sky130_fd_sc_hd__dlygate4sd3_1
Xhold697 team_03_WB.instance_to_wrap.core.register_file.registers_state\[268\] vssd1
+ vssd1 vccd1 vccd1 net2190 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07060__C1 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09966_ _05887_ net2660 net292 vssd1 vssd1 vccd1 vccd1 _02744_ sky130_fd_sc_hd__mux2_1
XANTENNA__07374__A net1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08917_ _04855_ _04856_ _04858_ _04857_ net942 net862 vssd1 vssd1 vccd1 vccd1 _04859_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__11608__B net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09897_ net321 _05419_ _05838_ vssd1 vssd1 vccd1 vccd1 _05839_ sky130_fd_sc_hd__a21bo_1
XANTENNA_fanout854_A net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout475_X net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10498__B1 net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10004__S net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08848_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[416\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[384\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[288\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[256\]
+ net990 net1078 vssd1 vssd1 vccd1 vccd1 _04790_ sky130_fd_sc_hd__mux4_1
XANTENNA__07363__B1 net1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08779_ net1050 team_03_WB.instance_to_wrap.core.register_file.registers_state\[322\]
+ net1002 team_03_WB.instance_to_wrap.core.register_file.registers_state\[354\] net1214
+ vssd1 vssd1 vccd1 vccd1 _04721_ sky130_fd_sc_hd__a221o_1
XFILLER_0_68_903 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout642_X net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10810_ net691 _05583_ net585 vssd1 vssd1 vccd1 vccd1 _06417_ sky130_fd_sc_hd__o21ai_2
XTAP_TAPCELL_ROW_0_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_711 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08409__S net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11790_ net2722 _06621_ net327 vssd1 vssd1 vccd1 vccd1 _01748_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_0_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07115__B1 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09655__A2 _05281_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11998__B1 net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08312__C1 net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10741_ net1673 net529 net524 _06362_ vssd1 vssd1 vccd1 vccd1 _02445_ sky130_fd_sc_hd__a22o_1
XANTENNA__07666__A1 net1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11343__B net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_2443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11462__A2 net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_2454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout907_X net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_939 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07130__A3 net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13460_ net1323 vssd1 vssd1 vccd1 vccd1 _01224_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_153_3510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10672_ _05429_ _06313_ vssd1 vssd1 vccd1 vccd1 _06314_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_153_3521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08933__A net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07418__A1 net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12411_ net1362 vssd1 vssd1 vccd1 vccd1 _00175_ sky130_fd_sc_hd__inv_2
XANTENNA__11214__A2 net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08615__B1 net1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13391_ net1416 vssd1 vssd1 vccd1 vccd1 _01155_ sky130_fd_sc_hd__inv_2
XFILLER_0_164_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09812__C1 _04777_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12455__A net1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07549__A _03459_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_527 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12342_ net1258 vssd1 vssd1 vccd1 vccd1 _00106_ sky130_fd_sc_hd__inv_2
XANTENNA__11765__A3 net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15061_ net1447 vssd1 vssd1 vccd1 vccd1 irq[0] sky130_fd_sc_hd__buf_2
X_12273_ net1265 vssd1 vssd1 vccd1 vccd1 _00037_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_79_1991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08918__A1 net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14012_ clknet_leaf_146_wb_clk_i _01776_ _00377_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[366\]
+ sky130_fd_sc_hd__dfrtp_1
X_11224_ _06456_ _06517_ vssd1 vssd1 vccd1 vccd1 _06683_ sky130_fd_sc_hd__nor2_1
XANTENNA__10725__A1 net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11155_ net630 _06654_ vssd1 vssd1 vccd1 vccd1 _06655_ sky130_fd_sc_hd__nor2_1
X_10106_ _02834_ _05916_ vssd1 vssd1 vccd1 vccd1 _05950_ sky130_fd_sc_hd__or2_4
X_11086_ _06454_ net2429 net416 vssd1 vssd1 vccd1 vccd1 _02262_ sky130_fd_sc_hd__mux2_1
XANTENNA__07715__C net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10489__B1 net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10037_ net20 net1040 net911 net2765 vssd1 vssd1 vccd1 vccd1 _02694_ sky130_fd_sc_hd__a22o_1
X_14914_ clknet_leaf_43_wb_clk_i _02669_ _01279_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_O\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__11237__C net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_125_2933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07354__B1 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09894__A2 _04323_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08551__C1 net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14845_ clknet_leaf_85_wb_clk_i _02609_ _01210_ vssd1 vssd1 vccd1 vccd1 net131 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_172_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1138 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_16 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11093__X _06623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08529__S0 net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11534__A net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14776_ clknet_leaf_89_wb_clk_i _02540_ _01141_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_I\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_105_23 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11988_ net273 net2517 net443 vssd1 vssd1 vccd1 vccd1 _01556_ sky130_fd_sc_hd__mux2_1
XFILLER_0_147_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11989__B1 net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07657__A1 net1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13727_ clknet_leaf_19_wb_clk_i _01491_ _00092_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[81\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11253__B net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10939_ team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[6\] net306 vssd1 vssd1
+ vccd1 vccd1 _06524_ sky130_fd_sc_hd__and2_1
XANTENNA__08854__B1 net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11453__A2 net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_173_3919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09939__A _03526_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13658_ clknet_leaf_141_wb_clk_i _01422_ _00023_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_171_602 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12609_ net1262 vssd1 vssd1 vccd1 vccd1 _00373_ sky130_fd_sc_hd__inv_2
XFILLER_0_144_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13589_ net1343 vssd1 vssd1 vccd1 vccd1 _01353_ sky130_fd_sc_hd__inv_2
XFILLER_0_143_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10413__B1 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11756__A3 net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10964__A1 _06542_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_134_wb_clk_i clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_134_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_121_99 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08909__A1 net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09031__B1 net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09820_ net565 _05134_ vssd1 vssd1 vccd1 vccd1 _05762_ sky130_fd_sc_hd__or2_1
Xfanout407 _06717_ vssd1 vssd1 vccd1 vccd1 net407 sky130_fd_sc_hd__buf_4
Xfanout418 _06610_ vssd1 vssd1 vccd1 vccd1 net418 sky130_fd_sc_hd__buf_8
Xfanout429 net430 vssd1 vssd1 vccd1 vccd1 net429 sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_129_Left_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07593__B1 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09751_ _04816_ _05692_ net666 vssd1 vssd1 vccd1 vccd1 _05693_ sky130_fd_sc_hd__o21a_1
X_06963_ net1121 _02903_ _02904_ vssd1 vssd1 vccd1 vccd1 _02905_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_33_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08702_ net1222 _04642_ _04643_ vssd1 vssd1 vccd1 vccd1 _04644_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_33_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09682_ _05296_ _05298_ _05597_ vssd1 vssd1 vccd1 vccd1 _05624_ sky130_fd_sc_hd__nand3_1
X_06894_ _02823_ _02831_ vssd1 vssd1 vccd1 vccd1 _02836_ sky130_fd_sc_hd__or2_1
XFILLER_0_154_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08542__C1 net1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08633_ net1053 team_03_WB.instance_to_wrap.core.register_file.registers_state\[454\]
+ net1006 team_03_WB.instance_to_wrap.core.register_file.registers_state\[486\] net1077
+ vssd1 vssd1 vccd1 vccd1 _04575_ sky130_fd_sc_hd__a221o_1
XANTENNA__11692__A2 net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout268_A _06541_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08564_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[61\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[29\]
+ net966 vssd1 vssd1 vccd1 vccd1 _04506_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_2037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_2048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07515_ net823 _03456_ net724 vssd1 vssd1 vccd1 vccd1 _03457_ sky130_fd_sc_hd__a21o_1
XANTENNA__10247__A3 _06086_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08495_ net864 _04433_ _04436_ vssd1 vssd1 vccd1 vccd1 _04437_ sky130_fd_sc_hd__o21ai_1
XANTENNA__08845__B1 net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11444__A2 net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout435_A net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_138_Left_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10652__A0 net1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1177_A net1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07446_ _03386_ _03387_ net817 vssd1 vssd1 vccd1 vccd1 _03388_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_88_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_378 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold1285_A team_03_WB.instance_to_wrap.CPU_DAT_O\[16\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout602_A net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07377_ net741 _03315_ _03316_ _03317_ _03318_ vssd1 vssd1 vccd1 vccd1 _03319_ sky130_fd_sc_hd__o32a_1
XFILLER_0_91_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_146_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1344_A net1346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09116_ net1051 team_03_WB.instance_to_wrap.core.register_file.registers_state\[846\]
+ net1001 team_03_WB.instance_to_wrap.core.register_file.registers_state\[878\] net1214
+ vssd1 vssd1 vccd1 vccd1 _05058_ sky130_fd_sc_hd__a221o_1
XFILLER_0_150_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11747__A3 net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08073__A1 net1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_871 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10955__A1 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_584 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07281__C1 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09047_ _04987_ _04988_ net855 vssd1 vssd1 vccd1 vccd1 _04989_ sky130_fd_sc_hd__o21a_1
XFILLER_0_128_1070 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1132_X net1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07259__S0 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold450 team_03_WB.instance_to_wrap.core.register_file.registers_state\[300\] vssd1
+ vssd1 vccd1 vccd1 net1943 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold461 team_03_WB.instance_to_wrap.core.register_file.registers_state\[703\] vssd1
+ vssd1 vccd1 vccd1 net1954 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout971_A net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold472 net177 vssd1 vssd1 vccd1 vccd1 net1965 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1042 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11904__B1 net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_147_Left_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09573__A1 net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_3022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold483 team_03_WB.instance_to_wrap.core.register_file.registers_state\[247\] vssd1
+ vssd1 vccd1 vccd1 net1976 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_3033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold494 team_03_WB.instance_to_wrap.core.register_file.registers_state\[446\] vssd1
+ vssd1 vccd1 vccd1 net1987 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11380__A1 net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout930 net932 vssd1 vssd1 vccd1 vccd1 net930 sky130_fd_sc_hd__buf_4
Xfanout941 net942 vssd1 vssd1 vccd1 vccd1 net941 sky130_fd_sc_hd__buf_4
XANTENNA__06926__A3 net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09949_ _03136_ net661 vssd1 vssd1 vccd1 vccd1 _05879_ sky130_fd_sc_hd__nor2_2
Xfanout952 net956 vssd1 vssd1 vccd1 vccd1 net952 sky130_fd_sc_hd__clkbuf_4
Xfanout963 net964 vssd1 vssd1 vccd1 vccd1 net963 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout857_X net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08128__A2 net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_146_3380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout974 _04086_ vssd1 vssd1 vccd1 vccd1 net974 sky130_fd_sc_hd__clkbuf_4
Xfanout985 net988 vssd1 vssd1 vccd1 vccd1 net985 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_5_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout996 net997 vssd1 vssd1 vccd1 vccd1 net996 sky130_fd_sc_hd__clkbuf_2
X_12960_ net1399 vssd1 vssd1 vccd1 vccd1 _00724_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_5_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11057__C _06545_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1150 team_03_WB.instance_to_wrap.core.register_file.registers_state\[659\] vssd1
+ vssd1 vccd1 vccd1 net2643 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08928__A net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09523__S net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1161 team_03_WB.instance_to_wrap.core.register_file.registers_state\[83\] vssd1
+ vssd1 vccd1 vccd1 net2654 sky130_fd_sc_hd__dlygate4sd3_1
X_11911_ _06612_ net2685 net367 vssd1 vssd1 vccd1 vccd1 _01631_ sky130_fd_sc_hd__mux2_1
Xhold1172 team_03_WB.instance_to_wrap.core.register_file.registers_state\[600\] vssd1
+ vssd1 vccd1 vccd1 net2665 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_142_3288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11683__A2 net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1183 team_03_WB.instance_to_wrap.core.register_file.registers_state\[638\] vssd1
+ vssd1 vccd1 vccd1 net2676 sky130_fd_sc_hd__dlygate4sd3_1
X_12891_ net1361 vssd1 vssd1 vccd1 vccd1 _00655_ sky130_fd_sc_hd__inv_2
XFILLER_0_169_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_142_3299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1194 team_03_WB.instance_to_wrap.core.register_file.registers_state\[191\] vssd1
+ vssd1 vccd1 vccd1 net2687 sky130_fd_sc_hd__dlygate4sd3_1
X_14630_ clknet_leaf_70_wb_clk_i _02394_ _00995_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[984\]
+ sky130_fd_sc_hd__dfstp_1
X_11842_ _06455_ net461 vssd1 vssd1 vccd1 vccd1 _06812_ sky130_fd_sc_hd__nand2_4
XTAP_TAPCELL_ROW_16_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09089__B1 net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_156_Left_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_120_2830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_2841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_610 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14561_ clknet_leaf_179_wb_clk_i _02325_ _00926_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[915\]
+ sky130_fd_sc_hd__dfrtp_1
X_11773_ net653 _06606_ net467 net333 net1956 vssd1 vssd1 vccd1 vccd1 _01764_ sky130_fd_sc_hd__a32o_1
XFILLER_0_138_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10643__A0 net1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13512_ net1321 vssd1 vssd1 vccd1 vccd1 _01276_ sky130_fd_sc_hd__inv_2
X_10724_ _05833_ net602 vssd1 vssd1 vccd1 vccd1 _06354_ sky130_fd_sc_hd__nand2_1
XFILLER_0_166_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14492_ clknet_leaf_149_wb_clk_i _02256_ _00857_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[846\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08663__A net1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13443_ net1423 vssd1 vssd1 vccd1 vccd1 _01207_ sky130_fd_sc_hd__inv_2
XFILLER_0_137_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_153_635 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10655_ team_03_WB.instance_to_wrap.core.control_logic.instruction\[6\] team_03_WB.instance_to_wrap.CPU_DAT_O\[6\]
+ net846 vssd1 vssd1 vccd1 vccd1 _02473_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11738__A3 net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08064__A1 net1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload17 clknet_leaf_5_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload17/Y sky130_fd_sc_hd__clkinv_4
X_13374_ net1415 vssd1 vssd1 vccd1 vccd1 _01138_ sky130_fd_sc_hd__inv_2
Xclkload28 clknet_leaf_173_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload28/Y sky130_fd_sc_hd__clkinv_4
X_10586_ net1666 net534 net601 _03023_ vssd1 vssd1 vccd1 vccd1 _02537_ sky130_fd_sc_hd__a22o_1
XANTENNA__10946__A1 team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[5\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15113_ net913 vssd1 vssd1 vccd1 vccd1 net246 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_118_2792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload39 clknet_leaf_185_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload39/Y sky130_fd_sc_hd__clkinv_2
XFILLER_0_152_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12325_ net1353 vssd1 vssd1 vccd1 vccd1 _00089_ sky130_fd_sc_hd__inv_2
XANTENNA__07811__A1 net1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_688 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_165_Left_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15044_ clknet_leaf_90_wb_clk_i _02764_ _01409_ vssd1 vssd1 vccd1 vccd1 net200 sky130_fd_sc_hd__dfrtp_1
X_12256_ net1430 vssd1 vssd1 vccd1 vccd1 _00020_ sky130_fd_sc_hd__inv_2
XANTENNA__06911__A net1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11529__A net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11207_ _06438_ net2163 net487 vssd1 vssd1 vccd1 vccd1 _02201_ sky130_fd_sc_hd__mux2_1
XANTENNA__10433__A net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12187_ net1537 vssd1 vssd1 vccd1 vccd1 _02366_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_166_3778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_166_3789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11138_ net276 net651 net708 net696 vssd1 vssd1 vccd1 vccd1 _06645_ sky130_fd_sc_hd__and4_1
XANTENNA__09941__B net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11069_ _06612_ net2647 net417 vssd1 vssd1 vccd1 vccd1 _02271_ sky130_fd_sc_hd__mux2_1
XANTENNA__07327__B1 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11123__B2 net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08524__C1 net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07742__A net1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07878__A1 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14828_ clknet_leaf_94_wb_clk_i net1671 _01193_ vssd1 vssd1 vccd1 vccd1 net149 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08827__B1 net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14759_ clknet_leaf_48_wb_clk_i _02523_ _01124_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_47_939 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07300_ team_03_WB.instance_to_wrap.core.decoder.inst\[29\] net826 vssd1 vssd1 vccd1
+ vccd1 _03242_ sky130_fd_sc_hd__nand2_2
XANTENNA__10634__A0 team_03_WB.instance_to_wrap.core.decoder.inst\[27\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08280_ net1063 _04218_ _04219_ _04221_ vssd1 vssd1 vccd1 vccd1 _04222_ sky130_fd_sc_hd__o31a_1
XFILLER_0_117_816 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_630 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07231_ net1191 net881 team_03_WB.instance_to_wrap.core.register_file.registers_state\[776\]
+ vssd1 vssd1 vccd1 vccd1 _03173_ sky130_fd_sc_hd__a21o_1
XFILLER_0_128_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_144_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11203__S net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07162_ _03075_ _03081_ _03102_ net612 vssd1 vssd1 vccd1 vccd1 _03104_ sky130_fd_sc_hd__a211o_2
XANTENNA__08055__A1 net1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07093_ _03032_ _03034_ net748 vssd1 vssd1 vccd1 vccd1 _03035_ sky130_fd_sc_hd__mux2_1
XANTENNA__09608__S net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09004__B1 net995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09555__A1 _04778_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_35_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11362__A1 net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07566__B1 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09803_ net322 _05403_ _05737_ _05740_ _05744_ vssd1 vssd1 vccd1 vccd1 _05745_ sky130_fd_sc_hd__a221o_1
XFILLER_0_10_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11901__A3 net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07995_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[560\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[528\]
+ net782 vssd1 vssd1 vccd1 vccd1 _03937_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout385_A net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11873__S net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09734_ net582 _05663_ _05664_ _05675_ vssd1 vssd1 vccd1 vccd1 _05676_ sky130_fd_sc_hd__a31o_2
X_06946_ _02862_ _02876_ _02887_ net719 vssd1 vssd1 vccd1 vccd1 _02888_ sky130_fd_sc_hd__o22a_4
Xclkbuf_leaf_31_wb_clk_i clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_31_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_2_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09665_ _02804_ _03139_ net535 _05604_ _05606_ vssd1 vssd1 vccd1 vccd1 _05607_ sky130_fd_sc_hd__o221ai_4
XANTENNA_fanout552_A _03105_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06877_ _02808_ _02818_ vssd1 vssd1 vccd1 vccd1 _02819_ sky130_fd_sc_hd__or2_2
XANTENNA_fanout1294_A net1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08616_ net865 _04556_ _04557_ _04555_ vssd1 vssd1 vccd1 vccd1 _04558_ sky130_fd_sc_hd__a31o_1
XFILLER_0_167_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09596_ _04778_ _05527_ _05531_ _05537_ vssd1 vssd1 vccd1 vccd1 _05538_ sky130_fd_sc_hd__o211a_1
XFILLER_0_139_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08547_ net917 _04487_ _04488_ net1218 vssd1 vssd1 vccd1 vccd1 _04489_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout340_X net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1082_X net1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout817_A net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08478_ net944 _04418_ _04419_ net856 vssd1 vssd1 vccd1 vccd1 _04420_ sky130_fd_sc_hd__o211a_1
XANTENNA__12090__A2 net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_706 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07429_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[788\] net795
+ net1041 _03370_ vssd1 vssd1 vccd1 vccd1 _03371_ sky130_fd_sc_hd__o211a_1
XFILLER_0_46_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout605_X net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1347_X net1347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_163_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10440_ team_03_WB.instance_to_wrap.core.pc.current_pc\[8\] net682 _06256_ _06258_
+ vssd1 vssd1 vccd1 vccd1 _02642_ sky130_fd_sc_hd__o22a_1
XFILLER_0_116_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_98_2386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10928__A1 net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_2397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10371_ _05983_ _05986_ _06088_ vssd1 vssd1 vccd1 vccd1 _06202_ sky130_fd_sc_hd__or3_1
XFILLER_0_131_852 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12110_ net1143 _06305_ _06821_ net844 vssd1 vssd1 vccd1 vccd1 _00000_ sky130_fd_sc_hd__a211o_1
XANTENNA__07827__A net1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13090_ net1287 vssd1 vssd1 vccd1 vccd1 _00854_ sky130_fd_sc_hd__inv_2
XFILLER_0_131_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout974_X net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_148_3420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09546__A1 net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12041_ _06609_ net2583 net355 vssd1 vssd1 vccd1 vccd1 _01505_ sky130_fd_sc_hd__mux2_1
XANTENNA__11349__A net1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold280 team_03_WB.instance_to_wrap.CPU_DAT_I\[14\] vssd1 vssd1 vccd1 vccd1 net1773
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold291 team_03_WB.instance_to_wrap.core.ru.state\[4\] vssd1 vssd1 vccd1 vccd1 net1784
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_1847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10156__A2 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_1858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07021__A2 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11068__B _06414_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_144_3328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_3339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout760 net761 vssd1 vssd1 vccd1 vccd1 net760 sky130_fd_sc_hd__buf_4
XANTENNA__11783__S net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout771 net773 vssd1 vssd1 vccd1 vccd1 net771 sky130_fd_sc_hd__clkbuf_4
Xfanout782 net790 vssd1 vssd1 vccd1 vccd1 net782 sky130_fd_sc_hd__clkbuf_2
X_13992_ clknet_leaf_8_wb_clk_i _01756_ _00357_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[346\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout793 net794 vssd1 vssd1 vccd1 vccd1 net793 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_161_3675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_14_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__07562__A net1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_161_3686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12943_ net1394 vssd1 vssd1 vccd1 vccd1 _00707_ sky130_fd_sc_hd__inv_2
XANTENNA__11084__A net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12874_ net1284 vssd1 vssd1 vccd1 vccd1 _00638_ sky130_fd_sc_hd__inv_2
XFILLER_0_73_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11825_ net656 _06656_ net474 net326 net2028 vssd1 vssd1 vccd1 vccd1 _01714_ sky130_fd_sc_hd__a32o_1
X_14613_ clknet_leaf_106_wb_clk_i _02377_ _00978_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[967\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_157_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11234__D net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14544_ clknet_leaf_161_wb_clk_i _02308_ _00909_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[898\]
+ sky130_fd_sc_hd__dfrtp_1
X_11756_ net648 _06581_ net454 net331 net2230 vssd1 vssd1 vccd1 vccd1 _01781_ sky130_fd_sc_hd__a32o_1
XFILLER_0_95_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09482__B1 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12081__A2 net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06906__A net1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10707_ net1677 net528 net523 _06343_ vssd1 vssd1 vccd1 vccd1 _02460_ sky130_fd_sc_hd__a22o_1
X_14475_ clknet_leaf_46_wb_clk_i _02239_ _00840_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[829\]
+ sky130_fd_sc_hd__dfrtp_1
X_11687_ _06729_ net382 net339 net1906 vssd1 vssd1 vccd1 vccd1 _01847_ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13426_ net1433 vssd1 vssd1 vccd1 vccd1 _01190_ sky130_fd_sc_hd__inv_2
XANTENNA__09776__X _05718_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10638_ net1147 net1961 net844 vssd1 vssd1 vccd1 vccd1 _02490_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload106 clknet_leaf_154_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload106/Y sky130_fd_sc_hd__clkinv_1
XFILLER_0_153_487 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10919__A1 team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[10\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload117 clknet_leaf_161_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload117/Y sky130_fd_sc_hd__clkinv_4
Xclkload128 clknet_leaf_141_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload128/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_52_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09785__A1 _03459_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkload139 clknet_leaf_134_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload139/Y sky130_fd_sc_hd__clkinv_2
X_13357_ net1318 vssd1 vssd1 vccd1 vccd1 _01121_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10569_ net1656 net534 net601 _05879_ vssd1 vssd1 vccd1 vccd1 _02554_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_168_3818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10395__A2 net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_168_3829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12308_ net1313 vssd1 vssd1 vccd1 vccd1 _00072_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13288_ net1341 vssd1 vssd1 vccd1 vccd1 _01052_ sky130_fd_sc_hd__inv_2
XFILLER_0_122_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09537__A1 net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11259__A net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15027_ clknet_leaf_103_wb_clk_i _02747_ _01392_ vssd1 vssd1 vccd1 vccd1 net183 sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_53_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_12239_ net1553 vssd1 vssd1 vccd1 vccd1 _01418_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11344__A1 net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07780_ _03715_ _03721_ net718 vssd1 vssd1 vccd1 vccd1 _03722_ sky130_fd_sc_hd__a21o_1
Xinput4 DAT_I[11] vssd1 vssd1 vccd1 vccd1 net4 sky130_fd_sc_hd__buf_1
XFILLER_0_36_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09450_ _05116_ _05118_ vssd1 vssd1 vccd1 vccd1 _05392_ sky130_fd_sc_hd__nor2_1
XFILLER_0_8_1120 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07720__B1 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08401_ _04341_ _04342_ net1223 vssd1 vssd1 vccd1 vccd1 _04343_ sky130_fd_sc_hd__o21a_1
X_09381_ _04354_ _05322_ vssd1 vssd1 vccd1 vccd1 _05323_ sky130_fd_sc_hd__nor2_1
XFILLER_0_164_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08332_ _04270_ _04271_ _04272_ _04273_ net861 net920 vssd1 vssd1 vccd1 vccd1 _04274_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__08276__A1 net1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08507__S net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_157_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10083__A1 _02954_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08263_ net871 _04196_ _04199_ vssd1 vssd1 vccd1 vccd1 _04205_ sky130_fd_sc_hd__or3_1
XFILLER_0_62_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11280__B1 net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07214_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[562\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[530\]
+ net756 vssd1 vssd1 vccd1 vccd1 _03156_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_171_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_92_wb_clk_i_A clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__08590__X _04532_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08194_ net1231 team_03_WB.instance_to_wrap.core.register_file.registers_state\[723\]
+ net957 team_03_WB.instance_to_wrap.core.register_file.registers_state\[755\] net935
+ vssd1 vssd1 vccd1 vccd1 _04136_ sky130_fd_sc_hd__o221a_1
XFILLER_0_6_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11868__S net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07236__C1 net1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_398 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07145_ net1103 team_03_WB.instance_to_wrap.core.register_file.registers_state\[64\]
+ vssd1 vssd1 vccd1 vccd1 _03087_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout300_A _06442_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1042_A net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07787__B1 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08984__C1 net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07076_ net1191 team_03_WB.instance_to_wrap.core.register_file.registers_state\[482\]
+ net882 _03017_ vssd1 vssd1 vccd1 vccd1 _03018_ sky130_fd_sc_hd__a31o_1
XFILLER_0_140_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_93_2283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_2294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1307_A net1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07539__B1 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08736__C1 net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09862__A _05278_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout290_X net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout767_A net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout388_X net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07978_ net1106 team_03_WB.instance_to_wrap.core.register_file.registers_state\[432\]
+ net901 vssd1 vssd1 vccd1 vccd1 _03920_ sky130_fd_sc_hd__or3_1
XFILLER_0_96_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09073__S net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09717_ _05648_ _05649_ _05657_ _05658_ vssd1 vssd1 vccd1 vccd1 _05659_ sky130_fd_sc_hd__o211ai_4
X_06929_ net1154 net1164 vssd1 vssd1 vccd1 vccd1 _02871_ sky130_fd_sc_hd__nor2_4
XANTENNA__11638__A2 net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout934_A net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11108__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09648_ net539 _05588_ vssd1 vssd1 vccd1 vccd1 _05590_ sky130_fd_sc_hd__nand2_1
XANTENNA__07937__S1 net1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11335__C net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07711__B1 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09579_ _05520_ vssd1 vssd1 vccd1 vccd1 _05521_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout722_X net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12728__A net1380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11610_ net1042 net702 _06803_ vssd1 vssd1 vccd1 vccd1 _06804_ sky130_fd_sc_hd__or3_4
XFILLER_0_136_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12590_ net1303 vssd1 vssd1 vccd1 vccd1 _00354_ sky130_fd_sc_hd__inv_2
XFILLER_0_93_864 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14716__Q team_03_WB.instance_to_wrap.core.decoder.inst\[13\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07475__C1 net1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11541_ net493 net622 _06651_ net482 net1982 vssd1 vssd1 vccd1 vccd1 _01974_ sky130_fd_sc_hd__a32o_1
XANTENNA__11351__B net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11810__A2 net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_137_3187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_137_3198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14260_ clknet_leaf_132_wb_clk_i _02024_ _00625_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[614\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08019__A1 net1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11472_ net2507 net394 _06771_ net512 vssd1 vssd1 vccd1 vccd1 _02027_ sky130_fd_sc_hd__a22o_1
XFILLER_0_52_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_936 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13211_ net1367 vssd1 vssd1 vccd1 vccd1 _00975_ sky130_fd_sc_hd__inv_2
XANTENNA__11778__S net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10423_ _06242_ _06244_ net285 vssd1 vssd1 vccd1 vccd1 _06245_ sky130_fd_sc_hd__mux2_1
XANTENNA__11023__B1 net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_2740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14191_ clknet_leaf_134_wb_clk_i _01955_ _00556_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[545\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_61_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13142_ net1259 vssd1 vssd1 vccd1 vccd1 _00906_ sky130_fd_sc_hd__inv_2
XANTENNA__07557__A net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input63_A gpio_in[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10354_ _06101_ _06187_ _06092_ vssd1 vssd1 vccd1 vccd1 _06188_ sky130_fd_sc_hd__and3b_1
XFILLER_0_131_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_111_2648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_2659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13073_ net1270 vssd1 vssd1 vccd1 vccd1 _00837_ sky130_fd_sc_hd__inv_2
X_10285_ _05973_ _06126_ vssd1 vssd1 vccd1 vccd1 _06127_ sky130_fd_sc_hd__nand2_1
XFILLER_0_20_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08727__C1 net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_163_3715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09772__A net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12024_ _06767_ net462 net360 net2742 vssd1 vssd1 vccd1 vccd1 _01521_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_163_3726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_168_Right_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13294__A net1328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_137_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11629__A2 net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13975_ clknet_leaf_112_wb_clk_i _01739_ _00340_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[329\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10837__A0 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11245__C net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12926_ net1409 vssd1 vssd1 vccd1 vccd1 _00690_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12857_ net1351 vssd1 vssd1 vccd1 vccd1 _00621_ sky130_fd_sc_hd__inv_2
XANTENNA__12638__A net1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11808_ net2656 _06633_ net329 vssd1 vssd1 vccd1 vccd1 _01730_ sky130_fd_sc_hd__mux2_1
X_12788_ net1313 vssd1 vssd1 vccd1 vccd1 _00552_ sky130_fd_sc_hd__inv_2
XFILLER_0_17_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_139_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09012__A _04953_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11261__B _06473_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11262__B1 net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11739_ net1892 net268 net336 vssd1 vssd1 vccd1 vccd1 _01797_ sky130_fd_sc_hd__mux2_1
X_14527_ clknet_leaf_170_wb_clk_i _02291_ _00892_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[881\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_71_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09947__A _03389_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_142_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07481__A2 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14458_ clknet_leaf_147_wb_clk_i _02222_ _00823_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[812\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_796 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_284 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07218__C1 net1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11014__B1 net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13469__A net1328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09758__B2 _04818_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13409_ net1416 vssd1 vssd1 vccd1 vccd1 _01173_ sky130_fd_sc_hd__inv_2
XFILLER_0_40_912 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14389_ clknet_leaf_105_wb_clk_i _02153_ _00754_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[743\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_113_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10368__A2 net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11565__A1 net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_141_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07233__A2 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_176_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__08430__A1 net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08950_ net852 _04884_ _04891_ vssd1 vssd1 vccd1 vccd1 _04892_ sky130_fd_sc_hd__and3_1
XFILLER_0_121_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08997__S net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07901_ net822 _03838_ _03840_ _03842_ net722 vssd1 vssd1 vccd1 vccd1 _03843_ sky130_fd_sc_hd__a41o_1
X_08881_ _04813_ _04814_ _04822_ vssd1 vssd1 vccd1 vccd1 _04823_ sky130_fd_sc_hd__o21ai_1
XPHY_EDGE_ROW_135_Right_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08194__B1 net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_102_Left_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07832_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[426\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[394\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[298\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[266\]
+ net760 net1124 vssd1 vssd1 vccd1 vccd1 _03774_ sky130_fd_sc_hd__mux4_1
XFILLER_0_155_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07941__B1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07763_ net1194 net883 team_03_WB.instance_to_wrap.core.register_file.registers_state\[780\]
+ vssd1 vssd1 vccd1 vccd1 _03705_ sky130_fd_sc_hd__a21o_1
XANTENNA__11436__B net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09502_ team_03_WB.instance_to_wrap.core.decoder.inst\[27\] net1021 net535 _05443_
+ vssd1 vssd1 vccd1 vccd1 _05444_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_2_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08497__A1 net1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07694_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[926\] net793
+ _03635_ vssd1 vssd1 vccd1 vccd1 _03636_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_79_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_154_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09433_ _04648_ _04923_ vssd1 vssd1 vccd1 vccd1 _05375_ sky130_fd_sc_hd__nor2_1
XFILLER_0_2_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_628 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10994__C _06418_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout348_A _06804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11452__A net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09364_ _05278_ _05281_ _05301_ _05193_ vssd1 vssd1 vccd1 vccd1 _05306_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_59_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_111_Left_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08315_ net1064 _04255_ _04256_ net1213 vssd1 vssd1 vccd1 vccd1 _04257_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_23_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10056__B2 team_03_WB.instance_to_wrap.CPU_DAT_O\[7\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09295_ net526 _03490_ _05144_ net609 vssd1 vssd1 vccd1 vccd1 _05237_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_43_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10068__A team_03_WB.instance_to_wrap.core.decoder.inst\[14\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout515_A net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09857__A _05784_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08246_ net1226 team_03_WB.instance_to_wrap.core.register_file.registers_state\[338\]
+ net950 team_03_WB.instance_to_wrap.core.register_file.registers_state\[370\] net1070
+ vssd1 vssd1 vccd1 vccd1 _04188_ sky130_fd_sc_hd__o221a_1
XFILLER_0_34_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_2323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_2334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11598__S net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_969 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08177_ net850 _04103_ _04118_ vssd1 vssd1 vccd1 vccd1 _04119_ sky130_fd_sc_hd__o21a_4
XANTENNA_fanout303_X net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1045_X net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11556__A1 net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_3084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08957__C1 net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07128_ net1109 team_03_WB.instance_to_wrap.core.register_file.registers_state\[704\]
+ net803 team_03_WB.instance_to_wrap.core.register_file.registers_state\[736\] net735
+ vssd1 vssd1 vccd1 vccd1 _03070_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_132_3095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08421__A1 net1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout884_A net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07059_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[674\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[642\]
+ net775 vssd1 vssd1 vccd1 vccd1 _03001_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput160 net160 vssd1 vssd1 vccd1 vccd1 DAT_O[31] sky130_fd_sc_hd__buf_2
XANTENNA_fanout1212_X net1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput171 net171 vssd1 vssd1 vccd1 vccd1 SEL_O[3] sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_120_Left_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput182 net182 vssd1 vssd1 vccd1 vccd1 gpio_oeb[17] sky130_fd_sc_hd__buf_2
Xoutput193 net193 vssd1 vssd1 vccd1 vccd1 gpio_oeb[28] sky130_fd_sc_hd__buf_2
X_10070_ _02800_ _02811_ _05908_ _05913_ net1144 vssd1 vssd1 vccd1 vccd1 _05914_ sky130_fd_sc_hd__o41a_2
XFILLER_0_100_376 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11049__D net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_102_Right_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10531__A2 net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout937_X net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13760_ clknet_leaf_191_wb_clk_i _01524_ _00125_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[114\]
+ sky130_fd_sc_hd__dfrtp_1
X_10972_ _02931_ _05923_ _02829_ net688 vssd1 vssd1 vccd1 vccd1 _06551_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__08488__A1 net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_67_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_168_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12711_ net1369 vssd1 vssd1 vccd1 vccd1 _00475_ sky130_fd_sc_hd__inv_2
XFILLER_0_85_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13691_ clknet_leaf_145_wb_clk_i _01455_ _00056_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[45\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10834__A3 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07160__A1 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_139_3227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_139_3238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12642_ net1296 vssd1 vssd1 vccd1 vccd1 _00406_ sky130_fd_sc_hd__inv_2
XFILLER_0_109_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12036__A2 net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08147__S net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_352 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11244__B1 net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_156_3574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12573_ net1389 vssd1 vssd1 vccd1 vccd1 _00337_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_156_3585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11524_ net280 net620 net703 net695 vssd1 vssd1 vccd1 vccd1 _06781_ sky130_fd_sc_hd__and4_1
XFILLER_0_68_1023 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14312_ clknet_leaf_14_wb_clk_i _02076_ _00677_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[666\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14243_ clknet_leaf_34_wb_clk_i _02007_ _00608_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[597\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11455_ net493 net622 _06580_ net392 net2086 vssd1 vssd1 vccd1 vccd1 _02038_ sky130_fd_sc_hd__a32o_1
XFILLER_0_40_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11301__S net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10406_ team_03_WB.instance_to_wrap.core.pc.current_pc\[14\] _06141_ vssd1 vssd1
+ vccd1 vccd1 _06231_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_22_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08948__C1 net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08412__A1 net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14174_ clknet_leaf_117_wb_clk_i _01938_ _00539_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[528\]
+ sky130_fd_sc_hd__dfrtp_1
X_11386_ net515 net643 _06745_ net403 net2254 vssd1 vssd1 vccd1 vccd1 _02087_ sky130_fd_sc_hd__a32o_1
XFILLER_0_1_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13125_ net1348 vssd1 vssd1 vccd1 vccd1 _00889_ sky130_fd_sc_hd__inv_2
X_10337_ team_03_WB.instance_to_wrap.core.pc.current_pc\[23\] _06147_ _06149_ team_03_WB.instance_to_wrap.core.pc.current_pc\[26\]
+ vssd1 vssd1 vccd1 vccd1 _06174_ sky130_fd_sc_hd__a31o_1
XFILLER_0_0_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06974__A1 net1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13056_ net1403 vssd1 vssd1 vccd1 vccd1 _00820_ sky130_fd_sc_hd__inv_2
X_10268_ _06107_ _06109_ _05979_ vssd1 vssd1 vccd1 vccd1 _06110_ sky130_fd_sc_hd__a21o_1
X_12007_ net1249 net654 net701 net466 vssd1 vssd1 vccd1 vccd1 _06817_ sky130_fd_sc_hd__or4b_4
XFILLER_0_84_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1330 net1438 vssd1 vssd1 vccd1 vccd1 net1330 sky130_fd_sc_hd__clkbuf_4
Xfanout1341 net1342 vssd1 vssd1 vccd1 vccd1 net1341 sky130_fd_sc_hd__buf_4
Xfanout1352 net1358 vssd1 vssd1 vccd1 vccd1 net1352 sky130_fd_sc_hd__buf_2
X_10199_ _04711_ _02774_ net676 vssd1 vssd1 vccd1 vccd1 _06041_ sky130_fd_sc_hd__mux2_1
XFILLER_0_139_1028 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10522__A2 net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_159_wb_clk_i clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_159_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xfanout1363 net1364 vssd1 vssd1 vccd1 vccd1 net1363 sky130_fd_sc_hd__clkbuf_4
Xfanout1374 net1376 vssd1 vssd1 vccd1 vccd1 net1374 sky130_fd_sc_hd__buf_4
XFILLER_0_75_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1385 net1387 vssd1 vssd1 vccd1 vccd1 net1385 sky130_fd_sc_hd__buf_4
XFILLER_0_89_901 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1396 net1398 vssd1 vssd1 vccd1 vccd1 net1396 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_128_2997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08479__A1 net1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09676__B1 net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13958_ clknet_leaf_72_wb_clk_i _01722_ _00323_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[312\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_159_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11483__B1 net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12909_ net1275 vssd1 vssd1 vccd1 vccd1 _00673_ sky130_fd_sc_hd__inv_2
X_13889_ clknet_leaf_180_wb_clk_i _01653_ _00254_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[243\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07151__A1 net1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12027__A2 net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10038__A1 net19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08100__B1 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08100_ net1173 team_03_WB.instance_to_wrap.core.register_file.registers_state\[346\]
+ net759 team_03_WB.instance_to_wrap.core.register_file.registers_state\[378\] net1124
+ vssd1 vssd1 vccd1 vccd1 _04042_ sky130_fd_sc_hd__o221a_1
XANTENNA__11786__A1 _06619_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09080_ net1240 team_03_WB.instance_to_wrap.core.register_file.registers_state\[333\]
+ net982 team_03_WB.instance_to_wrap.core.register_file.registers_state\[365\] net1077
+ vssd1 vssd1 vccd1 vccd1 _05022_ sky130_fd_sc_hd__o221a_1
XFILLER_0_72_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08031_ net1178 team_03_WB.instance_to_wrap.core.register_file.registers_state\[337\]
+ vssd1 vssd1 vccd1 vccd1 _03973_ sky130_fd_sc_hd__or2_1
Xinput40 gpio_in[15] vssd1 vssd1 vccd1 vccd1 net40 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_141_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13199__A net1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput51 gpio_in[26] vssd1 vssd1 vccd1 vccd1 net51 sky130_fd_sc_hd__clkbuf_1
Xinput62 gpio_in[6] vssd1 vssd1 vccd1 vccd1 net62 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_271 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold802 team_03_WB.instance_to_wrap.core.register_file.registers_state\[99\] vssd1
+ vssd1 vccd1 vccd1 net2295 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11211__S net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_720 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_399 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07197__A _03138_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput73 wbs_adr_i[15] vssd1 vssd1 vccd1 vccd1 net73 sky130_fd_sc_hd__clkbuf_1
Xinput84 wbs_adr_i[25] vssd1 vssd1 vccd1 vccd1 net84 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold813 team_03_WB.instance_to_wrap.core.register_file.registers_state\[535\] vssd1
+ vssd1 vccd1 vccd1 net2306 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold824 team_03_WB.instance_to_wrap.core.register_file.registers_state\[139\] vssd1
+ vssd1 vccd1 vccd1 net2317 sky130_fd_sc_hd__dlygate4sd3_1
Xinput95 wbs_adr_i[6] vssd1 vssd1 vccd1 vccd1 net95 sky130_fd_sc_hd__clkbuf_1
Xhold835 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[7\] vssd1 vssd1 vccd1
+ vccd1 net2328 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07628__C net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold846 team_03_WB.instance_to_wrap.core.register_file.registers_state\[510\] vssd1
+ vssd1 vccd1 vccd1 net2339 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_2220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold857 team_03_WB.instance_to_wrap.core.register_file.registers_state\[305\] vssd1
+ vssd1 vccd1 vccd1 net2350 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_2231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07611__C1 net1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09982_ _05861_ net1865 net288 vssd1 vssd1 vccd1 vccd1 _02732_ sky130_fd_sc_hd__mux2_1
Xhold868 team_03_WB.instance_to_wrap.core.register_file.registers_state\[895\] vssd1
+ vssd1 vccd1 vccd1 net2361 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10903__X _06495_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12831__A net1347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold879 team_03_WB.instance_to_wrap.core.register_file.registers_state\[478\] vssd1
+ vssd1 vccd1 vccd1 net2372 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06965__A1 net1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08933_ net1066 _04874_ vssd1 vssd1 vccd1 vccd1 _04875_ sky130_fd_sc_hd__nand2_1
XANTENNA__08520__S net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08167__B1 net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout298_A _06495_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10989__C net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12042__S net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08864_ net1208 _04805_ _04800_ net848 vssd1 vssd1 vccd1 vccd1 _04806_ sky130_fd_sc_hd__a211oi_1
XANTENNA__08262__S0 net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1005_A net1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07815_ net1017 _02835_ team_03_WB.instance_to_wrap.core.decoder.inst\[31\] vssd1
+ vssd1 vccd1 vccd1 _03757_ sky130_fd_sc_hd__o21a_1
X_08795_ _04735_ _04736_ vssd1 vssd1 vccd1 vccd1 _04737_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout465_A net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09116__C1 net1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_2182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_2193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07746_ net1194 team_03_WB.instance_to_wrap.core.register_file.registers_state\[76\]
+ net780 team_03_WB.instance_to_wrap.core.register_file.registers_state\[108\] net731
+ vssd1 vssd1 vccd1 vccd1 _03688_ sky130_fd_sc_hd__o221a_1
XFILLER_0_74_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07660__A _03601_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_3_2_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07677_ net1115 _03615_ _03616_ vssd1 vssd1 vccd1 vccd1 _03619_ sky130_fd_sc_hd__or3_1
XANTENNA_fanout632_A net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12278__A net1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08475__B net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1374_A net1376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09416_ net541 _04505_ _04478_ net559 vssd1 vssd1 vccd1 vccd1 _05358_ sky130_fd_sc_hd__a211o_1
XFILLER_0_149_354 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11182__A net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07693__A2 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_62_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09347_ _04148_ _05287_ vssd1 vssd1 vccd1 vccd1 _05289_ sky130_fd_sc_hd__nand2_1
XFILLER_0_81_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_62_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout420_X net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1162_X net1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11332__D net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout518_X net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_311 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_134_3124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09587__A net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_134_3135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07659__X _03601_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09278_ _04893_ _05219_ vssd1 vssd1 vccd1 vccd1 _05220_ sky130_fd_sc_hd__or2_1
XFILLER_0_106_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_958 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08229_ net1233 team_03_WB.instance_to_wrap.core.register_file.registers_state\[593\]
+ net960 team_03_WB.instance_to_wrap.core.register_file.registers_state\[625\] net919
+ vssd1 vssd1 vccd1 vccd1 _04171_ sky130_fd_sc_hd__o221a_1
XFILLER_0_160_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_151_3471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_151_3482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11240_ net499 net627 _06687_ net408 net2712 vssd1 vssd1 vccd1 vccd1 _02175_ sky130_fd_sc_hd__a32o_1
XANTENNA__10245__B _06086_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout887_X net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07602__C1 net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10960__S net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11171_ net625 _06664_ vssd1 vssd1 vccd1 vccd1 _06665_ sky130_fd_sc_hd__nor2_1
XANTENNA__12741__A net1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06956__A1 net1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10122_ _03640_ _05961_ vssd1 vssd1 vccd1 vccd1 _05964_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_140_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10912__D_N team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[11\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11357__A net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14930_ clknet_leaf_51_wb_clk_i _02685_ _01295_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_O\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_10053_ net3 net1039 net911 team_03_WB.instance_to_wrap.CPU_DAT_O\[10\] vssd1 vssd1
+ vccd1 vccd1 _02678_ sky130_fd_sc_hd__a22o_1
XANTENNA__08002__Y _03944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input26_A DAT_I[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11076__B net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14861_ clknet_leaf_59_wb_clk_i _02625_ _01226_ vssd1 vssd1 vccd1 vccd1 net117 sky130_fd_sc_hd__dfrtp_1
XANTENNA__07381__A1 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11791__S net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13812_ clknet_leaf_133_wb_clk_i _01576_ _00177_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[166\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_106_2547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_742 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14792_ clknet_leaf_94_wb_clk_i _02556_ _01157_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_I\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_106_2558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07570__A net1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_252 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_158_3614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13743_ clknet_leaf_136_wb_clk_i _01507_ _00108_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[97\]
+ sky130_fd_sc_hd__dfrtp_1
X_10955_ net511 net597 net264 net520 net1979 vssd1 vssd1 vccd1 vccd1 _02310_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_158_3625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07133__A1 net1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_123_2894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12009__A2 net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10886_ team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[16\] net307 net688 vssd1
+ vssd1 vccd1 vccd1 _06481_ sky130_fd_sc_hd__a21o_1
X_13674_ clknet_leaf_1_wb_clk_i _01438_ _00039_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07684__A2 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11217__A0 net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12625_ net1266 vssd1 vssd1 vccd1 vccd1 _00389_ sky130_fd_sc_hd__inv_2
XFILLER_0_39_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09497__A net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12556_ net1333 vssd1 vssd1 vccd1 vccd1 _00320_ sky130_fd_sc_hd__inv_2
XANTENNA__08633__A1 net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08605__S net992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09830__B1 net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06914__A net1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_170_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11507_ _06625_ net2653 net390 vssd1 vssd1 vccd1 vccd1 _01999_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07987__A3 net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07841__C1 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12487_ net1369 vssd1 vssd1 vccd1 vccd1 _00251_ sky130_fd_sc_hd__inv_2
XFILLER_0_112_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_777 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_46 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold109 team_03_WB.instance_to_wrap.core.register_file.registers_state\[970\] vssd1
+ vssd1 vccd1 vccd1 net1602 sky130_fd_sc_hd__dlygate4sd3_1
X_11438_ net280 net620 net703 net827 vssd1 vssd1 vccd1 vccd1 _06759_ sky130_fd_sc_hd__and4_1
X_14226_ clknet_leaf_168_wb_clk_i _01990_ _00591_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[580\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_145_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10155__B net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14157_ clknet_leaf_188_wb_clk_i _01921_ _00522_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[511\]
+ sky130_fd_sc_hd__dfrtp_1
X_11369_ net713 net298 net697 vssd1 vssd1 vccd1 vccd1 _06737_ sky130_fd_sc_hd__and3_1
XANTENNA__07295__S1 net1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10743__A2 net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06947__B2 team_03_WB.instance_to_wrap.core.decoder.inst\[24\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13108_ net1308 vssd1 vssd1 vccd1 vccd1 _00872_ sky130_fd_sc_hd__inv_2
X_14088_ clknet_leaf_18_wb_clk_i _01852_ _00453_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[442\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11267__A net1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13039_ net1338 vssd1 vssd1 vccd1 vccd1 _00803_ sky130_fd_sc_hd__inv_2
Xfanout1160 net1161 vssd1 vssd1 vccd1 vccd1 net1160 sky130_fd_sc_hd__buf_4
Xfanout1171 net1180 vssd1 vssd1 vccd1 vccd1 net1171 sky130_fd_sc_hd__clkbuf_4
Xfanout1182 net1183 vssd1 vssd1 vccd1 vccd1 net1182 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__07372__A1 _03313_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1193 net1199 vssd1 vssd1 vccd1 vccd1 net1193 sky130_fd_sc_hd__clkbuf_4
X_15083__1469 vssd1 vssd1 vccd1 vccd1 _15083__1469/HI net1469 sky130_fd_sc_hd__conb_1
X_07600_ net1111 team_03_WB.instance_to_wrap.core.register_file.registers_state\[505\]
+ net902 _03541_ net1159 vssd1 vssd1 vccd1 vccd1 _03542_ sky130_fd_sc_hd__o311a_1
X_08580_ net1049 team_03_WB.instance_to_wrap.core.register_file.registers_state\[669\]
+ net1000 team_03_WB.instance_to_wrap.core.register_file.registers_state\[701\] net922
+ vssd1 vssd1 vccd1 vccd1 _04522_ sky130_fd_sc_hd__a221o_1
XFILLER_0_89_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07531_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[6\] net799
+ net732 _03472_ vssd1 vssd1 vccd1 vccd1 _03473_ sky130_fd_sc_hd__o211a_1
XANTENNA__11456__B1 net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_159_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08295__B net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11206__S net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1155 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07462_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[437\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[405\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[309\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[277\]
+ net772 net1130 vssd1 vssd1 vccd1 vccd1 _03404_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_83_2090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_159_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09201_ net607 _04071_ vssd1 vssd1 vccd1 vccd1 _05143_ sky130_fd_sc_hd__or2_1
XANTENNA__11208__A0 net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07393_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[831\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[799\]
+ net758 vssd1 vssd1 vccd1 vccd1 _03335_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_56_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_56_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_134_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11759__A1 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09132_ _04829_ net322 _05072_ _05073_ _04823_ vssd1 vssd1 vccd1 vccd1 _05074_ sky130_fd_sc_hd__a221o_1
XFILLER_0_17_536 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_wire590_X net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08515__S net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07427__A2 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_161_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09063_ net1081 _05001_ _05004_ net849 vssd1 vssd1 vccd1 vccd1 _05005_ sky130_fd_sc_hd__a31o_1
XANTENNA__10991__D net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08014_ net1115 _03954_ _03955_ vssd1 vssd1 vccd1 vccd1 _03956_ sky130_fd_sc_hd__or3_1
XFILLER_0_60_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold610 team_03_WB.instance_to_wrap.core.register_file.registers_state\[458\] vssd1
+ vssd1 vccd1 vccd1 net2103 sky130_fd_sc_hd__dlygate4sd3_1
Xhold621 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[29\] vssd1 vssd1 vccd1
+ vccd1 net2114 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_230 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10065__B net1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold632 team_03_WB.instance_to_wrap.core.register_file.registers_state\[764\] vssd1
+ vssd1 vccd1 vccd1 net2125 sky130_fd_sc_hd__dlygate4sd3_1
Xhold643 team_03_WB.instance_to_wrap.core.register_file.registers_state\[678\] vssd1
+ vssd1 vccd1 vccd1 net2136 sky130_fd_sc_hd__dlygate4sd3_1
Xhold654 team_03_WB.instance_to_wrap.core.register_file.registers_state\[178\] vssd1
+ vssd1 vccd1 vccd1 net2147 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold665 team_03_WB.instance_to_wrap.core.register_file.registers_state\[827\] vssd1
+ vssd1 vccd1 vccd1 net2158 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12561__A net1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold676 team_03_WB.instance_to_wrap.core.register_file.registers_state\[697\] vssd1
+ vssd1 vccd1 vccd1 net2169 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1122_A _02786_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07060__B1 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold687 team_03_WB.instance_to_wrap.core.register_file.registers_state\[503\] vssd1
+ vssd1 vccd1 vccd1 net2180 sky130_fd_sc_hd__dlygate4sd3_1
Xhold698 team_03_WB.instance_to_wrap.core.register_file.registers_state\[736\] vssd1
+ vssd1 vccd1 vccd1 net2191 sky130_fd_sc_hd__dlygate4sd3_1
X_09965_ _03756_ net661 vssd1 vssd1 vccd1 vccd1 _05887_ sky130_fd_sc_hd__nor2_1
X_08916_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[876\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[844\]
+ net979 vssd1 vssd1 vccd1 vccd1 _04858_ sky130_fd_sc_hd__mux2_1
X_09896_ net1130 _02804_ _05836_ _05837_ vssd1 vssd1 vccd1 vccd1 _05838_ sky130_fd_sc_hd__o211a_1
XANTENNA__09888__B1 _04820_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1008_X net1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11695__B1 net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout370_X net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08847_ net1056 team_03_WB.instance_to_wrap.core.register_file.registers_state\[448\]
+ net1009 team_03_WB.instance_to_wrap.core.register_file.registers_state\[480\] net1078
+ vssd1 vssd1 vccd1 vccd1 _04789_ sky130_fd_sc_hd__a221o_1
XANTENNA__07363__A1 net1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout847_A _06303_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout468_X net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08778_ net862 _04718_ _04719_ _04717_ vssd1 vssd1 vccd1 vccd1 _04720_ sky130_fd_sc_hd__a31o_1
XFILLER_0_169_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_169_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07729_ net1197 team_03_WB.instance_to_wrap.core.register_file.registers_state\[973\]
+ net786 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1005\] net1156
+ vssd1 vssd1 vccd1 vccd1 _03671_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_0_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout635_X net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07115__A1 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_3_3_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_3_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_0_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08312__B1 net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1377_X net1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10740_ team_03_WB.instance_to_wrap.core.pc.current_pc\[11\] _05676_ net605 vssd1
+ vssd1 vccd1 vccd1 _06362_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_0_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_302 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11343__C net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08863__A1 net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_2444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_2455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10671_ _06311_ _05583_ _05563_ vssd1 vssd1 vccd1 vccd1 _06313_ sky130_fd_sc_hd__or3b_1
XANTENNA_fanout802_X net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_153_3511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_153_3522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_311 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12736__A net1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12410_ net1372 vssd1 vssd1 vccd1 vccd1 _00174_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_11_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13390_ net1433 vssd1 vssd1 vccd1 vccd1 _01154_ sky130_fd_sc_hd__inv_2
XFILLER_0_153_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08615__A1 net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12341_ net1272 vssd1 vssd1 vccd1 vccd1 _00105_ sky130_fd_sc_hd__inv_2
XFILLER_0_63_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07549__B _03489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07823__C1 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_161_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15060_ net1446 vssd1 vssd1 vccd1 vccd1 gpio_out[37] sky130_fd_sc_hd__buf_2
XFILLER_0_106_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12272_ net1411 vssd1 vssd1 vccd1 vccd1 _00036_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_79_1992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14011_ clknet_leaf_123_wb_clk_i _01775_ _00376_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[365\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11786__S net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11223_ _06513_ net2273 net489 vssd1 vssd1 vccd1 vccd1 _02187_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_594 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11154_ net1249 net832 _06478_ net671 vssd1 vssd1 vccd1 vccd1 _06654_ sky130_fd_sc_hd__or4_1
X_10105_ team_03_WB.instance_to_wrap.core.pc.current_pc\[1\] net675 vssd1 vssd1 vccd1
+ vccd1 _05949_ sky130_fd_sc_hd__nand2_1
X_11085_ _06620_ net2466 net417 vssd1 vssd1 vccd1 vccd1 _02263_ sky130_fd_sc_hd__mux2_1
X_10036_ net21 net1038 net910 net1650 vssd1 vssd1 vccd1 vccd1 _02695_ sky130_fd_sc_hd__o22a_1
X_14913_ clknet_leaf_43_wb_clk_i _02668_ _01278_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_O\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA_input29_X net29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11686__B1 net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08551__B1 net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14844_ clknet_leaf_87_wb_clk_i net1864 _01209_ vssd1 vssd1 vccd1 vccd1 net130 sky130_fd_sc_hd__dfrtp_1
XANTENNA__08396__A net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06909__A net1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08529__S1 net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11534__B net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14775_ clknet_leaf_95_wb_clk_i _02539_ _01140_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_I\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_11987_ _06468_ net2554 net443 vssd1 vssd1 vccd1 vccd1 _01557_ sky130_fd_sc_hd__mux2_1
XANTENNA__08303__B1 net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13726_ clknet_leaf_121_wb_clk_i _01490_ _00091_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[80\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_458 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10938_ net295 net1991 net521 vssd1 vssd1 vccd1 vccd1 _02313_ sky130_fd_sc_hd__mux2_1
XANTENNA__11253__C net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10661__A1 team_03_WB.instance_to_wrap.CPU_DAT_O\[0\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_155_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09939__B net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10869_ net685 _05833_ vssd1 vssd1 vccd1 vccd1 _06467_ sky130_fd_sc_hd__nand2_1
X_13657_ clknet_leaf_161_wb_clk_i _01421_ _00022_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12646__A net1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_368 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07299__X _03241_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11550__A net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12608_ net1399 vssd1 vssd1 vccd1 vccd1 _00372_ sky130_fd_sc_hd__inv_2
XANTENNA__08335__S net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13588_ net1346 vssd1 vssd1 vccd1 vccd1 _01352_ sky130_fd_sc_hd__inv_2
XFILLER_0_170_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10413__A1 net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08082__A2 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12539_ net1361 vssd1 vssd1 vccd1 vccd1 _00303_ sky130_fd_sc_hd__inv_2
XFILLER_0_170_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09955__A _03942_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_151_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14209_ clknet_leaf_180_wb_clk_i _01973_ _00574_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[563\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_268 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_174_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_174_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__07042__B1 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout408 _06684_ vssd1 vssd1 vccd1 vccd1 net408 sky130_fd_sc_hd__buf_8
Xfanout419 _06610_ vssd1 vssd1 vccd1 vccd1 net419 sky130_fd_sc_hd__buf_4
Xclkbuf_leaf_103_wb_clk_i clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_103_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__07593__A1 net1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09750_ _03727_ net591 vssd1 vssd1 vccd1 vccd1 _05692_ sky130_fd_sc_hd__nor2_1
X_06962_ net1167 _02901_ _02902_ vssd1 vssd1 vccd1 vccd1 _02904_ sky130_fd_sc_hd__and3_1
XANTENNA__09961__Y _05885_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08701_ net1066 _04640_ _04641_ vssd1 vssd1 vccd1 vccd1 _04643_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_33_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09681_ net581 _05501_ _05612_ _05622_ vssd1 vssd1 vccd1 vccd1 _05623_ sky130_fd_sc_hd__a31o_2
XANTENNA__11677__B1 net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06893_ team_03_WB.instance_to_wrap.core.control_logic.instruction\[6\] _02809_ vssd1
+ vssd1 vccd1 vccd1 _02835_ sky130_fd_sc_hd__nor2_1
XANTENNA__08542__B1 net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08632_ net1053 team_03_WB.instance_to_wrap.core.register_file.registers_state\[326\]
+ net1006 team_03_WB.instance_to_wrap.core.register_file.registers_state\[358\] net1215
+ vssd1 vssd1 vccd1 vccd1 _04574_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_85_2130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11429__A0 net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08563_ net431 net424 _04503_ vssd1 vssd1 vccd1 vccd1 _04505_ sky130_fd_sc_hd__nor3_1
XANTENNA__09098__A1 net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_81_2038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07514_ _03451_ _03455_ _03454_ net1121 vssd1 vssd1 vccd1 vccd1 _03456_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__09689__X _05631_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_2049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08494_ net856 _04434_ _04435_ vssd1 vssd1 vccd1 vccd1 _04436_ sky130_fd_sc_hd__or3_1
XFILLER_0_9_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_162_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10652__A1 team_03_WB.instance_to_wrap.CPU_DAT_O\[9\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_9_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07445_ net1115 _03383_ _03384_ vssd1 vssd1 vccd1 vccd1 _03387_ sky130_fd_sc_hd__or3_1
XFILLER_0_58_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout330_A _06810_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08753__B net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1072_A net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07376_ net1175 team_03_WB.instance_to_wrap.core.register_file.registers_state\[191\]
+ net889 net1125 vssd1 vssd1 vccd1 vccd1 _03318_ sky130_fd_sc_hd__a211o_1
XFILLER_0_174_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_161_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09115_ net1051 team_03_WB.instance_to_wrap.core.register_file.registers_state\[974\]
+ net1001 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1006\] net1075
+ vssd1 vssd1 vccd1 vccd1 _05057_ sky130_fd_sc_hd__a221o_1
XFILLER_0_45_675 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11601__A0 _06527_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_143_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10955__A2 net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1337_A net1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_883 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_347 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09046_ net1236 team_03_WB.instance_to_wrap.core.register_file.registers_state\[143\]
+ net971 team_03_WB.instance_to_wrap.core.register_file.registers_state\[175\] net939
+ vssd1 vssd1 vccd1 vccd1 _04988_ sky130_fd_sc_hd__o221a_1
XFILLER_0_5_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout797_A net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold440 team_03_WB.instance_to_wrap.core.register_file.registers_state\[904\] vssd1
+ vssd1 vccd1 vccd1 net1933 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09022__A1 net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07259__S1 net1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1125_X net1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold451 team_03_WB.instance_to_wrap.core.register_file.registers_state\[62\] vssd1
+ vssd1 vccd1 vccd1 net1944 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10707__A2 net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11904__A1 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold462 team_03_WB.instance_to_wrap.core.register_file.registers_state\[694\] vssd1
+ vssd1 vccd1 vccd1 net1955 sky130_fd_sc_hd__dlygate4sd3_1
Xhold473 team_03_WB.instance_to_wrap.core.register_file.registers_state\[675\] vssd1
+ vssd1 vccd1 vccd1 net1966 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07033__B1 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_3023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold484 team_03_WB.instance_to_wrap.core.register_file.registers_state\[907\] vssd1
+ vssd1 vccd1 vccd1 net1977 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08230__C1 net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_3034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold495 team_03_WB.instance_to_wrap.core.register_file.registers_state\[430\] vssd1
+ vssd1 vccd1 vccd1 net1988 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout585_X net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout964_A net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout920 net922 vssd1 vssd1 vccd1 vccd1 net920 sky130_fd_sc_hd__buf_4
XANTENNA__07584__A1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout931 net932 vssd1 vssd1 vccd1 vccd1 net931 sky130_fd_sc_hd__clkbuf_2
XANTENNA__11380__A2 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09948_ _05878_ net1811 net292 vssd1 vssd1 vccd1 vccd1 _02753_ sky130_fd_sc_hd__mux2_1
Xfanout942 net943 vssd1 vssd1 vccd1 vccd1 net942 sky130_fd_sc_hd__buf_4
Xfanout953 net955 vssd1 vssd1 vccd1 vccd1 net953 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_146_3370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout964 net965 vssd1 vssd1 vccd1 vccd1 net964 sky130_fd_sc_hd__clkbuf_4
Xfanout975 net976 vssd1 vssd1 vccd1 vccd1 net975 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_146_3381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout986 net987 vssd1 vssd1 vccd1 vccd1 net986 sky130_fd_sc_hd__clkbuf_4
X_09879_ _05635_ _05813_ _05820_ vssd1 vssd1 vccd1 vccd1 _05821_ sky130_fd_sc_hd__o21ba_2
XTAP_TAPCELL_ROW_5_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11057__D net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout997 _04085_ vssd1 vssd1 vccd1 vccd1 net997 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout752_X net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1140 team_03_WB.instance_to_wrap.core.register_file.registers_state\[203\] vssd1
+ vssd1 vccd1 vccd1 net2633 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1151 team_03_WB.instance_to_wrap.core.register_file.registers_state\[842\] vssd1
+ vssd1 vccd1 vccd1 net2644 sky130_fd_sc_hd__dlygate4sd3_1
X_11910_ _06611_ net2467 net367 vssd1 vssd1 vccd1 vccd1 _01632_ sky130_fd_sc_hd__mux2_1
Xhold1162 team_03_WB.instance_to_wrap.core.register_file.registers_state\[781\] vssd1
+ vssd1 vccd1 vccd1 net2655 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1173 team_03_WB.instance_to_wrap.core.register_file.registers_state\[513\] vssd1
+ vssd1 vccd1 vccd1 net2666 sky130_fd_sc_hd__dlygate4sd3_1
X_12890_ net1373 vssd1 vssd1 vccd1 vccd1 _00654_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_142_3289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1184 team_03_WB.instance_to_wrap.core.register_file.registers_state\[839\] vssd1
+ vssd1 vccd1 vccd1 net2677 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1195 team_03_WB.instance_to_wrap.core.register_file.registers_state\[705\] vssd1
+ vssd1 vccd1 vccd1 net2688 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10891__A1 net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09089__A1 net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11841_ _06679_ net477 net325 net2524 vssd1 vssd1 vccd1 vccd1 _01698_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_16_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_211 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09599__X _05541_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_2831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_120_2842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14560_ clknet_leaf_192_wb_clk_i _02324_ _00925_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[914\]
+ sky130_fd_sc_hd__dfrtp_1
X_11772_ _06605_ net468 net333 net2632 vssd1 vssd1 vccd1 vccd1 _01765_ sky130_fd_sc_hd__a22o_1
XANTENNA__12093__B1 net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_704 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10723_ team_03_WB.instance_to_wrap.core.pc.current_pc\[19\] net602 vssd1 vssd1 vccd1
+ vccd1 _06353_ sky130_fd_sc_hd__or2_1
X_13511_ net1321 vssd1 vssd1 vccd1 vccd1 _01275_ sky130_fd_sc_hd__inv_2
XANTENNA__11840__B1 net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14491_ clknet_leaf_125_wb_clk_i _02255_ _00856_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[845\]
+ sky130_fd_sc_hd__dfrtp_1
X_13442_ net1423 vssd1 vssd1 vccd1 vccd1 _01206_ sky130_fd_sc_hd__inv_2
XFILLER_0_138_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10654_ net1252 team_03_WB.instance_to_wrap.CPU_DAT_O\[7\] net846 vssd1 vssd1 vccd1
+ vccd1 _02474_ sky130_fd_sc_hd__mux2_1
XANTENNA_input93_A wbs_adr_i[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_647 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13373_ net1416 vssd1 vssd1 vccd1 vccd1 _01137_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10585_ net1600 net534 net601 net593 vssd1 vssd1 vccd1 vccd1 _02538_ sky130_fd_sc_hd__a22o_1
Xclkload18 clknet_leaf_6_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload18/Y sky130_fd_sc_hd__clkinv_4
Xclkload29 clknet_leaf_174_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload29/X sky130_fd_sc_hd__clkbuf_8
X_15112_ net1485 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[17] sky130_fd_sc_hd__buf_2
X_15082__1468 vssd1 vssd1 vccd1 vccd1 _15082__1468/HI net1468 sky130_fd_sc_hd__conb_1
XFILLER_0_152_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_118_2793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12324_ net1374 vssd1 vssd1 vccd1 vccd1 _00088_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_1_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_1_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_23_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15043_ clknet_leaf_82_wb_clk_i _02763_ _01408_ vssd1 vssd1 vccd1 vccd1 net199 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12255_ net1348 vssd1 vssd1 vccd1 vccd1 _00019_ sky130_fd_sc_hd__inv_2
XFILLER_0_142_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_43_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_50_199 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06911__B net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11206_ _06434_ net2414 net487 vssd1 vssd1 vccd1 vccd1 _02202_ sky130_fd_sc_hd__mux2_1
XANTENNA__07024__B1 net1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12186_ net1538 vssd1 vssd1 vccd1 vccd1 _02367_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_166_3779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11137_ net2034 net415 _06644_ net515 vssd1 vssd1 vccd1 vccd1 _02235_ sky130_fd_sc_hd__a22o_1
XANTENNA__08119__A3 net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11068_ net837 _06414_ vssd1 vssd1 vccd1 vccd1 _06612_ sky130_fd_sc_hd__nor2_2
XANTENNA__11123__A2 net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08524__B1 net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08838__B net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10019_ net80 net79 net82 net81 vssd1 vssd1 vccd1 vccd1 _05897_ sky130_fd_sc_hd__or4_1
X_14827_ clknet_leaf_90_wb_clk_i net1697 _01192_ vssd1 vssd1 vccd1 vccd1 net148 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_149_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12084__B1 net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14758_ clknet_leaf_54_wb_clk_i _02522_ _01123_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08827__A1 net1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_157_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13709_ clknet_leaf_182_wb_clk_i _01473_ _00074_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[63\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_117_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11831__B1 net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14689_ clknet_leaf_59_wb_clk_i _02453_ _01054_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.ADR_I\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_156_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_759 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07230_ net1096 team_03_WB.instance_to_wrap.core.register_file.registers_state\[808\]
+ net896 vssd1 vssd1 vccd1 vccd1 _03172_ sky130_fd_sc_hd__or3_1
XFILLER_0_27_642 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_82_wb_clk_i_A clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_172_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07161_ _03075_ _03081_ _03102_ vssd1 vssd1 vccd1 vccd1 _03103_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_82_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07092_ net1198 team_03_WB.instance_to_wrap.core.register_file.registers_state\[737\]
+ net884 _03033_ vssd1 vssd1 vccd1 vccd1 _03034_ sky130_fd_sc_hd__a31o_1
XFILLER_0_112_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09004__A1 net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08438__S0 net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11898__B1 net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07636__C net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07566__A1 net1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11362__A2 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09802_ net537 _05741_ _05743_ vssd1 vssd1 vccd1 vccd1 _05744_ sky130_fd_sc_hd__o21ai_1
X_07994_ net1203 team_03_WB.instance_to_wrap.core.register_file.registers_state\[720\]
+ net786 team_03_WB.instance_to_wrap.core.register_file.registers_state\[752\] net752
+ vssd1 vssd1 vccd1 vccd1 _03936_ sky130_fd_sc_hd__o221a_1
XANTENNA__10570__B1 net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09733_ _05673_ _05674_ _05668_ vssd1 vssd1 vccd1 vccd1 _05675_ sky130_fd_sc_hd__a21o_1
X_06945_ _02881_ _02886_ net823 vssd1 vssd1 vccd1 vccd1 _02887_ sky130_fd_sc_hd__mux2_1
XANTENNA__07318__A1 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout280_A _06409_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout378_A _06812_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12050__S net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09664_ _03170_ _04207_ net664 _05605_ vssd1 vssd1 vccd1 vccd1 _05606_ sky130_fd_sc_hd__a22o_1
X_06876_ _02814_ net1017 vssd1 vssd1 vccd1 vccd1 _02818_ sky130_fd_sc_hd__or2_4
X_08615_ net1058 team_03_WB.instance_to_wrap.core.register_file.registers_state\[197\]
+ net1012 team_03_WB.instance_to_wrap.core.register_file.registers_state\[229\] net931
+ vssd1 vssd1 vccd1 vccd1 _04557_ sky130_fd_sc_hd__a221o_1
X_09595_ net573 _05535_ _05536_ _04832_ _05534_ vssd1 vssd1 vccd1 vccd1 _05537_ sky130_fd_sc_hd__a311o_1
Xclkbuf_leaf_71_wb_clk_i clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_71_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout545_A _03106_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08818__A1 net1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12075__B1 net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08546_ net1049 team_03_WB.instance_to_wrap.core.register_file.registers_state\[702\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[670\] net1000 net933
+ vssd1 vssd1 vccd1 vccd1 _04488_ sky130_fd_sc_hd__o221a_1
XANTENNA__07177__S0 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10625__A1 team_03_WB.instance_to_wrap.CPU_DAT_O\[4\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_08477_ net1048 team_03_WB.instance_to_wrap.core.register_file.registers_state\[667\]
+ net999 team_03_WB.instance_to_wrap.core.register_file.registers_state\[699\] net929
+ vssd1 vssd1 vccd1 vccd1 _04419_ sky130_fd_sc_hd__a221o_1
XANTENNA__11822__B1 net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout712_A net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout333_X net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1075_X net1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11190__A net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07428_ net1084 team_03_WB.instance_to_wrap.core.register_file.registers_state\[820\]
+ net889 vssd1 vssd1 vccd1 vccd1 _03370_ sky130_fd_sc_hd__or3_1
XFILLER_0_18_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_165_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_162_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_455 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout500_X net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07359_ net1172 team_03_WB.instance_to_wrap.core.register_file.registers_state\[860\]
+ net759 team_03_WB.instance_to_wrap.core.register_file.registers_state\[892\] net1124
+ vssd1 vssd1 vccd1 vccd1 _03301_ sky130_fd_sc_hd__o221a_1
XFILLER_0_163_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_98_2387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1242_X net1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_2398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10928__A2 net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10370_ _06200_ _06201_ team_03_WB.instance_to_wrap.core.pc.current_pc\[21\] net677
+ vssd1 vssd1 vccd1 vccd1 _02655_ sky130_fd_sc_hd__o2bb2a_1
XPHY_EDGE_ROW_149_Right_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11050__B2 net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08703__S net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10805__Y _06413_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_1940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09029_ net1244 team_03_WB.instance_to_wrap.core.register_file.registers_state\[592\]
+ net989 team_03_WB.instance_to_wrap.core.register_file.registers_state\[624\] net930
+ vssd1 vssd1 vccd1 vccd1 _04971_ sky130_fd_sc_hd__o221a_1
XFILLER_0_103_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_148_3410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_148_3421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12040_ net1250 net656 _06463_ net473 vssd1 vssd1 vccd1 vccd1 _06818_ sky130_fd_sc_hd__or4b_4
Xhold270 net221 vssd1 vssd1 vccd1 vccd1 net1763 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_113_2690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11889__B1 net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11349__B net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold281 _02585_ vssd1 vssd1 vccd1 vccd1 net1774 sky130_fd_sc_hd__dlygate4sd3_1
Xhold292 team_03_WB.instance_to_wrap.CPU_DAT_O\[25\] vssd1 vssd1 vccd1 vccd1 net1785
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_72_1848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08754__B1 net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_1859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10821__X _06426_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10561__B1 net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_144_3329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_127_wb_clk_i_A clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout750 net754 vssd1 vssd1 vccd1 vccd1 net750 sky130_fd_sc_hd__buf_4
Xfanout761 net773 vssd1 vssd1 vccd1 vccd1 net761 sky130_fd_sc_hd__buf_2
XFILLER_0_102_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout772 net773 vssd1 vssd1 vccd1 vccd1 net772 sky130_fd_sc_hd__buf_2
XANTENNA__07309__A1 net1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout783 net790 vssd1 vssd1 vccd1 vccd1 net783 sky130_fd_sc_hd__clkbuf_4
X_13991_ clknet_leaf_113_wb_clk_i _01755_ _00356_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[345\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout794 net795 vssd1 vssd1 vccd1 vccd1 net794 sky130_fd_sc_hd__buf_4
XANTENNA__11365__A net1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_161_3676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12942_ net1310 vssd1 vssd1 vccd1 vccd1 _00706_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_161_3687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11084__B net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12873_ net1253 vssd1 vssd1 vccd1 vccd1 _00637_ sky130_fd_sc_hd__inv_2
X_14612_ clknet_leaf_132_wb_clk_i _02376_ _00977_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[966\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__12066__A0 _06528_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07989__S net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11824_ _06655_ net462 net323 net2350 vssd1 vssd1 vccd1 vccd1 _01715_ sky130_fd_sc_hd__a22o_1
XFILLER_0_139_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14543_ clknet_leaf_135_wb_clk_i _02307_ _00908_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[897\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11813__B1 net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11755_ net647 _06580_ net454 net331 net2248 vssd1 vssd1 vccd1 vccd1 _01782_ sky130_fd_sc_hd__a32o_1
XANTENNA__11304__S net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06906__B net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10706_ _06341_ _06342_ net606 vssd1 vssd1 vccd1 vccd1 _06343_ sky130_fd_sc_hd__mux2_1
XFILLER_0_127_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14474_ clknet_leaf_6_wb_clk_i _02238_ _00839_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[828\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_153_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11686_ _06728_ net381 net339 net1797 vssd1 vssd1 vccd1 vccd1 _01848_ sky130_fd_sc_hd__a22o_1
XFILLER_0_126_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13425_ net1421 vssd1 vssd1 vccd1 vccd1 _01189_ sky130_fd_sc_hd__inv_2
X_10637_ team_03_WB.instance_to_wrap.core.decoder.inst\[24\] team_03_WB.instance_to_wrap.CPU_DAT_O\[24\]
+ _06303_ vssd1 vssd1 vccd1 vccd1 _02491_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08037__A2 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkload107 clknet_leaf_155_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload107/Y sky130_fd_sc_hd__clkinv_2
XANTENNA__10919__A2 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkload118 clknet_leaf_162_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload118/Y sky130_fd_sc_hd__inv_8
XFILLER_0_140_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_153_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkload129 clknet_leaf_142_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload129/Y sky130_fd_sc_hd__clkinv_2
X_10568_ net1696 net531 net598 _05878_ vssd1 vssd1 vccd1 vccd1 _02555_ sky130_fd_sc_hd__a22o_1
XANTENNA__09785__A2 _04619_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13356_ net1318 vssd1 vssd1 vccd1 vccd1 _01120_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_116_Right_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_667 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06922__A team_03_WB.instance_to_wrap.core.decoder.inst\[24\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_166_wb_clk_i_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_87_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_168_3819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12307_ net1256 vssd1 vssd1 vccd1 vccd1 _00071_ sky130_fd_sc_hd__inv_2
XFILLER_0_121_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13287_ net1343 vssd1 vssd1 vccd1 vccd1 _01051_ sky130_fd_sc_hd__inv_2
X_10499_ net1594 net1030 net907 net1562 vssd1 vssd1 vccd1 vccd1 _02610_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_15_Left_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15026_ clknet_leaf_104_wb_clk_i _02746_ _01391_ vssd1 vssd1 vccd1 vccd1 net182 sky130_fd_sc_hd__dfrtp_1
X_12238_ net2727 vssd1 vssd1 vccd1 vccd1 _01419_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__11259__B _06468_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07456__C net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11344__A2 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12169_ net1635 vssd1 vssd1 vccd1 vccd1 _02384_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__11895__A3 net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08849__A net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07753__A net1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput5 DAT_I[12] vssd1 vssd1 vccd1 vccd1 net5 sky130_fd_sc_hd__clkbuf_1
XANTENNA__11275__A net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07181__C1 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_1132 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07720__A1 net1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_21 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12057__A0 _06623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08400_ net1246 team_03_WB.instance_to_wrap.core.register_file.registers_state\[729\]
+ net991 team_03_WB.instance_to_wrap.core.register_file.registers_state\[761\] net947
+ vssd1 vssd1 vccd1 vccd1 _04342_ sky130_fd_sc_hd__o221a_1
X_09380_ _03566_ _05158_ vssd1 vssd1 vccd1 vccd1 _05322_ sky130_fd_sc_hd__xor2_1
XFILLER_0_47_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08331_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[629\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[597\]
+ net968 vssd1 vssd1 vccd1 vccd1 _04273_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_3_7_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09399__B _04475_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07484__B1 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08262_ _04200_ _04201_ _04202_ _04203_ net859 net934 vssd1 vssd1 vccd1 vccd1 _04204_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__11280__A1 net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07213_ net1114 _03153_ _03154_ vssd1 vssd1 vccd1 vccd1 _03155_ sky130_fd_sc_hd__or3_1
X_08193_ net1231 team_03_WB.instance_to_wrap.core.register_file.registers_state\[595\]
+ net957 team_03_WB.instance_to_wrap.core.register_file.registers_state\[627\] net918
+ vssd1 vssd1 vccd1 vccd1 _04135_ sky130_fd_sc_hd__o221a_1
XFILLER_0_15_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07144_ net735 _03082_ _03083_ _03084_ _03085_ vssd1 vssd1 vccd1 vccd1 _03086_ sky130_fd_sc_hd__a32o_1
XFILLER_0_125_680 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07787__A1 net1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07331__S0 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08984__B1 net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07075_ net1095 team_03_WB.instance_to_wrap.core.register_file.registers_state\[450\]
+ vssd1 vssd1 vccd1 vccd1 _03017_ sky130_fd_sc_hd__and2_1
XANTENNA__12045__S net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_2284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_2295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07539__A1 net1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout495_A net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09862__B _05281_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10543__B1 net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1202_A net1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11886__A3 net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout283_X net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout662_A net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07977_ _03916_ _03918_ net1167 vssd1 vssd1 vccd1 vccd1 _03919_ sky130_fd_sc_hd__o21a_1
X_09716_ _04832_ _05548_ vssd1 vssd1 vccd1 vccd1 _05658_ sky130_fd_sc_hd__or2_1
X_06928_ net1158 net1120 vssd1 vssd1 vccd1 vccd1 _02870_ sky130_fd_sc_hd__nand2_4
XFILLER_0_93_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09700__A2 net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15081__1467 vssd1 vssd1 vccd1 vccd1 _15081__1467/HI net1467 sky130_fd_sc_hd__conb_1
X_09647_ net1120 _02804_ net535 _05588_ vssd1 vssd1 vccd1 vccd1 _05589_ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout450_X net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06859_ team_03_WB.instance_to_wrap.core.control_logic.instruction\[6\] team_03_WB.instance_to_wrap.core.control_logic.instruction\[5\]
+ team_03_WB.instance_to_wrap.core.control_logic.instruction\[4\] vssd1 vssd1 vccd1
+ vccd1 _02801_ sky130_fd_sc_hd__and3b_2
XANTENNA__07172__C1 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07711__A1 net1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout927_A net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09578_ net570 _05399_ vssd1 vssd1 vccd1 vccd1 _05520_ sky130_fd_sc_hd__nand2_1
XANTENNA__08494__A net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_155_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08529_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[447\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[415\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[319\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[287\]
+ net952 net1070 vssd1 vssd1 vccd1 vccd1 _04471_ sky130_fd_sc_hd__mux4_1
XANTENNA__08267__A2 _04079_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout715_X net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07475__B1 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11540_ net502 net629 _06650_ net483 net1705 vssd1 vssd1 vccd1 vccd1 _01975_ sky130_fd_sc_hd__a32o_1
XFILLER_0_93_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11351__C net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_162_230 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_3188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11471_ net658 _06596_ vssd1 vssd1 vccd1 vccd1 _06771_ sky130_fd_sc_hd__nor2_1
XANTENNA__10816__X _06422_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09216__A1 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_740 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10422_ _06064_ _06243_ vssd1 vssd1 vccd1 vccd1 _06244_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_151_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13210_ net1377 vssd1 vssd1 vccd1 vccd1 _00974_ sky130_fd_sc_hd__inv_2
XANTENNA__11023__A1 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_2730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14190_ clknet_leaf_124_wb_clk_i _01954_ _00555_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[544\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_115_2741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07778__A1 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14732__Q team_03_WB.instance_to_wrap.core.decoder.inst\[29\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10353_ _06104_ _06089_ vssd1 vssd1 vccd1 vccd1 _06187_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_33_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13141_ net1292 vssd1 vssd1 vccd1 vccd1 _00905_ sky130_fd_sc_hd__inv_2
XANTENNA__10782__B1 net1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_374 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13072_ net1412 vssd1 vssd1 vccd1 vccd1 _00836_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_111_2649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input56_A gpio_in[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10284_ _06125_ _06123_ vssd1 vssd1 vccd1 vccd1 _06126_ sky130_fd_sc_hd__nand2b_1
XANTENNA__11794__S net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08727__B1 net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12023_ net641 _06585_ net474 net362 net2388 vssd1 vssd1 vccd1 vccd1 _01522_ sky130_fd_sc_hd__a32o_1
XFILLER_0_104_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_163_3716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_163_3727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10534__B1 net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11877__A3 net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07573__A net1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout580 _02992_ vssd1 vssd1 vccd1 vccd1 net580 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11095__A net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13974_ clknet_leaf_178_wb_clk_i _01738_ _00339_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[328\]
+ sky130_fd_sc_hd__dfrtp_1
X_12925_ net1383 vssd1 vssd1 vccd1 vccd1 _00689_ sky130_fd_sc_hd__inv_2
XFILLER_0_158_503 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07702__A1 net1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11245__D net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12039__B1 net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12856_ net1381 vssd1 vssd1 vccd1 vccd1 _00620_ sky130_fd_sc_hd__inv_2
XFILLER_0_158_547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11807_ net2409 _06632_ net330 vssd1 vssd1 vccd1 vccd1 _01731_ sky130_fd_sc_hd__mux2_1
XFILLER_0_127_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12787_ net1271 vssd1 vssd1 vccd1 vccd1 _00551_ sky130_fd_sc_hd__inv_2
XFILLER_0_154_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07466__B1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11262__A1 net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14526_ clknet_leaf_114_wb_clk_i _02290_ _00891_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[880\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_25_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11261__C net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11738_ net597 net264 net473 _06808_ net1844 vssd1 vssd1 vccd1 vccd1 _01798_ sky130_fd_sc_hd__a32o_1
XFILLER_0_3_1051 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10158__B net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07561__S0 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09947__B net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14457_ clknet_leaf_175_wb_clk_i _02221_ _00822_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[811\]
+ sky130_fd_sc_hd__dfrtp_1
X_11669_ net2674 net265 net344 vssd1 vssd1 vccd1 vccd1 _01864_ sky130_fd_sc_hd__mux2_1
XFILLER_0_142_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11014__A1 net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07748__A net1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13408_ net1415 vssd1 vssd1 vccd1 vccd1 _01172_ sky130_fd_sc_hd__inv_2
XFILLER_0_98_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09758__A2 _04922_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08415__C1 net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14388_ clknet_leaf_133_wb_clk_i _02152_ _00753_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[742\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11565__A2 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_795 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13339_ net1334 vssd1 vssd1 vccd1 vccd1 _01103_ sky130_fd_sc_hd__inv_2
XANTENNA__10174__A team_03_WB.instance_to_wrap.core.decoder.inst\[30\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09963__A _03723_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08981__A3 _04922_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15009_ clknet_leaf_51_wb_clk_i net57 _01374_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_07900_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[271\] net781
+ _03841_ vssd1 vssd1 vccd1 vccd1 _03842_ sky130_fd_sc_hd__a21o_1
X_08880_ net556 _04770_ net537 _04819_ vssd1 vssd1 vccd1 vccd1 _04822_ sky130_fd_sc_hd__o31a_1
XANTENNA__10902__A team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[13\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10525__B1 net1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07831_ _03769_ _03770_ _03772_ net1123 vssd1 vssd1 vccd1 vccd1 _03773_ sky130_fd_sc_hd__o22a_1
XFILLER_0_138_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07941__A1 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11209__S net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07762_ net1098 team_03_WB.instance_to_wrap.core.register_file.registers_state\[812\]
+ net897 vssd1 vssd1 vccd1 vccd1 _03704_ sky130_fd_sc_hd__or3_1
XANTENNA__11436__C net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09501_ _03823_ _04444_ vssd1 vssd1 vccd1 vccd1 _05443_ sky130_fd_sc_hd__or2_1
XFILLER_0_79_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07693_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[958\] net767
+ net1014 vssd1 vssd1 vccd1 vccd1 _03635_ sky130_fd_sc_hd__o21a_1
XFILLER_0_2_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09432_ _05372_ _05373_ net558 vssd1 vssd1 vccd1 vccd1 _05374_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09203__A net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10994__D net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09363_ _05291_ _05303_ _05304_ _05288_ vssd1 vssd1 vccd1 vccd1 _05305_ sky130_fd_sc_hd__o211a_1
XFILLER_0_19_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10056__A2 net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08314_ net1237 team_03_WB.instance_to_wrap.core.register_file.registers_state\[856\]
+ net973 team_03_WB.instance_to_wrap.core.register_file.registers_state\[888\] net1219
+ vssd1 vssd1 vccd1 vccd1 _04256_ sky130_fd_sc_hd__o221a_1
XFILLER_0_47_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09294_ _05226_ _05228_ vssd1 vssd1 vccd1 vccd1 _05236_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_23_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10068__B team_03_WB.instance_to_wrap.core.decoder.inst\[13\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08245_ net859 _04183_ _04186_ vssd1 vssd1 vccd1 vccd1 _04187_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_90_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_160_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09857__B _05798_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout410_A _06684_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1152_A net1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_95_2324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout508_A net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_2335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_734 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09749__A2 _05570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08176_ net1207 _04110_ _04117_ net850 vssd1 vssd1 vccd1 vccd1 _04118_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_42_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11556__A2 net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07127_ net1198 team_03_WB.instance_to_wrap.core.register_file.registers_state\[672\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[640\] net785 net735
+ vssd1 vssd1 vccd1 vccd1 _03069_ sky130_fd_sc_hd__a221o_1
XANTENNA__08957__B1 net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_3085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_3096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10764__B1 net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1038_X net1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07058_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[546\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[514\]
+ net775 vssd1 vssd1 vccd1 vccd1 _03000_ sky130_fd_sc_hd__mux2_1
Xoutput150 net150 vssd1 vssd1 vccd1 vccd1 DAT_O[22] sky130_fd_sc_hd__buf_2
XANTENNA_fanout877_A net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput161 net161 vssd1 vssd1 vccd1 vccd1 DAT_O[3] sky130_fd_sc_hd__buf_2
Xoutput172 net172 vssd1 vssd1 vccd1 vccd1 STB_O sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout498_X net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11908__A net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput183 net183 vssd1 vssd1 vccd1 vccd1 gpio_oeb[18] sky130_fd_sc_hd__buf_2
XANTENNA__10516__B1 net1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput194 net194 vssd1 vssd1 vccd1 vccd1 gpio_oeb[29] sky130_fd_sc_hd__buf_2
XANTENNA_fanout1205_X net1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09921__A2 _05453_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11119__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10819__A1 net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10971_ net267 net2232 net520 vssd1 vssd1 vccd1 vccd1 _02307_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout832_X net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09685__B2 _04178_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11643__A net1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12710_ net1299 vssd1 vssd1 vccd1 vccd1 _00474_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_67_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13690_ clknet_leaf_142_wb_clk_i _01454_ _00055_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[44\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_139_3228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14727__Q team_03_WB.instance_to_wrap.core.decoder.inst\[24\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_139_3239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12641_ net1290 vssd1 vssd1 vccd1 vccd1 _00405_ sky130_fd_sc_hd__inv_2
XFILLER_0_167_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10047__A2 net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11244__A1 net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07448__B1 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12572_ net1416 vssd1 vssd1 vccd1 vccd1 _00336_ sky130_fd_sc_hd__inv_2
XANTENNA__08645__C1 net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_156_3575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_156_3586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07999__A1 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14311_ clknet_leaf_110_wb_clk_i _02075_ _00676_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[665\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11789__S net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11523_ net2262 net482 _06780_ net493 vssd1 vssd1 vccd1 vccd1 _01985_ sky130_fd_sc_hd__a22o_1
XFILLER_0_163_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12474__A net1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14242_ clknet_leaf_184_wb_clk_i _02006_ _00607_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[596\]
+ sky130_fd_sc_hd__dfrtp_1
X_11454_ net500 net627 _06579_ net395 net2203 vssd1 vssd1 vccd1 vccd1 _02039_ sky130_fd_sc_hd__a32o_1
XFILLER_0_33_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10204__C1 _02994_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10405_ net284 _06229_ vssd1 vssd1 vccd1 vccd1 _06230_ sky130_fd_sc_hd__and2_1
X_11385_ net715 net269 net700 vssd1 vssd1 vccd1 vccd1 _06745_ sky130_fd_sc_hd__and3_1
X_14173_ clknet_leaf_26_wb_clk_i _01937_ _00538_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[527\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_68_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06959__C1 net1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13124_ net1385 vssd1 vssd1 vccd1 vccd1 _00888_ sky130_fd_sc_hd__inv_2
X_10336_ _06172_ _06173_ team_03_WB.instance_to_wrap.core.pc.current_pc\[27\] net679
+ vssd1 vssd1 vccd1 vccd1 _02661_ sky130_fd_sc_hd__o2bb2a_1
X_10267_ _05979_ _06108_ vssd1 vssd1 vccd1 vccd1 _06109_ sky130_fd_sc_hd__nor2_1
X_13055_ net1349 vssd1 vssd1 vccd1 vccd1 _00819_ sky130_fd_sc_hd__inv_2
XANTENNA__08176__A1 net1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1320 net1330 vssd1 vssd1 vccd1 vccd1 net1320 sky130_fd_sc_hd__buf_2
X_12006_ net266 net2684 net444 vssd1 vssd1 vccd1 vccd1 _01538_ sky130_fd_sc_hd__mux2_1
XFILLER_0_139_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1331 net1339 vssd1 vssd1 vccd1 vccd1 net1331 sky130_fd_sc_hd__buf_4
X_10198_ team_03_WB.instance_to_wrap.core.pc.current_pc\[4\] net660 _06038_ _02889_
+ vssd1 vssd1 vccd1 vccd1 _06040_ sky130_fd_sc_hd__o211a_1
Xfanout1342 net1346 vssd1 vssd1 vccd1 vccd1 net1342 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07384__C1 net1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1353 net1354 vssd1 vssd1 vccd1 vccd1 net1353 sky130_fd_sc_hd__buf_4
XFILLER_0_79_1153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1364 net1437 vssd1 vssd1 vccd1 vccd1 net1364 sky130_fd_sc_hd__buf_2
Xfanout1375 net1376 vssd1 vssd1 vccd1 vccd1 net1375 sky130_fd_sc_hd__buf_4
Xfanout1386 net1387 vssd1 vssd1 vccd1 vccd1 net1386 sky130_fd_sc_hd__buf_4
XFILLER_0_89_913 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1397 net1398 vssd1 vssd1 vccd1 vccd1 net1397 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_128_2998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13957_ clknet_leaf_37_wb_clk_i _01721_ _00322_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[311\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09676__A1 _03391_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07136__C1 net1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12908_ net1314 vssd1 vssd1 vccd1 vccd1 _00672_ sky130_fd_sc_hd__inv_2
XANTENNA__11483__A1 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07687__B1 net1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08338__S net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13888_ clknet_leaf_190_wb_clk_i _01652_ _00253_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[242\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_128_wb_clk_i clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_128_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_159_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_523 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12839_ net1400 vssd1 vssd1 vccd1 vccd1 _00603_ sky130_fd_sc_hd__inv_2
XANTENNA__10169__A _04893_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_174_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_158_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10038__A2 net1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08862__A net1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08100__A1 net1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10996__C_N _06422_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14509_ clknet_leaf_189_wb_clk_i _02273_ _00874_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[863\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_142_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08030_ net811 _03967_ _03968_ _03971_ vssd1 vssd1 vccd1 vccd1 _03972_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_115_959 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput30 DAT_I[6] vssd1 vssd1 vccd1 vccd1 net30 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_4_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput41 gpio_in[16] vssd1 vssd1 vccd1 vccd1 net41 sky130_fd_sc_hd__clkbuf_1
Xinput52 gpio_in[27] vssd1 vssd1 vccd1 vccd1 net52 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_141_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput63 gpio_in[7] vssd1 vssd1 vccd1 vccd1 net63 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_130_907 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_935 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_255 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold803 team_03_WB.instance_to_wrap.core.register_file.registers_state\[786\] vssd1
+ vssd1 vccd1 vccd1 net2296 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_283 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold814 team_03_WB.instance_to_wrap.core.register_file.registers_state\[449\] vssd1
+ vssd1 vccd1 vccd1 net2307 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_732 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput74 wbs_adr_i[16] vssd1 vssd1 vccd1 vccd1 net74 sky130_fd_sc_hd__clkbuf_1
Xinput85 wbs_adr_i[26] vssd1 vssd1 vccd1 vccd1 net85 sky130_fd_sc_hd__clkbuf_1
Xhold825 team_03_WB.instance_to_wrap.core.register_file.registers_state\[867\] vssd1
+ vssd1 vccd1 vccd1 net2318 sky130_fd_sc_hd__dlygate4sd3_1
X_15080__1466 vssd1 vssd1 vccd1 vccd1 _15080__1466/HI net1466 sky130_fd_sc_hd__conb_1
XANTENNA__10746__B1 net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput96 wbs_adr_i[7] vssd1 vssd1 vccd1 vccd1 net96 sky130_fd_sc_hd__clkbuf_1
Xhold836 team_03_WB.instance_to_wrap.core.register_file.registers_state\[487\] vssd1
+ vssd1 vccd1 vccd1 net2329 sky130_fd_sc_hd__dlygate4sd3_1
Xhold847 team_03_WB.instance_to_wrap.core.register_file.registers_state\[329\] vssd1
+ vssd1 vccd1 vccd1 net2340 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_90_2221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_620 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_776 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_2232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold858 team_03_WB.instance_to_wrap.core.register_file.registers_state\[379\] vssd1
+ vssd1 vccd1 vccd1 net2351 sky130_fd_sc_hd__dlygate4sd3_1
X_09981_ _05852_ _05858_ _05082_ vssd1 vssd1 vccd1 vccd1 _05891_ sky130_fd_sc_hd__or3b_1
Xhold869 team_03_WB.instance_to_wrap.core.register_file.registers_state\[579\] vssd1
+ vssd1 vccd1 vccd1 net2362 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09039__S0 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08932_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[427\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[395\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[299\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[267\]
+ net977 net1071 vssd1 vssd1 vccd1 vccd1 _04874_ sky130_fd_sc_hd__mux4_1
XFILLER_0_122_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08167__A1 net1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10989__D net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08863_ net1067 _04801_ _04804_ vssd1 vssd1 vccd1 vccd1 _04805_ sky130_fd_sc_hd__a21o_1
XANTENNA__08262__S1 net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07914__A1 net1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07814_ net718 _03739_ _03748_ _03755_ vssd1 vssd1 vccd1 vccd1 _03756_ sky130_fd_sc_hd__a2bb2o_4
X_08794_ net1050 team_03_WB.instance_to_wrap.core.register_file.registers_state\[706\]
+ net1002 team_03_WB.instance_to_wrap.core.register_file.registers_state\[738\] net925
+ vssd1 vssd1 vccd1 vccd1 _04736_ sky130_fd_sc_hd__a221o_1
XFILLER_0_74_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09116__B1 net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_88_2183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07745_ net731 _03683_ _03684_ _03685_ _03686_ vssd1 vssd1 vccd1 vccd1 _03687_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_88_2194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07127__C1 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout360_A _06817_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout458_A net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09204__Y _05146_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07678__B1 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11474__B2 net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07676_ net1161 _03617_ vssd1 vssd1 vccd1 vccd1 _03618_ sky130_fd_sc_hd__or2_1
XFILLER_0_79_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_45_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09415_ _04416_ _04533_ net548 vssd1 vssd1 vccd1 vccd1 _05357_ sky130_fd_sc_hd__mux2_1
XANTENNA__08475__C _04415_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_366 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12018__A3 net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout625_A net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1367_A net1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09346_ _04148_ _05287_ vssd1 vssd1 vccd1 vccd1 _05288_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_62_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08627__C1 net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_134_3125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_134_3136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09277_ _03759_ _05218_ vssd1 vssd1 vccd1 vccd1 _05219_ sky130_fd_sc_hd__xor2_1
XANTENNA_fanout413_X net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_786 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11402__S net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1155_X net1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08228_ _04166_ _04169_ net1081 vssd1 vssd1 vccd1 vccd1 _04170_ sky130_fd_sc_hd__a21o_1
XFILLER_0_172_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_222 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_151_3472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout994_A _04086_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_151_3483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08159_ net1061 _04098_ _04099_ vssd1 vssd1 vccd1 vccd1 _04101_ sky130_fd_sc_hd__or3_1
XANTENNA__09052__C1 net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10737__B1 net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11170_ net710 _06503_ net694 vssd1 vssd1 vccd1 vccd1 _06664_ sky130_fd_sc_hd__or3_1
XANTENNA_fanout782_X net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10121_ _05962_ vssd1 vssd1 vccd1 vccd1 _05963_ sky130_fd_sc_hd__inv_2
XFILLER_0_100_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10542__A net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10052_ net4 net1036 net909 team_03_WB.instance_to_wrap.CPU_DAT_O\[11\] vssd1 vssd1
+ vccd1 vccd1 _02679_ sky130_fd_sc_hd__o22a_1
XANTENNA__11357__B _06468_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11701__A2 net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14860_ clknet_leaf_57_wb_clk_i net1903 _01225_ vssd1 vssd1 vccd1 vccd1 net116 sky130_fd_sc_hd__dfrtp_1
X_13811_ clknet_leaf_109_wb_clk_i _01575_ _00176_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[165\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input19_A DAT_I[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14791_ clknet_leaf_90_wb_clk_i _02555_ _01156_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_I\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_106_2548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11373__A net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_27_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13742_ clknet_leaf_131_wb_clk_i _01506_ _00107_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[96\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_158_3615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11465__B2 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10954_ net834 _06536_ vssd1 vssd1 vccd1 vccd1 _06537_ sky130_fd_sc_hd__and2_1
XFILLER_0_97_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_787 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_158_3626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_123_2895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13673_ clknet_leaf_77_wb_clk_i _01437_ _00038_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_10885_ team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[16\] net305 vssd1
+ vssd1 vccd1 vccd1 _06480_ sky130_fd_sc_hd__and2_1
XFILLER_0_39_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12624_ net1401 vssd1 vssd1 vccd1 vccd1 _00388_ sky130_fd_sc_hd__inv_2
XANTENNA__08618__C1 net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11768__A2 net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09497__B net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12555_ net1288 vssd1 vssd1 vccd1 vccd1 _00319_ sky130_fd_sc_hd__inv_2
XANTENNA__08094__B1 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09830__A1 net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11312__S net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11506_ _06624_ net2333 net390 vssd1 vssd1 vccd1 vccd1 _02000_ sky130_fd_sc_hd__mux2_1
XANTENNA__10440__A2 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07841__B1 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12486_ net1293 vssd1 vssd1 vccd1 vccd1 _00250_ sky130_fd_sc_hd__inv_2
XFILLER_0_112_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14225_ clknet_leaf_139_wb_clk_i _01989_ _00590_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[579\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09189__A3 _04565_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_789 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11437_ net2449 net392 _06758_ net492 vssd1 vssd1 vccd1 vccd1 _02049_ sky130_fd_sc_hd__a22o_1
XFILLER_0_80_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_58 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08397__A1 net1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14156_ clknet_leaf_20_wb_clk_i _01920_ _00521_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[510\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06930__A net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11368_ net504 net632 _06736_ net402 net1768 vssd1 vssd1 vccd1 vccd1 _02096_ sky130_fd_sc_hd__a32o_1
XFILLER_0_81_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14920__Q team_03_WB.instance_to_wrap.CPU_DAT_O\[7\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_13107_ net1265 vssd1 vssd1 vccd1 vccd1 _00871_ sky130_fd_sc_hd__inv_2
X_10319_ net282 _06159_ net678 vssd1 vssd1 vccd1 vccd1 _06160_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_0_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10452__A _05925_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14087_ clknet_leaf_109_wb_clk_i _01851_ _00452_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[441\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08149__A1 net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11299_ net1042 _06449_ net650 _06463_ vssd1 vssd1 vccd1 vccd1 _06717_ sky130_fd_sc_hd__or4_4
XANTENNA__11267__B net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13038_ net1305 vssd1 vssd1 vccd1 vccd1 _00802_ sky130_fd_sc_hd__inv_2
XANTENNA__09897__A1 net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11153__B1 net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1150 net1151 vssd1 vssd1 vccd1 vccd1 net1150 sky130_fd_sc_hd__buf_4
XANTENNA__11982__S net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1161 net1169 vssd1 vssd1 vccd1 vccd1 net1161 sky130_fd_sc_hd__buf_4
Xfanout1172 net1174 vssd1 vssd1 vccd1 vccd1 net1172 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10900__B1 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1183 net1190 vssd1 vssd1 vccd1 vccd1 net1183 sky130_fd_sc_hd__buf_2
Xfanout1194 net1195 vssd1 vssd1 vccd1 vccd1 net1194 sky130_fd_sc_hd__buf_2
XANTENNA__07761__A net1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09649__A1 _03428_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10598__S net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14989_ clknet_leaf_66_wb_clk_i net37 _01354_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07109__C1 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11283__A net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11456__A1 net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07530_ net1103 team_03_WB.instance_to_wrap.core.register_file.registers_state\[38\]
+ net899 vssd1 vssd1 vccd1 vccd1 _03472_ sky130_fd_sc_hd__or3_1
XFILLER_0_152_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_798 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07755__S0 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07461_ net1183 team_03_WB.instance_to_wrap.core.register_file.registers_state\[469\]
+ net769 team_03_WB.instance_to_wrap.core.register_file.registers_state\[501\] net1152
+ vssd1 vssd1 vccd1 vccd1 _03403_ sky130_fd_sc_hd__o221a_1
XANTENNA__09959__Y _05884_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_83_2080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_2091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09200_ _02954_ _05107_ _05141_ vssd1 vssd1 vccd1 vccd1 _05142_ sky130_fd_sc_hd__a21oi_4
X_07392_ net1082 team_03_WB.instance_to_wrap.core.register_file.registers_state\[959\]
+ net888 vssd1 vssd1 vccd1 vccd1 _03334_ sky130_fd_sc_hd__or3_1
XFILLER_0_173_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09131_ net583 _02953_ net580 vssd1 vssd1 vccd1 vccd1 _05073_ sky130_fd_sc_hd__and3_2
XTAP_TAPCELL_ROW_40_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08085__B1 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11222__S net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09062_ net921 _05003_ _05002_ net1219 vssd1 vssd1 vccd1 vccd1 _05004_ sky130_fd_sc_hd__a211o_1
XFILLER_0_142_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_96_wb_clk_i clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_96_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_5_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_7_Left_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08013_ net1177 team_03_WB.instance_to_wrap.core.register_file.registers_state\[593\]
+ net765 team_03_WB.instance_to_wrap.core.register_file.registers_state\[625\] net727
+ vssd1 vssd1 vccd1 vccd1 _03955_ sky130_fd_sc_hd__o221a_1
XFILLER_0_8_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09034__C1 net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold600 team_03_WB.instance_to_wrap.core.register_file.registers_state\[566\] vssd1
+ vssd1 vccd1 vccd1 net2093 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12842__A net1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold611 team_03_WB.instance_to_wrap.core.register_file.registers_state\[892\] vssd1
+ vssd1 vccd1 vccd1 net2104 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_25_wb_clk_i clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_25_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__10065__C net1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08388__A1 net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold622 team_03_WB.instance_to_wrap.core.register_file.registers_state\[243\] vssd1
+ vssd1 vccd1 vccd1 net2115 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold633 team_03_WB.instance_to_wrap.core.register_file.registers_state\[189\] vssd1
+ vssd1 vccd1 vccd1 net2126 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold644 team_03_WB.instance_to_wrap.core.register_file.registers_state\[684\] vssd1
+ vssd1 vccd1 vccd1 net2137 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06840__A team_03_WB.instance_to_wrap.core.decoder.inst\[26\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold655 team_03_WB.instance_to_wrap.core.register_file.registers_state\[748\] vssd1
+ vssd1 vccd1 vccd1 net2148 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11392__B1 net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold666 team_03_WB.instance_to_wrap.core.register_file.registers_state\[190\] vssd1
+ vssd1 vccd1 vccd1 net2159 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold677 team_03_WB.instance_to_wrap.core.register_file.registers_state\[771\] vssd1
+ vssd1 vccd1 vccd1 net2170 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_38_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07060__A1 net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold688 team_03_WB.instance_to_wrap.core.register_file.registers_state\[737\] vssd1
+ vssd1 vccd1 vccd1 net2181 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11458__A net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12053__S net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09964_ _05886_ net1833 net291 vssd1 vssd1 vccd1 vccd1 _02745_ sky130_fd_sc_hd__mux2_1
Xhold699 team_03_WB.instance_to_wrap.core.register_file.registers_state\[381\] vssd1
+ vssd1 vccd1 vccd1 net2192 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1115_A net1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08915_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[1004\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[972\]
+ net979 vssd1 vssd1 vccd1 vccd1 _04857_ sky130_fd_sc_hd__mux2_1
XANTENNA__07374__C net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09895_ _04031_ _04323_ net536 vssd1 vssd1 vccd1 vccd1 _05837_ sky130_fd_sc_hd__or3_1
XANTENNA__10498__A2 net1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08846_ net1056 team_03_WB.instance_to_wrap.core.register_file.registers_state\[320\]
+ net1009 team_03_WB.instance_to_wrap.core.register_file.registers_state\[352\] net1216
+ vssd1 vssd1 vccd1 vccd1 _04788_ sky130_fd_sc_hd__a221o_1
XANTENNA__07899__B1 _02872_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08560__A1 net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout742_A net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08777_ net1050 team_03_WB.instance_to_wrap.core.register_file.registers_state\[194\]
+ net1003 team_03_WB.instance_to_wrap.core.register_file.registers_state\[226\] net924
+ vssd1 vssd1 vccd1 vccd1 _04719_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout363_X net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07728_ net1197 team_03_WB.instance_to_wrap.core.register_file.registers_state\[845\]
+ net786 team_03_WB.instance_to_wrap.core.register_file.registers_state\[877\] net1134
+ vssd1 vssd1 vccd1 vccd1 _03670_ sky130_fd_sc_hd__o221a_1
XANTENNA__11447__B2 net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08312__A1 net1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11998__A2 net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout530_X net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07659_ team_03_WB.instance_to_wrap.core.decoder.inst\[14\] net1015 _03107_ vssd1
+ vssd1 vccd1 vccd1 _03601_ sky130_fd_sc_hd__a21o_2
XANTENNA__07520__C1 net1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11343__D net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_2445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_314 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout628_X net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_2456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09598__A _05539_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10670_ _05583_ _06311_ vssd1 vssd1 vccd1 vccd1 _06312_ sky130_fd_sc_hd__nor2_1
XFILLER_0_36_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_153_3512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_153_3523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09902__D_N _05583_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09329_ _05246_ _05250_ _05269_ _05244_ _05241_ vssd1 vssd1 vccd1 vccd1 _05271_ sky130_fd_sc_hd__a311o_2
XTAP_TAPCELL_ROW_11_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09812__A1 _03024_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_168_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12340_ net1303 vssd1 vssd1 vccd1 vccd1 _00104_ sky130_fd_sc_hd__inv_2
XFILLER_0_62_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07823__B1 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_170_3870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout997_X net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10971__S net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12271_ net1394 vssd1 vssd1 vccd1 vccd1 _00035_ sky130_fd_sc_hd__inv_2
XFILLER_0_160_372 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12752__A net1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_33_wb_clk_i_A clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09576__B1 _05516_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14010_ clknet_leaf_145_wb_clk_i _01774_ _00375_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[364\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_79_1993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11222_ net270 net2303 net486 vssd1 vssd1 vccd1 vccd1 _02188_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_951 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09671__S0 net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11153_ net490 net646 _06653_ net412 net1972 vssd1 vssd1 vccd1 vccd1 _02228_ sky130_fd_sc_hd__a32o_1
X_10104_ _02811_ _02816_ _02830_ _02833_ vssd1 vssd1 vccd1 vccd1 _05948_ sky130_fd_sc_hd__a211o_4
XFILLER_0_101_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11084_ net832 net275 vssd1 vssd1 vccd1 vccd1 _06620_ sky130_fd_sc_hd__and2_2
XANTENNA__11135__B1 net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14912_ clknet_leaf_55_wb_clk_i _00006_ _01277_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.ru.state\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_10035_ net22 net1037 net909 net2391 vssd1 vssd1 vccd1 vccd1 _02696_ sky130_fd_sc_hd__o22a_1
XANTENNA__10489__A2 net1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08551__A1 net1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14843_ clknet_leaf_81_wb_clk_i net1639 _01208_ vssd1 vssd1 vccd1 vccd1 net129 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_125_2946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output125_A net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06909__B net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11307__S net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11534__C net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14774_ clknet_leaf_103_wb_clk_i _02538_ _01139_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_I\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_11986_ net274 net2575 net443 vssd1 vssd1 vccd1 vccd1 _01558_ sky130_fd_sc_hd__mux2_1
XANTENNA__11989__A2 net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13725_ clknet_leaf_29_wb_clk_i _01489_ _00090_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[79\]
+ sky130_fd_sc_hd__dfrtp_1
X_10937_ net688 _06521_ _06522_ _06520_ vssd1 vssd1 vccd1 vccd1 _06523_ sky130_fd_sc_hd__o31a_4
XFILLER_0_86_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_908 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12927__A net1347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13656_ clknet_leaf_172_wb_clk_i _01420_ _00021_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_155_133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10868_ team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[19\] net307 net685 vssd1
+ vssd1 vccd1 vccd1 _06466_ sky130_fd_sc_hd__a21o_1
XFILLER_0_128_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06925__A net1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_72_wb_clk_i_A clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_27_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09301__A _03489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14915__Q team_03_WB.instance_to_wrap.CPU_DAT_O\[2\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_112_1076 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12607_ net1285 vssd1 vssd1 vccd1 vccd1 _00371_ sky130_fd_sc_hd__inv_2
XFILLER_0_155_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13587_ net1345 vssd1 vssd1 vccd1 vccd1 _01351_ sky130_fd_sc_hd__inv_2
XANTENNA__10949__A0 _06532_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10799_ team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[30\] net305 _06407_ net691
+ vssd1 vssd1 vccd1 vccd1 _06408_ sky130_fd_sc_hd__o211a_1
XFILLER_0_54_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12538_ net1372 vssd1 vssd1 vccd1 vccd1 _00302_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11977__S net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12469_ net1290 vssd1 vssd1 vccd1 vccd1 _00233_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09955__B net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09567__B1 _04816_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14208_ clknet_leaf_190_wb_clk_i _01972_ _00573_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[562\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08351__S net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11374__B1 net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14139_ clknet_leaf_134_wb_clk_i _01903_ _00504_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[493\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10182__A team_03_WB.instance_to_wrap.core.decoder.inst\[28\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout409 _06684_ vssd1 vssd1 vccd1 vccd1 net409 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09971__A _03205_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06961_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[421\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[389\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[293\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[261\]
+ net787 net1135 vssd1 vssd1 vccd1 vccd1 _02903_ sky130_fd_sc_hd__mux4_1
X_08700_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[424\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[392\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[296\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[264\]
+ net975 net1075 vssd1 vssd1 vccd1 vccd1 _04642_ sky130_fd_sc_hd__mux4_1
XFILLER_0_20_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09680_ _05621_ _05616_ _05620_ vssd1 vssd1 vccd1 vccd1 _05622_ sky130_fd_sc_hd__or3b_2
XTAP_TAPCELL_ROW_33_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06892_ _02816_ _02830_ _02833_ vssd1 vssd1 vccd1 vccd1 _02834_ sky130_fd_sc_hd__nor3_1
XANTENNA__08542__A1 net1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_143_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_143_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_08631_ net863 _04571_ _04572_ _04570_ vssd1 vssd1 vccd1 vccd1 _04573_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_85_2120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11217__S net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08562_ _04503_ vssd1 vssd1 vccd1 vccd1 _04504_ sky130_fd_sc_hd__inv_2
XANTENNA__08874__X _04816_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_2039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07513_ net1135 _03453_ net1168 vssd1 vssd1 vccd1 vccd1 _03455_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_162_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08493_ net1242 team_03_WB.instance_to_wrap.core.register_file.registers_state\[219\]
+ net985 team_03_WB.instance_to_wrap.core.register_file.registers_state\[251\] net945
+ vssd1 vssd1 vccd1 vccd1 _04435_ sky130_fd_sc_hd__o221a_1
XFILLER_0_146_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07444_ net1161 _03385_ vssd1 vssd1 vccd1 vccd1 _03386_ sky130_fd_sc_hd__or2_1
XFILLER_0_18_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09211__A net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10357__A net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07375_ net1084 net889 team_03_WB.instance_to_wrap.core.register_file.registers_state\[159\]
+ vssd1 vssd1 vccd1 vccd1 _03317_ sky130_fd_sc_hd__o21a_1
XFILLER_0_88_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12048__S net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout323_A _06811_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1065_A net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09114_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[942\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[910\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[814\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[782\]
+ net978 net1075 vssd1 vssd1 vccd1 vccd1 _05056_ sky130_fd_sc_hd__mux4_1
XFILLER_0_5_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_687 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07281__A1 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10955__A3 net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09045_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[15\] net998
+ net921 _04986_ vssd1 vssd1 vccd1 vccd1 _04987_ sky130_fd_sc_hd__o211a_1
XFILLER_0_103_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1232_A net1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_748 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold430 team_03_WB.instance_to_wrap.core.register_file.registers_state\[241\] vssd1
+ vssd1 vccd1 vccd1 net1923 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold441 team_03_WB.instance_to_wrap.core.register_file.registers_state\[445\] vssd1
+ vssd1 vccd1 vccd1 net1934 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout692_A net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold452 team_03_WB.instance_to_wrap.core.register_file.registers_state\[567\] vssd1
+ vssd1 vccd1 vccd1 net1945 sky130_fd_sc_hd__dlygate4sd3_1
Xhold463 team_03_WB.instance_to_wrap.core.register_file.registers_state\[354\] vssd1
+ vssd1 vccd1 vccd1 net1956 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11188__A net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold474 net155 vssd1 vssd1 vccd1 vccd1 net1967 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10092__A _05563_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08230__B1 net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_3024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1020_X net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold485 team_03_WB.instance_to_wrap.core.register_file.registers_state\[110\] vssd1
+ vssd1 vccd1 vccd1 net1978 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1118_X net1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold496 team_03_WB.instance_to_wrap.core.register_file.registers_state\[385\] vssd1
+ vssd1 vccd1 vccd1 net1989 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_117_wb_clk_i_A clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout910 _05907_ vssd1 vssd1 vccd1 vccd1 net910 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_74_1890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout921 net922 vssd1 vssd1 vccd1 vccd1 net921 sky130_fd_sc_hd__buf_4
X_09947_ _03389_ net662 vssd1 vssd1 vccd1 vccd1 _05878_ sky130_fd_sc_hd__nor2_1
Xfanout932 _04088_ vssd1 vssd1 vccd1 vccd1 net932 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout480_X net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout943 net948 vssd1 vssd1 vccd1 vccd1 net943 sky130_fd_sc_hd__buf_2
Xfanout954 net955 vssd1 vssd1 vccd1 vccd1 net954 sky130_fd_sc_hd__buf_2
XANTENNA_fanout578_X net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout957_A net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_146_3371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout965 net974 vssd1 vssd1 vccd1 vccd1 net965 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_146_3382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout976 net978 vssd1 vssd1 vccd1 vccd1 net976 sky130_fd_sc_hd__clkbuf_4
X_09878_ net351 _05404_ _05815_ _05817_ _05819_ vssd1 vssd1 vccd1 vccd1 _05820_ sky130_fd_sc_hd__a2111o_1
Xfanout987 net988 vssd1 vssd1 vccd1 vccd1 net987 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_5_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1130 team_03_WB.instance_to_wrap.core.register_file.registers_state\[726\] vssd1
+ vssd1 vccd1 vccd1 net2623 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout998 net999 vssd1 vssd1 vccd1 vccd1 net998 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_5_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1141 team_03_WB.instance_to_wrap.core.register_file.registers_state\[156\] vssd1
+ vssd1 vccd1 vccd1 net2634 sky130_fd_sc_hd__dlygate4sd3_1
X_08829_ _04080_ _04770_ vssd1 vssd1 vccd1 vccd1 _04771_ sky130_fd_sc_hd__nor2_1
Xhold1152 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[15\] vssd1 vssd1
+ vccd1 vccd1 net2645 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1163 team_03_WB.instance_to_wrap.core.register_file.registers_state\[320\] vssd1
+ vssd1 vccd1 vccd1 net2656 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_203 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout745_X net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1174 team_03_WB.instance_to_wrap.core.register_file.registers_state\[666\] vssd1
+ vssd1 vccd1 vccd1 net2667 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1185 team_03_WB.instance_to_wrap.core.register_file.registers_state\[80\] vssd1
+ vssd1 vccd1 vccd1 net2678 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1196 team_03_WB.instance_to_wrap.core.register_file.registers_state\[68\] vssd1
+ vssd1 vccd1 vccd1 net2689 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_174_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11840_ _06678_ net471 net325 net1914 vssd1 vssd1 vccd1 vccd1 _01699_ sky130_fd_sc_hd__a22o_1
XANTENNA__10891__A2 net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_2832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11771_ net656 _06604_ net473 net333 net2171 vssd1 vssd1 vccd1 vccd1 _01766_ sky130_fd_sc_hd__a32o_1
XFILLER_0_166_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_120_2843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07639__A3 net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13510_ net1322 vssd1 vssd1 vccd1 vccd1 _01274_ sky130_fd_sc_hd__inv_2
X_10722_ net1564 net527 net522 _06352_ vssd1 vssd1 vccd1 vccd1 _02454_ sky130_fd_sc_hd__a22o_1
XFILLER_0_138_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_165_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09685__A1_N net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14490_ clknet_leaf_148_wb_clk_i _02254_ _00855_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[844\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08436__S net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_172_3910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13441_ net1423 vssd1 vssd1 vccd1 vccd1 _01205_ sky130_fd_sc_hd__inv_2
X_10653_ net1251 team_03_WB.instance_to_wrap.CPU_DAT_O\[8\] net847 vssd1 vssd1 vccd1
+ vccd1 _02475_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_153_659 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input86_A wbs_adr_i[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_687 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13372_ net1415 vssd1 vssd1 vccd1 vccd1 _01136_ sky130_fd_sc_hd__inv_2
XFILLER_0_152_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10584_ net1713 net532 net599 _02888_ vssd1 vssd1 vccd1 vccd1 _02539_ sky130_fd_sc_hd__a22o_1
XFILLER_0_24_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkload19 clknet_leaf_7_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload19/Y sky130_fd_sc_hd__bufinv_16
X_15111_ net913 vssd1 vssd1 vccd1 vccd1 net245 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_140_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11797__S net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_156_wb_clk_i_A clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_2_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12323_ net1371 vssd1 vssd1 vccd1 vccd1 _00087_ sky130_fd_sc_hd__inv_2
XANTENNA__07847__Y _03789_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_2794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09549__B1 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15042_ clknet_leaf_87_wb_clk_i _02762_ _01407_ vssd1 vssd1 vccd1 vccd1 net198 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_160_180 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12254_ net1392 vssd1 vssd1 vccd1 vccd1 _00018_ sky130_fd_sc_hd__inv_2
XANTENNA__11356__B1 net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11205_ _06430_ net2420 net489 vssd1 vssd1 vccd1 vccd1 _02203_ sky130_fd_sc_hd__mux2_1
XANTENNA__07024__A1 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12185_ net1541 vssd1 vssd1 vccd1 vccd1 _02368_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_102_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11136_ net277 net657 net707 net699 vssd1 vssd1 vccd1 vccd1 _06644_ sky130_fd_sc_hd__and4_1
XPHY_EDGE_ROW_79_Left_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11067_ _06611_ net2595 net416 vssd1 vssd1 vccd1 vccd1 _02272_ sky130_fd_sc_hd__mux2_1
XANTENNA__08524__A1 net1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10018_ _05892_ _05893_ _05894_ _05895_ vssd1 vssd1 vccd1 vccd1 _05896_ sky130_fd_sc_hd__or4_1
XANTENNA__07742__C net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14826_ clknet_leaf_104_wb_clk_i net1657 _01191_ vssd1 vssd1 vccd1 vccd1 net146 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_99_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14757_ clknet_leaf_53_wb_clk_i _02521_ _01122_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12084__A1 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12657__A net1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11969_ net639 _06746_ net473 net366 net2378 vssd1 vssd1 vccd1 vccd1 _01574_ sky130_fd_sc_hd__a32o_1
XANTENNA__11561__A net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13708_ clknet_leaf_18_wb_clk_i _01472_ _00073_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[62\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_88_Left_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11831__A1 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14688_ clknet_leaf_57_wb_clk_i _02452_ _01053_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.ADR_I\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_157_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_678 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13639_ net1434 vssd1 vssd1 vccd1 vccd1 _01403_ sky130_fd_sc_hd__inv_2
XFILLER_0_132_67 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10177__A _04922_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_486 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07160_ net819 _03091_ _03101_ vssd1 vssd1 vccd1 vccd1 _03102_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_55_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_171_456 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11595__A0 net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_350 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07091_ net1102 team_03_WB.instance_to_wrap.core.register_file.registers_state\[705\]
+ vssd1 vssd1 vccd1 vccd1 _03033_ sky130_fd_sc_hd__and2_1
XFILLER_0_48_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11500__S net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_11__f_wb_clk_i_A clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08438__S1 net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08212__B1 net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_97_Left_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_35_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11898__A1 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09801_ _03490_ _04592_ net667 _05742_ vssd1 vssd1 vccd1 vccd1 _05743_ sky130_fd_sc_hd__a22o_1
XANTENNA__09960__A0 _05884_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_598 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07993_ net1203 team_03_WB.instance_to_wrap.core.register_file.registers_state\[592\]
+ net786 team_03_WB.instance_to_wrap.core.register_file.registers_state\[624\] net735
+ vssd1 vssd1 vccd1 vccd1 _03935_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_52_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09732_ _02953_ net573 _05442_ net352 vssd1 vssd1 vccd1 vccd1 _05674_ sky130_fd_sc_hd__a31o_1
X_06944_ _02882_ _02883_ _02885_ _02884_ net750 net813 vssd1 vssd1 vccd1 vccd1 _02886_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_2_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09663_ net538 _05604_ vssd1 vssd1 vccd1 vccd1 _05605_ sky130_fd_sc_hd__nand2_1
X_06875_ _02794_ team_03_WB.instance_to_wrap.core.control_logic.instruction\[3\] _02805_
+ team_03_WB.instance_to_wrap.core.control_logic.instruction\[5\] team_03_WB.instance_to_wrap.core.control_logic.instruction\[6\]
+ vssd1 vssd1 vccd1 vccd1 _02817_ sky130_fd_sc_hd__a2111oi_2
XANTENNA_fanout273_A _06473_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08614_ net1058 team_03_WB.instance_to_wrap.core.register_file.registers_state\[69\]
+ net1012 team_03_WB.instance_to_wrap.core.register_file.registers_state\[101\] net947
+ vssd1 vssd1 vccd1 vccd1 _04556_ sky130_fd_sc_hd__a221o_1
XFILLER_0_96_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09594_ net569 _05407_ vssd1 vssd1 vccd1 vccd1 _05536_ sky130_fd_sc_hd__nand2_1
X_08545_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[574\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[542\]
+ net955 vssd1 vssd1 vccd1 vccd1 _04487_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout440_A _06819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1182_A net1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout538_A net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11471__A net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07177__S1 net1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11822__A1 net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08476_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[571\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[539\]
+ net987 vssd1 vssd1 vccd1 vccd1 _04418_ sky130_fd_sc_hd__mux2_1
XFILLER_0_147_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11190__B net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07427_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[916\] net795
+ net1014 _03368_ vssd1 vssd1 vccd1 vccd1 _03369_ sky130_fd_sc_hd__o211a_1
XFILLER_0_174_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout326_X net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout705_A net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_40_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_40_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_119_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1068_X net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07358_ net1083 team_03_WB.instance_to_wrap.core.register_file.registers_state\[700\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[668\] net792 net739
+ vssd1 vssd1 vccd1 vccd1 _03300_ sky130_fd_sc_hd__o221a_1
XFILLER_0_73_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11586__A0 net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_98_2388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_2399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10928__A3 net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08451__B1 net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11050__A2 net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07289_ net1201 team_03_WB.instance_to_wrap.core.register_file.registers_state\[201\]
+ net788 team_03_WB.instance_to_wrap.core.register_file.registers_state\[233\] net750
+ vssd1 vssd1 vccd1 vccd1 _03231_ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout1235_X net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11410__S net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_76_1930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09028_ _04964_ _04969_ net873 vssd1 vssd1 vccd1 vccd1 _04970_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_76_1941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07827__C net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11338__B1 net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout695_X net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_148_3411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold260 net191 vssd1 vssd1 vccd1 vccd1 net1753 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_148_3422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11889__A1 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1402_X net1402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold271 team_03_WB.instance_to_wrap.core.register_file.registers_state\[992\] vssd1
+ vssd1 vccd1 vccd1 net1764 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11349__C _06438_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_2691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10010__A0 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold282 team_03_WB.instance_to_wrap.core.register_file.registers_state\[308\] vssd1
+ vssd1 vccd1 vccd1 net1775 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_72_1849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold293 net217 vssd1 vssd1 vccd1 vccd1 net1786 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout862_X net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout740 net742 vssd1 vssd1 vccd1 vccd1 net740 sky130_fd_sc_hd__buf_4
Xfanout751 net754 vssd1 vssd1 vccd1 vccd1 net751 sky130_fd_sc_hd__buf_2
XANTENNA__15118__A net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout762 net763 vssd1 vssd1 vccd1 vccd1 net762 sky130_fd_sc_hd__clkbuf_4
X_13990_ clknet_leaf_72_wb_clk_i _01754_ _00355_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[344\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout773 _02851_ vssd1 vssd1 vccd1 vccd1 net773 sky130_fd_sc_hd__clkbuf_4
Xfanout784 net790 vssd1 vssd1 vccd1 vccd1 net784 sky130_fd_sc_hd__buf_2
XFILLER_0_137_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout795 _02850_ vssd1 vssd1 vccd1 vccd1 net795 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11365__B net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12941_ net1311 vssd1 vssd1 vccd1 vccd1 _00705_ sky130_fd_sc_hd__inv_2
XFILLER_0_99_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_161_3677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_161_3688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12872_ net1295 vssd1 vssd1 vccd1 vccd1 _00636_ sky130_fd_sc_hd__inv_2
X_14611_ clknet_leaf_100_wb_clk_i _02375_ _00976_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[965\]
+ sky130_fd_sc_hd__dfstp_1
X_11823_ net646 _06653_ net451 net323 net1757 vssd1 vssd1 vccd1 vccd1 _01716_ sky130_fd_sc_hd__a32o_1
XFILLER_0_139_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_554 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11381__A net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14542_ clknet_leaf_125_wb_clk_i _02306_ _00907_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[896\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11813__A1 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11754_ net652 _06579_ net458 net332 net2293 vssd1 vssd1 vccd1 vccd1 _01783_ sky130_fd_sc_hd__a32o_1
XANTENNA__09482__A2 _04503_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_7__f_wb_clk_i_A clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10705_ team_03_WB.instance_to_wrap.core.pc.current_pc\[26\] _06315_ vssd1 vssd1
+ vccd1 vccd1 _06342_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_153_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14473_ clknet_leaf_76_wb_clk_i _02237_ _00838_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[827\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_626 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11685_ _06727_ net381 net339 net1860 vssd1 vssd1 vccd1 vccd1 _01849_ sky130_fd_sc_hd__a22o_1
X_13424_ net1421 vssd1 vssd1 vccd1 vccd1 _01188_ sky130_fd_sc_hd__inv_2
X_10636_ team_03_WB.instance_to_wrap.core.decoder.inst\[25\] net1785 net845 vssd1
+ vssd1 vccd1 vccd1 _02492_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11577__A0 net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload108 clknet_leaf_156_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload108/Y sky130_fd_sc_hd__clkinv_1
XFILLER_0_63_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_590 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07245__A1 net1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkload119 clknet_leaf_163_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload119/Y sky130_fd_sc_hd__clkinv_8
X_13355_ net1315 vssd1 vssd1 vccd1 vccd1 _01119_ sky130_fd_sc_hd__inv_2
X_10567_ net1670 net532 net599 _05877_ vssd1 vssd1 vccd1 vccd1 _02556_ sky130_fd_sc_hd__a22o_1
XANTENNA__09785__A3 _04820_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06922__B net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11320__S net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12306_ net1397 vssd1 vssd1 vccd1 vccd1 _00070_ sky130_fd_sc_hd__inv_2
X_13286_ net1343 vssd1 vssd1 vccd1 vccd1 _01050_ sky130_fd_sc_hd__inv_2
XANTENNA__11329__A0 net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10498_ net133 net1030 net907 net1612 vssd1 vssd1 vccd1 vccd1 _02611_ sky130_fd_sc_hd__a22o_1
X_15025_ clknet_leaf_130_wb_clk_i _02745_ _01390_ vssd1 vssd1 vccd1 vccd1 net181 sky130_fd_sc_hd__dfrtp_1
X_12237_ net1627 vssd1 vssd1 vccd1 vccd1 _01420_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__11259__C net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10001__A0 _05886_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08745__A1 net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12168_ net1522 vssd1 vssd1 vccd1 vccd1 _02385_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__10552__A1 net1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07953__C1 net1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11119_ _06633_ net2683 net418 vssd1 vssd1 vccd1 vccd1 _02242_ sky130_fd_sc_hd__mux2_1
XFILLER_0_127_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12099_ _06796_ net480 net442 net2099 vssd1 vssd1 vccd1 vccd1 _01448_ sky130_fd_sc_hd__a22o_1
XFILLER_0_127_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09026__A net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput6 DAT_I[13] vssd1 vssd1 vccd1 vccd1 net6 sky130_fd_sc_hd__buf_1
XANTENNA_clkbuf_3_4_0_wb_clk_i_X clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07705__C1 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11990__S net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14809_ clknet_leaf_104_wb_clk_i net1667 _01174_ vssd1 vssd1 vccd1 vccd1 net158 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_143_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_143_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11291__A net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08330_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[565\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[533\]
+ net972 vssd1 vssd1 vccd1 vccd1 _04272_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11804__A1 net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_99 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07484__A1 net1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08261_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[1010\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[978\]
+ net951 vssd1 vssd1 vccd1 vccd1 _04203_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09967__Y _05888_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11280__A2 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07212_ net1170 team_03_WB.instance_to_wrap.core.register_file.registers_state\[594\]
+ net756 team_03_WB.instance_to_wrap.core.register_file.registers_state\[626\] net725
+ vssd1 vssd1 vccd1 vccd1 _03154_ sky130_fd_sc_hd__o221a_1
XFILLER_0_172_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08192_ _04128_ _04133_ net872 vssd1 vssd1 vccd1 vccd1 _04134_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07143_ net1198 team_03_WB.instance_to_wrap.core.register_file.registers_state\[128\]
+ net885 net1155 vssd1 vssd1 vccd1 vccd1 _03085_ sky130_fd_sc_hd__o211a_1
XFILLER_0_42_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11230__S net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08984__A1 net1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07331__S1 net1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07074_ net1095 team_03_WB.instance_to_wrap.core.register_file.registers_state\[322\]
+ net796 team_03_WB.instance_to_wrap.core.register_file.registers_state\[354\] net1154
+ vssd1 vssd1 vccd1 vccd1 _03016_ sky130_fd_sc_hd__a221oi_1
XTAP_TAPCELL_ROW_93_2285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_2296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_7_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08197__C1 net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1028_A net1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_7_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08736__A1 net1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout390_A _06778_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout488_A _06680_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11740__B1 _06808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11466__A net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12061__S net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07976_ net1111 team_03_WB.instance_to_wrap.core.register_file.registers_state\[496\]
+ net901 _03917_ net1156 vssd1 vssd1 vccd1 vccd1 _03918_ sky130_fd_sc_hd__o311a_1
X_09715_ _04777_ _05650_ _05656_ vssd1 vssd1 vccd1 vccd1 _05657_ sky130_fd_sc_hd__a21oi_2
X_06927_ net1132 net1164 vssd1 vssd1 vccd1 vccd1 _02869_ sky130_fd_sc_hd__nor2_4
XANTENNA_fanout655_A net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout276_X net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1397_A net1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09646_ _03428_ _04295_ vssd1 vssd1 vccd1 vccd1 _05588_ sky130_fd_sc_hd__or2_1
X_06858_ team_03_WB.instance_to_wrap.core.control_logic.instruction\[3\] team_03_WB.instance_to_wrap.core.control_logic.instruction\[2\]
+ team_03_WB.instance_to_wrap.core.control_logic.instruction\[1\] team_03_WB.instance_to_wrap.core.control_logic.instruction\[0\]
+ vssd1 vssd1 vccd1 vccd1 _02800_ sky130_fd_sc_hd__nand4b_4
X_09577_ _05315_ _05431_ vssd1 vssd1 vccd1 vccd1 _05519_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12297__A net1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout443_X net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout822_A net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1185_X net1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10059__B1 net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11405__S net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08528_ net1227 team_03_WB.instance_to_wrap.core.register_file.registers_state\[479\]
+ net956 team_03_WB.instance_to_wrap.core.register_file.registers_state\[511\] net1210
+ vssd1 vssd1 vccd1 vccd1 _04470_ sky130_fd_sc_hd__o221a_1
XFILLER_0_65_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08267__A3 _04207_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07475__A1 net1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_167_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08459_ net850 _04400_ vssd1 vssd1 vccd1 vccd1 _04401_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_14_Right_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout708_X net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_163_743 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_516 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_899 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_3189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11470_ net491 net620 _06595_ net392 net2320 vssd1 vssd1 vccd1 vccd1 _02028_ sky130_fd_sc_hd__a32o_1
XFILLER_0_92_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_162_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_163_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10421_ _06012_ _06014_ vssd1 vssd1 vccd1 vccd1 _06243_ sky130_fd_sc_hd__nand2_1
XANTENNA__07227__A1 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11023__A2 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_2731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_2742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13140_ net1308 vssd1 vssd1 vccd1 vccd1 _00904_ sky130_fd_sc_hd__inv_2
X_10352_ team_03_WB.instance_to_wrap.core.pc.current_pc\[23\] _06147_ vssd1 vssd1
+ vccd1 vccd1 _06186_ sky130_fd_sc_hd__nor2_1
XFILLER_0_104_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13071_ net1338 vssd1 vssd1 vccd1 vccd1 _00835_ sky130_fd_sc_hd__inv_2
X_10283_ _05973_ _06124_ vssd1 vssd1 vccd1 vccd1 _06125_ sky130_fd_sc_hd__nand2_1
XANTENNA__12760__A net1376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08188__C1 net1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08727__A1 net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09545__S net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12022_ _06766_ net455 net359 net2186 vssd1 vssd1 vccd1 vccd1 _01523_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_163_3717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_1125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input49_A gpio_in[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_163_3728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10551__Y _06294_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_23_Right_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_4_10__f_wb_clk_i_X clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11731__B1 _06808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout570 net572 vssd1 vssd1 vccd1 vccd1 net570 sky130_fd_sc_hd__buf_2
Xfanout581 net582 vssd1 vssd1 vccd1 vccd1 net581 sky130_fd_sc_hd__buf_4
XANTENNA__11095__B net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13973_ clknet_leaf_129_wb_clk_i _01737_ _00338_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[327\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09152__A1 net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12924_ net1411 vssd1 vssd1 vccd1 vccd1 _00688_ sky130_fd_sc_hd__inv_2
XANTENNA__07702__A2 net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12855_ net1390 vssd1 vssd1 vccd1 vccd1 _00619_ sky130_fd_sc_hd__inv_2
XANTENNA__11315__S net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_559 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11806_ net2315 net263 net329 vssd1 vssd1 vccd1 vccd1 _01732_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12786_ net1397 vssd1 vssd1 vccd1 vccd1 _00550_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_32_Right_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07466__A1 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14525_ clknet_leaf_166_wb_clk_i _02289_ _00890_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[879\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_166_570 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11262__A2 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11737_ net2026 net269 net336 vssd1 vssd1 vccd1 vccd1 _01799_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12935__A net1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07561__S1 net1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14456_ clknet_leaf_5_wb_clk_i _02220_ _00821_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[810\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_142_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11668_ net2385 _06629_ net345 vssd1 vssd1 vccd1 vccd1 _01865_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13407_ net1322 vssd1 vssd1 vccd1 vccd1 _01171_ sky130_fd_sc_hd__inv_2
XANTENNA__14923__Q team_03_WB.instance_to_wrap.CPU_DAT_O\[10\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__07218__A1 net1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10619_ net1643 team_03_WB.instance_to_wrap.CPU_DAT_O\[10\] net841 vssd1 vssd1 vccd1
+ vccd1 _02509_ sky130_fd_sc_hd__mux2_1
XANTENNA__11014__A2 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14387_ clknet_leaf_106_wb_clk_i _02151_ _00752_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[741\]
+ sky130_fd_sc_hd__dfrtp_1
X_11599_ _06518_ net2249 net449 vssd1 vssd1 vccd1 vccd1 _01930_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07769__A2 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_180 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13338_ net1315 vssd1 vssd1 vccd1 vccd1 _01102_ sky130_fd_sc_hd__inv_2
XFILLER_0_11_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_1025 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10174__B net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06977__B1 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11970__B1 net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11985__S net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13269_ net1276 vssd1 vssd1 vccd1 vccd1 _01033_ sky130_fd_sc_hd__inv_2
XANTENNA__12670__A net1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09963__B net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_41_Right_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15008_ clknet_leaf_63_wb_clk_i net56 _01373_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10902__B net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11722__B1 _06808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07830_ net1175 team_03_WB.instance_to_wrap.core.register_file.registers_state\[490\]
+ net880 _03771_ vssd1 vssd1 vccd1 vccd1 _03772_ sky130_fd_sc_hd__a31o_1
XFILLER_0_47_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07761_ net1094 team_03_WB.instance_to_wrap.core.register_file.registers_state\[940\]
+ net897 vssd1 vssd1 vccd1 vccd1 _03703_ sky130_fd_sc_hd__or3_1
XANTENNA__11436__D net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09500_ _05441_ vssd1 vssd1 vccd1 vccd1 _05442_ sky130_fd_sc_hd__inv_2
XFILLER_0_91_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_155_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07692_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[798\] net793
+ _03633_ vssd1 vssd1 vccd1 vccd1 _03634_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_78_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07154__B1 net1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09431_ _05013_ _05070_ vssd1 vssd1 vccd1 vccd1 _05373_ sky130_fd_sc_hd__nor2_1
XFILLER_0_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_50_Right_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_1078 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09362_ _05283_ _05289_ vssd1 vssd1 vccd1 vccd1 _05304_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_47_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07004__A team_03_WB.instance_to_wrap.core.decoder.inst\[13\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08313_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[824\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[792\]
+ net972 vssd1 vssd1 vccd1 vccd1 _04255_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_170_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09293_ _05222_ _05233_ _05234_ _05220_ vssd1 vssd1 vccd1 vccd1 _05235_ sky130_fd_sc_hd__o211a_1
XANTENNA__08654__B1 net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10068__C team_03_WB.instance_to_wrap.core.decoder.inst\[12\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08244_ net854 _04184_ _04185_ vssd1 vssd1 vccd1 vccd1 _04186_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_43_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06843__A net1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07209__A1 net1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_95_2325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_2336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08175_ _04114_ _04116_ net1081 vssd1 vssd1 vccd1 vccd1 _04117_ sky130_fd_sc_hd__a21o_1
XANTENNA__12056__S net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout403_A _06718_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_6__f_wb_clk_i_X clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_6_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08957__A1 net1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07126_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[512\] net785
+ net752 _03067_ vssd1 vssd1 vccd1 vccd1 _03068_ sky130_fd_sc_hd__a211o_1
XFILLER_0_15_487 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_3086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10764__A1 net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10084__B _05142_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11961__B1 net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07057_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[930\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[898\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[802\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[770\]
+ net776 net1132 vssd1 vssd1 vccd1 vccd1 _02999_ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout1312_A net1330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput140 net140 vssd1 vssd1 vccd1 vccd1 DAT_O[13] sky130_fd_sc_hd__buf_2
Xoutput151 net151 vssd1 vssd1 vccd1 vccd1 DAT_O[23] sky130_fd_sc_hd__clkbuf_4
Xoutput162 net162 vssd1 vssd1 vccd1 vccd1 DAT_O[4] sky130_fd_sc_hd__buf_2
Xoutput173 net173 vssd1 vssd1 vccd1 vccd1 WE_O sky130_fd_sc_hd__clkbuf_4
XFILLER_0_100_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput184 net184 vssd1 vssd1 vccd1 vccd1 gpio_oeb[19] sky130_fd_sc_hd__buf_2
XANTENNA__11908__B net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput195 net195 vssd1 vssd1 vccd1 vccd1 gpio_oeb[30] sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout393_X net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout772_A net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11196__A net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout560_X net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07959_ net1147 net1019 net684 vssd1 vssd1 vccd1 vccd1 _03901_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout658_X net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10819__A2 net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10970_ _06547_ _06548_ _06549_ vssd1 vssd1 vccd1 vccd1 _06550_ sky130_fd_sc_hd__a21oi_4
XANTENNA__08342__C1 net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_2590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09629_ _03314_ _04415_ vssd1 vssd1 vccd1 vccd1 _05571_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_67_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10091__A_N _05583_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout825_X net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_502 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_139_3229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12640_ net1396 vssd1 vssd1 vccd1 vccd1 _00404_ sky130_fd_sc_hd__inv_2
XFILLER_0_167_356 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07448__A1 net1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08645__B1 net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12571_ net1361 vssd1 vssd1 vccd1 vccd1 _00335_ sky130_fd_sc_hd__inv_2
XANTENNA__11244__A2 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_156_3576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14310_ clknet_leaf_73_wb_clk_i _02074_ _00675_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[664\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_156_3587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07849__A net1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11522_ _06405_ net622 net703 net695 vssd1 vssd1 vccd1 vccd1 _06780_ sky130_fd_sc_hd__and4_1
XFILLER_0_110_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_776 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14241_ clknet_leaf_180_wb_clk_i _02005_ _00606_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[595\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11453_ net2305 net392 _06765_ net501 vssd1 vssd1 vccd1 vccd1 _02040_ sky130_fd_sc_hd__a22o_1
XANTENNA__08948__A1 net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10404_ _06070_ _06079_ vssd1 vssd1 vccd1 vccd1 _06229_ sky130_fd_sc_hd__xnor2_1
X_14172_ clknet_leaf_154_wb_clk_i _01936_ _00537_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[526\]
+ sky130_fd_sc_hd__dfrtp_1
X_11384_ net508 net636 _06744_ net402 net2136 vssd1 vssd1 vccd1 vccd1 _02088_ sky130_fd_sc_hd__a32o_1
XANTENNA__10755__A1 _05757_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06959__B1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11952__B1 net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13123_ net1373 vssd1 vssd1 vccd1 vccd1 _00887_ sky130_fd_sc_hd__inv_2
X_10335_ net283 _06151_ _06169_ net679 vssd1 vssd1 vccd1 vccd1 _06173_ sky130_fd_sc_hd__o31a_1
XANTENNA__07620__A1 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13054_ net1410 vssd1 vssd1 vccd1 vccd1 _00818_ sky130_fd_sc_hd__inv_2
X_10266_ _03528_ _05978_ vssd1 vssd1 vccd1 vccd1 _06108_ sky130_fd_sc_hd__and2_1
XFILLER_0_44_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11704__B1 net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12005_ net267 net2485 net445 vssd1 vssd1 vccd1 vccd1 _01539_ sky130_fd_sc_hd__mux2_1
Xfanout1310 net1312 vssd1 vssd1 vccd1 vccd1 net1310 sky130_fd_sc_hd__buf_4
Xfanout1321 net1324 vssd1 vssd1 vccd1 vccd1 net1321 sky130_fd_sc_hd__buf_4
Xfanout1332 net1339 vssd1 vssd1 vccd1 vccd1 net1332 sky130_fd_sc_hd__buf_4
Xfanout1343 net1344 vssd1 vssd1 vccd1 vccd1 net1343 sky130_fd_sc_hd__buf_4
X_10197_ team_03_WB.instance_to_wrap.core.pc.current_pc\[4\] net660 _06038_ vssd1
+ vssd1 vccd1 vccd1 _06039_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07384__B1 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1354 net1358 vssd1 vssd1 vccd1 vccd1 net1354 sky130_fd_sc_hd__buf_4
XANTENNA__11180__B2 net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1365 net1367 vssd1 vssd1 vccd1 vccd1 net1365 sky130_fd_sc_hd__buf_4
XFILLER_0_79_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1376 net1381 vssd1 vssd1 vccd1 vccd1 net1376 sky130_fd_sc_hd__buf_4
Xfanout1387 net1393 vssd1 vssd1 vccd1 vccd1 net1387 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09125__A1 net1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1398 net1408 vssd1 vssd1 vccd1 vccd1 net1398 sky130_fd_sc_hd__buf_2
XFILLER_0_89_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_128_2999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07136__B1 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13956_ clknet_leaf_36_wb_clk_i _01720_ _00321_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[310\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09676__A2 _04119_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06928__A net1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14918__Q team_03_WB.instance_to_wrap.CPU_DAT_O\[5\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_12907_ net1281 vssd1 vssd1 vccd1 vccd1 _00671_ sky130_fd_sc_hd__inv_2
XANTENNA__11483__A2 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13887_ clknet_leaf_20_wb_clk_i _01651_ _00252_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[241\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_124_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07151__A3 net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_908 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12838_ net1293 vssd1 vssd1 vccd1 vccd1 _00602_ sky130_fd_sc_hd__inv_2
XFILLER_0_115_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10169__B net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_507 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_68 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12769_ net1271 vssd1 vssd1 vccd1 vccd1 _00533_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_168_wb_clk_i clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_168_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_71_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14508_ clknet_leaf_16_wb_clk_i _02272_ _00873_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[862\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_142_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput20 DAT_I[26] vssd1 vssd1 vccd1 vccd1 net20 sky130_fd_sc_hd__buf_1
XFILLER_0_86_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10185__A _03430_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14439_ clknet_leaf_110_wb_clk_i _02203_ _00804_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[793\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput31 DAT_I[7] vssd1 vssd1 vccd1 vccd1 net31 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_142_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput42 gpio_in[17] vssd1 vssd1 vccd1 vccd1 net42 sky130_fd_sc_hd__clkbuf_1
Xinput53 gpio_in[28] vssd1 vssd1 vccd1 vccd1 net53 sky130_fd_sc_hd__clkbuf_1
Xinput64 gpio_in[8] vssd1 vssd1 vccd1 vccd1 net64 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_130_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold804 team_03_WB.instance_to_wrap.core.register_file.registers_state\[755\] vssd1
+ vssd1 vccd1 vccd1 net2297 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput75 wbs_adr_i[17] vssd1 vssd1 vccd1 vccd1 net75 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_80_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10746__A1 net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput86 wbs_adr_i[27] vssd1 vssd1 vccd1 vccd1 net86 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_141_267 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold815 team_03_WB.instance_to_wrap.core.register_file.registers_state\[919\] vssd1
+ vssd1 vccd1 vccd1 net2308 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_295 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_744 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold826 team_03_WB.instance_to_wrap.core.register_file.registers_state\[367\] vssd1
+ vssd1 vccd1 vccd1 net2319 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput97 wbs_adr_i[8] vssd1 vssd1 vccd1 vccd1 net97 sky130_fd_sc_hd__clkbuf_1
XANTENNA__11943__B1 net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold837 team_03_WB.instance_to_wrap.core.register_file.registers_state\[663\] vssd1
+ vssd1 vccd1 vccd1 net2330 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13496__A net1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07611__A1 net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold848 team_03_WB.instance_to_wrap.core.register_file.registers_state\[631\] vssd1
+ vssd1 vccd1 vccd1 net2341 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_2222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09980_ _03103_ net1663 net294 vssd1 vssd1 vccd1 vccd1 _02733_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_90_2233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold859 team_03_WB.instance_to_wrap.core.register_file.registers_state\[640\] vssd1
+ vssd1 vccd1 vccd1 net2352 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09039__S1 net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08931_ net1051 team_03_WB.instance_to_wrap.core.register_file.registers_state\[459\]
+ net1001 team_03_WB.instance_to_wrap.core.register_file.registers_state\[491\] net1075
+ vssd1 vssd1 vccd1 vccd1 _04873_ sky130_fd_sc_hd__a221o_1
XFILLER_0_58_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09364__A1 _05278_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08862_ net1223 _04802_ _04803_ vssd1 vssd1 vccd1 vccd1 _04804_ sky130_fd_sc_hd__and3_1
XANTENNA__07781__X _03723_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08572__C1 net1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07813_ net824 _03754_ net723 vssd1 vssd1 vccd1 vccd1 _03755_ sky130_fd_sc_hd__a21oi_1
X_08793_ net1050 team_03_WB.instance_to_wrap.core.register_file.registers_state\[578\]
+ net1002 team_03_WB.instance_to_wrap.core.register_file.registers_state\[610\] net940
+ vssd1 vssd1 vccd1 vccd1 _04735_ sky130_fd_sc_hd__a221o_1
XANTENNA__09116__A1 net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07744_ net1194 team_03_WB.instance_to_wrap.core.register_file.registers_state\[172\]
+ net898 net1133 vssd1 vssd1 vccd1 vccd1 _03686_ sky130_fd_sc_hd__a211oi_1
XTAP_TAPCELL_ROW_88_2184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09214__A _02937_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08875__B1 net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11474__A2 net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07675_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[446\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[414\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[318\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[286\]
+ net767 net1127 vssd1 vssd1 vccd1 vccd1 _03617_ sky130_fd_sc_hd__mux4_1
X_09414_ net320 vssd1 vssd1 vccd1 vccd1 _05356_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout1095_A net1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_490 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09345_ _03137_ _05286_ vssd1 vssd1 vccd1 vccd1 _05287_ sky130_fd_sc_hd__xor2_1
XANTENNA__08627__B1 net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout520_A _06395_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06844__Y _02787_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout618_A net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_941 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1262_A net1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08772__B net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_151 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_33_Left_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10434__B1 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07669__A net1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_134_3126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09276_ _03244_ _03790_ _05145_ net609 vssd1 vssd1 vccd1 vccd1 _05218_ sky130_fd_sc_hd__a31o_1
XFILLER_0_118_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_134_3137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_798 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08227_ net1061 _04167_ _04168_ net1211 vssd1 vssd1 vccd1 vccd1 _04169_ sky130_fd_sc_hd__a211o_1
XANTENNA__07388__B net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1050_X net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout406_X net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1148_X net1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_151_3473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_23_wb_clk_i_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_160_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_151_3484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08158_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[436\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[404\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[308\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[276\]
+ net961 net1071 vssd1 vssd1 vccd1 vccd1 _04100_ sky130_fd_sc_hd__mux4_1
XANTENNA__09052__B1 net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10198__C1 _02889_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11934__A0 net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout987_A net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07109_ net1100 team_03_WB.instance_to_wrap.core.register_file.registers_state\[193\]
+ net799 team_03_WB.instance_to_wrap.core.register_file.registers_state\[225\] net731
+ vssd1 vssd1 vccd1 vccd1 _03051_ sky130_fd_sc_hd__a221oi_1
XANTENNA__07602__A1 net1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08089_ _04029_ _04030_ net610 vssd1 vssd1 vccd1 vccd1 _04031_ sky130_fd_sc_hd__mux2_2
XANTENNA_fanout1315_X net1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09095__S net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10120_ _03640_ _05961_ vssd1 vssd1 vccd1 vccd1 _05962_ sky130_fd_sc_hd__and2b_1
XANTENNA_fanout775_X net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_490 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_42_Left_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08789__S0 net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10051_ net5 net1037 net910 net2768 vssd1 vssd1 vccd1 vccd1 _02680_ sky130_fd_sc_hd__o22a_1
XANTENNA__11357__C net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout942_X net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09107__A1 net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13810_ clknet_leaf_117_wb_clk_i _01574_ _00175_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[164\]
+ sky130_fd_sc_hd__dfrtp_1
X_14790_ clknet_leaf_105_wb_clk_i _02554_ _01155_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_I\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08315__C1 net1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_2549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13741_ clknet_leaf_189_wb_clk_i _01505_ _00106_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[95\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10953_ _06533_ _06534_ _06535_ _06399_ vssd1 vssd1 vccd1 vccd1 _06536_ sky130_fd_sc_hd__o211a_4
XANTENNA__11465__A2 net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07570__C net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_158_3616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_158_3627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11941__X _06815_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_168_654 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1046 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_123_2896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13672_ clknet_leaf_8_wb_clk_i _01436_ _00037_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_79_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10884_ net495 net596 _06479_ net518 net1749 vssd1 vssd1 vccd1 vccd1 _02323_ sky130_fd_sc_hd__a32o_1
XFILLER_0_167_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_687 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_51_Left_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12623_ net1336 vssd1 vssd1 vccd1 vccd1 _00387_ sky130_fd_sc_hd__inv_2
XFILLER_0_38_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_62_wb_clk_i_A clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_94_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08618__B1 net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12554_ net1279 vssd1 vssd1 vccd1 vccd1 _00318_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_14_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09830__A2 _04711_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11505_ _06623_ net2703 net389 vssd1 vssd1 vccd1 vccd1 _02001_ sky130_fd_sc_hd__mux2_1
XANTENNA__06914__C net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07841__A1 net1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_151_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12485_ net1353 vssd1 vssd1 vccd1 vccd1 _00249_ sky130_fd_sc_hd__inv_2
XFILLER_0_124_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input71_X net71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14224_ clknet_leaf_156_wb_clk_i _01988_ _00589_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[578\]
+ sky130_fd_sc_hd__dfrtp_1
X_11436_ _06405_ net618 net703 net827 vssd1 vssd1 vccd1 vccd1 _06758_ sky130_fd_sc_hd__and4_1
XANTENNA__10728__A1 _05632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11925__A0 _06623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_638 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07054__C1 net1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14155_ clknet_leaf_38_wb_clk_i _01919_ _00520_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[509\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_145_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11367_ net713 net271 net698 vssd1 vssd1 vccd1 vccd1 _06736_ sky130_fd_sc_hd__and3_1
XFILLER_0_10_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06930__B net1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13106_ net1396 vssd1 vssd1 vccd1 vccd1 _00870_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_60_Left_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10318_ _06153_ _06158_ vssd1 vssd1 vccd1 vccd1 _06159_ sky130_fd_sc_hd__nand2_1
X_14086_ clknet_leaf_28_wb_clk_i _01850_ _00451_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[440\]
+ sky130_fd_sc_hd__dfrtp_1
X_11298_ net514 net645 _06716_ net410 net2191 vssd1 vssd1 vccd1 vccd1 _02146_ sky130_fd_sc_hd__a32o_1
XANTENNA__10452__B net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13037_ net1292 vssd1 vssd1 vccd1 vccd1 _00801_ sky130_fd_sc_hd__inv_2
X_10249_ _03426_ _06090_ vssd1 vssd1 vccd1 vccd1 _06091_ sky130_fd_sc_hd__nand2_1
XFILLER_0_119_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11153__A1 net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11267__C net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1140 net1141 vssd1 vssd1 vccd1 vccd1 net1140 sky130_fd_sc_hd__buf_2
Xfanout1151 net1159 vssd1 vssd1 vccd1 vccd1 net1151 sky130_fd_sc_hd__clkbuf_4
Xfanout1162 net1169 vssd1 vssd1 vccd1 vccd1 net1162 sky130_fd_sc_hd__buf_4
XANTENNA__10900__A1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1173 net1174 vssd1 vssd1 vccd1 vccd1 net1173 sky130_fd_sc_hd__clkbuf_2
Xfanout1184 net1190 vssd1 vssd1 vccd1 vccd1 net1184 sky130_fd_sc_hd__buf_2
XANTENNA__06929__Y _02871_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1195 net1199 vssd1 vssd1 vccd1 vccd1 net1195 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_135_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07109__B1 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14988_ clknet_leaf_64_wb_clk_i net36 _01353_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12102__B1 net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_232 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11283__B _06523_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13939_ clknet_leaf_108_wb_clk_i _01703_ _00304_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[293\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09969__A _03241_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07755__S1 net1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07460_ net1183 team_03_WB.instance_to_wrap.core.register_file.registers_state\[341\]
+ net770 team_03_WB.instance_to_wrap.core.register_file.registers_state\[373\] net1128
+ vssd1 vssd1 vccd1 vccd1 _03402_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_83_2081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07391_ net821 _03324_ _03327_ _03332_ vssd1 vssd1 vccd1 vccd1 _03333_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_29_354 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11503__S net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09130_ _04895_ _04956_ _05014_ _05071_ net555 net566 vssd1 vssd1 vccd1 vccd1 _05072_
+ sky130_fd_sc_hd__mux4_2
XANTENNA__11759__A3 net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08085__A1 net1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_77 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09282__B1 _02937_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_40_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08624__A3 _04565_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09061_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[559\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[527\]
+ net971 vssd1 vssd1 vccd1 vccd1 _05003_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08012_ net1177 team_03_WB.instance_to_wrap.core.register_file.registers_state\[721\]
+ net764 team_03_WB.instance_to_wrap.core.register_file.registers_state\[753\] net742
+ vssd1 vssd1 vccd1 vccd1 _03954_ sky130_fd_sc_hd__o221a_1
XFILLER_0_72_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold601 team_03_WB.instance_to_wrap.core.register_file.registers_state\[98\] vssd1
+ vssd1 vccd1 vccd1 net2094 sky130_fd_sc_hd__dlygate4sd3_1
Xhold612 team_03_WB.instance_to_wrap.core.register_file.registers_state\[240\] vssd1
+ vssd1 vccd1 vccd1 net2105 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10065__D team_03_WB.instance_to_wrap.core.decoder.inst\[19\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold623 team_03_WB.instance_to_wrap.core.register_file.registers_state\[829\] vssd1
+ vssd1 vccd1 vccd1 net2116 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07045__C1 net1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold634 team_03_WB.instance_to_wrap.core.register_file.registers_state\[328\] vssd1
+ vssd1 vccd1 vccd1 net2127 sky130_fd_sc_hd__dlygate4sd3_1
Xhold645 team_03_WB.instance_to_wrap.core.register_file.registers_state\[693\] vssd1
+ vssd1 vccd1 vccd1 net2138 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07596__B1 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold656 team_03_WB.instance_to_wrap.core.register_file.registers_state\[44\] vssd1
+ vssd1 vccd1 vccd1 net2149 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11392__A1 net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold667 team_03_WB.instance_to_wrap.core.register_file.registers_state\[746\] vssd1
+ vssd1 vccd1 vccd1 net2160 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08793__C1 net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_107_wb_clk_i_A clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_4_Right_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold678 team_03_WB.instance_to_wrap.core.register_file.registers_state\[356\] vssd1
+ vssd1 vccd1 vccd1 net2171 sky130_fd_sc_hd__dlygate4sd3_1
X_09963_ _03723_ net661 vssd1 vssd1 vccd1 vccd1 _05886_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_38_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold689 team_03_WB.instance_to_wrap.core.register_file.registers_state\[505\] vssd1
+ vssd1 vccd1 vccd1 net2182 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_65_wb_clk_i clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_65_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_08914_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[940\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[908\]
+ net979 vssd1 vssd1 vccd1 vccd1 _04856_ sky130_fd_sc_hd__mux2_1
X_09894_ _04031_ _04323_ net664 _05835_ vssd1 vssd1 vccd1 vccd1 _05836_ sky130_fd_sc_hd__a22o_1
XANTENNA__10930__X _06517_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1010_A net1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09888__A2 _03109_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1108_A net1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1040 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08845_ _04783_ _04786_ net868 vssd1 vssd1 vccd1 vccd1 _04787_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07899__A1 net1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07443__S0 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11695__A2 net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout470_A net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout568_A net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08776_ net1055 team_03_WB.instance_to_wrap.core.register_file.registers_state\[66\]
+ net1002 team_03_WB.instance_to_wrap.core.register_file.registers_state\[98\] net940
+ vssd1 vssd1 vccd1 vccd1 _04718_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_108_Left_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07727_ _03663_ _03668_ net1140 vssd1 vssd1 vccd1 vccd1 _03669_ sky130_fd_sc_hd__o21a_1
XANTENNA__11447__A2 net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout735_A net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout356_X net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1098_X net1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07658_ _03585_ _03586_ _03599_ net723 vssd1 vssd1 vccd1 vccd1 _03600_ sky130_fd_sc_hd__a22o_4
XTAP_TAPCELL_ROW_0_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_0_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08783__A net1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07520__B1 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_101_2446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout523_X net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout902_A net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07589_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[25\] net787
+ net752 _03530_ vssd1 vssd1 vccd1 vccd1 _03531_ sky130_fd_sc_hd__a211o_1
XANTENNA__10818__A net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10407__B1 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_153_3513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09328_ _05246_ _05250_ _05269_ _05244_ vssd1 vssd1 vccd1 vccd1 _05270_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_153_3524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_819 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09259_ net589 _05200_ vssd1 vssd1 vccd1 vccd1 _05201_ sky130_fd_sc_hd__or2_1
XANTENNA_clkbuf_leaf_146_wb_clk_i_A clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__07823__A1 net1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_170_3860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_170_3871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_117_Left_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12270_ net1274 vssd1 vssd1 vccd1 vccd1 _00034_ sky130_fd_sc_hd__inv_2
XANTENNA__08722__S net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_530 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout892_X net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11907__B1 net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09576__A1 net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11221_ net2178 net486 _06682_ net495 vssd1 vssd1 vccd1 vccd1 _02189_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_79_1994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07587__A0 _03526_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07051__A2 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11152_ net703 net273 net695 vssd1 vssd1 vccd1 vccd1 _06653_ sky130_fd_sc_hd__and3_1
X_10103_ net683 net286 vssd1 vssd1 vccd1 vccd1 _05947_ sky130_fd_sc_hd__nand2_1
XFILLER_0_105_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11083_ _06619_ net2101 net417 vssd1 vssd1 vccd1 vccd1 _02264_ sky130_fd_sc_hd__mux2_1
XANTENNA__11135__A1 net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input31_A DAT_I[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14911_ clknet_leaf_55_wb_clk_i _00005_ _01276_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.ru.state\[5\]
+ sky130_fd_sc_hd__dfrtp_4
X_10034_ net23 net1038 net910 net1808 vssd1 vssd1 vccd1 vccd1 _02697_ sky130_fd_sc_hd__o22a_1
XANTENNA__11686__A2 net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10894__A0 net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14842_ clknet_leaf_87_wb_clk_i _02606_ _01207_ vssd1 vssd1 vccd1 vccd1 net128 sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_125_2936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08169__S net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08839__B1 net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14773_ clknet_leaf_104_wb_clk_i _02537_ _01138_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_I\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_11985_ _06446_ net2606 net446 vssd1 vssd1 vccd1 vccd1 _01559_ sky130_fd_sc_hd__mux2_1
XANTENNA__11534__D net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10646__A0 net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10936_ team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[7\] net312 _05845_ net318
+ vssd1 vssd1 vccd1 vccd1 _06522_ sky130_fd_sc_hd__and4_1
XFILLER_0_129_805 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13724_ clknet_leaf_148_wb_clk_i _01488_ _00089_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[78\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_185_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_169_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13655_ clknet_leaf_96_wb_clk_i _01419_ _00020_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[9\]
+ sky130_fd_sc_hd__dfrtp_2
X_10867_ team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[19\] net306 vssd1
+ vssd1 vccd1 vccd1 _06465_ sky130_fd_sc_hd__and2_1
XANTENNA__11323__S net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_156_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12606_ net1414 vssd1 vssd1 vccd1 vccd1 _00370_ sky130_fd_sc_hd__inv_2
X_13586_ net1345 vssd1 vssd1 vccd1 vccd1 _01350_ sky130_fd_sc_hd__inv_2
XANTENNA__08980__X _04922_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10798_ net311 net310 net317 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[30\]
+ vssd1 vssd1 vccd1 vccd1 _06407_ sky130_fd_sc_hd__a31o_1
XFILLER_0_112_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12537_ net1365 vssd1 vssd1 vccd1 vccd1 _00301_ sky130_fd_sc_hd__inv_2
XFILLER_0_152_852 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12468_ net1304 vssd1 vssd1 vccd1 vccd1 _00232_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11419_ _06499_ net2302 net398 vssd1 vssd1 vccd1 vccd1 _02062_ sky130_fd_sc_hd__mux2_1
XANTENNA__11559__A net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14207_ clknet_leaf_21_wb_clk_i _01971_ _00572_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[561\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_111_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12007__X _06817_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12399_ net1394 vssd1 vssd1 vccd1 vccd1 _00163_ sky130_fd_sc_hd__inv_2
XANTENNA__11374__A1 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14138_ clknet_leaf_144_wb_clk_i _01902_ _00503_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[492\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10182__B net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11993__S net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09971__B net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14069_ clknet_leaf_107_wb_clk_i _01833_ _00434_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[423\]
+ sky130_fd_sc_hd__dfrtp_1
X_06960_ net1112 team_03_WB.instance_to_wrap.core.register_file.registers_state\[453\]
+ net802 team_03_WB.instance_to_wrap.core.register_file.registers_state\[485\] net1135
+ vssd1 vssd1 vccd1 vccd1 _02902_ sky130_fd_sc_hd__a221o_1
XANTENNA__08527__C1 net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06891_ _02799_ _02832_ vssd1 vssd1 vccd1 vccd1 _02833_ sky130_fd_sc_hd__nand2_1
XANTENNA__11677__A2 net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08630_ net1054 team_03_WB.instance_to_wrap.core.register_file.registers_state\[198\]
+ net1007 team_03_WB.instance_to_wrap.core.register_file.registers_state\[230\] net927
+ vssd1 vssd1 vccd1 vccd1 _04572_ sky130_fd_sc_hd__a221o_1
XFILLER_0_55_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_85_2121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07750__B1 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08561_ net851 _04502_ _04491_ vssd1 vssd1 vccd1 vccd1 _04503_ sky130_fd_sc_hd__o21a_4
XANTENNA__10637__A0 team_03_WB.instance_to_wrap.core.decoder.inst\[24\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_183_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_183_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_07512_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[423\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[391\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[295\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[263\]
+ net786 net1135 vssd1 vssd1 vccd1 vccd1 _03454_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_18_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08492_ net1242 team_03_WB.instance_to_wrap.core.register_file.registers_state\[91\]
+ net985 team_03_WB.instance_to_wrap.core.register_file.registers_state\[123\] net929
+ vssd1 vssd1 vccd1 vccd1 _04434_ sky130_fd_sc_hd__o221a_1
XFILLER_0_49_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_112_wb_clk_i clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_112_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_71_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07443_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[436\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[404\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[308\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[276\]
+ net764 net1125 vssd1 vssd1 vccd1 vccd1 _03385_ sky130_fd_sc_hd__mux4_1
XFILLER_0_92_706 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11233__S net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07374_ net1175 team_03_WB.instance_to_wrap.core.register_file.registers_state\[63\]
+ net880 vssd1 vssd1 vccd1 vccd1 _03316_ sky130_fd_sc_hd__and3_1
XFILLER_0_73_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_146_178 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07012__A net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09113_ _05049_ _05054_ net873 vssd1 vssd1 vccd1 vccd1 _05055_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10925__X _06513_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1058_A net1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09044_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[47\] net971
+ vssd1 vssd1 vccd1 vccd1 _04986_ sky130_fd_sc_hd__or2_1
XANTENNA__09007__B1 net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14841__Q net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold420 team_03_WB.instance_to_wrap.core.register_file.registers_state\[297\] vssd1
+ vssd1 vccd1 vccd1 net1913 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12064__S net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold431 team_03_WB.instance_to_wrap.core.register_file.registers_state\[384\] vssd1
+ vssd1 vccd1 vccd1 net1924 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold442 team_03_WB.instance_to_wrap.core.register_file.registers_state\[187\] vssd1
+ vssd1 vccd1 vccd1 net1935 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08766__C1 net1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold453 team_03_WB.instance_to_wrap.core.register_file.registers_state\[436\] vssd1
+ vssd1 vccd1 vccd1 net1946 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11904__A3 net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07033__A2 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08230__A1 net1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold464 team_03_WB.instance_to_wrap.core.register_file.registers_state\[689\] vssd1
+ vssd1 vccd1 vccd1 net1957 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11188__B net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold475 team_03_WB.instance_to_wrap.core.register_file.registers_state\[509\] vssd1
+ vssd1 vccd1 vccd1 net1968 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_3025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold486 team_03_WB.instance_to_wrap.core.register_file.registers_state\[900\] vssd1
+ vssd1 vccd1 vccd1 net1979 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout685_A net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout900 net904 vssd1 vssd1 vccd1 vccd1 net900 sky130_fd_sc_hd__clkbuf_4
Xfanout911 _05906_ vssd1 vssd1 vccd1 vccd1 net911 sky130_fd_sc_hd__buf_2
XFILLER_0_1_991 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold497 team_03_WB.instance_to_wrap.core.register_file.registers_state\[429\] vssd1
+ vssd1 vccd1 vccd1 net1990 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout922 net923 vssd1 vssd1 vccd1 vccd1 net922 sky130_fd_sc_hd__clkbuf_4
X_09946_ _05877_ net1734 net292 vssd1 vssd1 vccd1 vccd1 _02754_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_74_1891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1013_X net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout933 net934 vssd1 vssd1 vccd1 vccd1 net933 sky130_fd_sc_hd__buf_4
Xfanout944 net948 vssd1 vssd1 vccd1 vccd1 net944 sky130_fd_sc_hd__clkbuf_4
Xfanout955 net956 vssd1 vssd1 vccd1 vccd1 net955 sky130_fd_sc_hd__buf_4
XANTENNA__07682__A net1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout966 net969 vssd1 vssd1 vccd1 vccd1 net966 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_146_3372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout977 net978 vssd1 vssd1 vccd1 vccd1 net977 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_146_3383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09877_ _03604_ _05069_ _05818_ vssd1 vssd1 vccd1 vccd1 _05819_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout852_A _04096_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout473_X net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1120 team_03_WB.instance_to_wrap.core.register_file.registers_state\[151\] vssd1
+ vssd1 vccd1 vccd1 net2613 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout988 net994 vssd1 vssd1 vccd1 vccd1 net988 sky130_fd_sc_hd__clkbuf_4
Xfanout999 net1000 vssd1 vssd1 vccd1 vccd1 net999 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_5_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11408__S net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1131 team_03_WB.instance_to_wrap.core.register_file.registers_state\[662\] vssd1
+ vssd1 vccd1 vccd1 net2624 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1142 team_03_WB.instance_to_wrap.core.register_file.registers_state\[214\] vssd1
+ vssd1 vccd1 vccd1 net2635 sky130_fd_sc_hd__dlygate4sd3_1
X_08828_ _04769_ _04768_ _04754_ _04748_ vssd1 vssd1 vccd1 vccd1 _04770_ sky130_fd_sc_hd__a2bb2o_4
Xhold1153 team_03_WB.instance_to_wrap.core.register_file.registers_state\[477\] vssd1
+ vssd1 vccd1 vccd1 net2646 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1164 team_03_WB.instance_to_wrap.core.register_file.registers_state\[144\] vssd1
+ vssd1 vccd1 vccd1 net2657 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1175 net175 vssd1 vssd1 vccd1 vccd1 net2668 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_79_Right_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1186 team_03_WB.instance_to_wrap.core.register_file.registers_state\[837\] vssd1
+ vssd1 vccd1 vccd1 net2679 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout640_X net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08759_ net1065 _04697_ _04700_ vssd1 vssd1 vccd1 vccd1 _04701_ sky130_fd_sc_hd__a21oi_1
Xhold1197 team_03_WB.instance_to_wrap.core.register_file.registers_state\[708\] vssd1
+ vssd1 vccd1 vccd1 net2690 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_135_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10891__A3 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout738_X net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11770_ net658 _06603_ net479 net334 net2225 vssd1 vssd1 vccd1 vccd1 _01767_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_120_2833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12093__A2 net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_2844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10721_ team_03_WB.instance_to_wrap.core.pc.current_pc\[20\] _05623_ net602 vssd1
+ vssd1 vccd1 vccd1 _06352_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_172_3900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout905_X net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11840__A2 net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_172_3911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13440_ net1405 vssd1 vssd1 vccd1 vccd1 _01204_ sky130_fd_sc_hd__inv_2
X_10652_ net1250 team_03_WB.instance_to_wrap.CPU_DAT_O\[9\] net845 vssd1 vssd1 vccd1
+ vccd1 _02476_ sky130_fd_sc_hd__mux2_1
XANTENNA__09246__B1 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_125_Left_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13371_ net1321 vssd1 vssd1 vccd1 vccd1 _01135_ sky130_fd_sc_hd__inv_2
X_10583_ net1644 net531 net598 _02921_ vssd1 vssd1 vccd1 vccd1 _02540_ sky130_fd_sc_hd__a22o_1
XFILLER_0_24_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15110_ net912 vssd1 vssd1 vccd1 vccd1 net244 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_35_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12322_ net1360 vssd1 vssd1 vccd1 vccd1 _00086_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_88_Right_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10800__B1 net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input79_A wbs_adr_i[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_2795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15041_ clknet_leaf_84_wb_clk_i _02761_ _01406_ vssd1 vssd1 vccd1 vccd1 net197 sky130_fd_sc_hd__dfrtp_1
XANTENNA__11379__A net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12253_ net1389 vssd1 vssd1 vccd1 vccd1 _00017_ sky130_fd_sc_hd__inv_2
XFILLER_0_160_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11356__A1 net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09013__A3 _04953_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08757__C1 net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11204_ _06426_ net2425 net487 vssd1 vssd1 vccd1 vccd1 _02204_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_1134 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12184_ net1514 vssd1 vssd1 vccd1 vccd1 _02369_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__07655__S0 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11135_ net497 net649 _06643_ net413 net1959 vssd1 vssd1 vccd1 vccd1 _02236_ sky130_fd_sc_hd__a32o_1
XANTENNA__08509__C1 net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11066_ net833 net280 vssd1 vssd1 vccd1 vccd1 _06611_ sky130_fd_sc_hd__and2_2
XANTENNA__11164__C_N net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11318__S net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_97_Right_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10017_ net71 net70 net73 net72 vssd1 vssd1 vccd1 vccd1 _05895_ sky130_fd_sc_hd__or4_1
XFILLER_0_92_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14825_ clknet_leaf_90_wb_clk_i net1780 _01190_ vssd1 vssd1 vccd1 vccd1 net145 sky130_fd_sc_hd__dfrtp_1
XANTENNA__12938__A net1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14756_ clknet_leaf_50_wb_clk_i net1620 _01121_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_11968_ net643 _06745_ net479 net366 net1937 vssd1 vssd1 vccd1 vccd1 _01575_ sky130_fd_sc_hd__a32o_1
XANTENNA__09312__A net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13707_ clknet_leaf_46_wb_clk_i _01471_ _00072_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[61\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11292__B1 net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07496__C1 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10919_ team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[10\] net307 net685 vssd1
+ vssd1 vccd1 vccd1 _06508_ sky130_fd_sc_hd__a21oi_2
X_14687_ clknet_leaf_64_wb_clk_i _02451_ _01052_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.ADR_I\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_11899_ net623 _06708_ net454 net371 net2346 vssd1 vssd1 vccd1 vccd1 _01642_ sky130_fd_sc_hd__a32o_1
XFILLER_0_46_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_157_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13638_ net1428 vssd1 vssd1 vccd1 vccd1 _01402_ sky130_fd_sc_hd__inv_2
XFILLER_0_116_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10177__B net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_156_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09788__A1 net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11988__S net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_901 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13569_ net1429 vssd1 vssd1 vccd1 vccd1 _01333_ sky130_fd_sc_hd__inv_2
XFILLER_0_125_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07799__B1 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08996__C1 net1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07090_ net1198 team_03_WB.instance_to_wrap.core.register_file.registers_state\[609\]
+ net884 _03031_ vssd1 vssd1 vccd1 vccd1 _03032_ sky130_fd_sc_hd__a31o_1
XFILLER_0_81_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_140_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_822 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11289__A net1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_160_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_wire274_X net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09800_ net540 _05741_ vssd1 vssd1 vccd1 vccd1 _05742_ sky130_fd_sc_hd__nand2_1
X_07992_ net1140 _03933_ net723 vssd1 vssd1 vccd1 vccd1 _03934_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10570__A2 net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07971__B1 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_1011 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_163_Right_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09731_ net584 _05672_ vssd1 vssd1 vccd1 vccd1 _05673_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_52_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06943_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[868\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[836\]
+ net776 vssd1 vssd1 vccd1 vccd1 _02885_ sky130_fd_sc_hd__mux2_1
XANTENNA__11228__S net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10132__S net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09662_ _03170_ _04207_ vssd1 vssd1 vccd1 vccd1 _05604_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_2_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06874_ team_03_WB.instance_to_wrap.core.control_logic.instruction\[6\] team_03_WB.instance_to_wrap.core.control_logic.instruction\[5\]
+ _02794_ vssd1 vssd1 vccd1 vccd1 _02816_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_2_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07723__B1 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08613_ _04553_ _04554_ net858 vssd1 vssd1 vccd1 vccd1 _04555_ sky130_fd_sc_hd__o21a_1
XANTENNA__07007__A net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09593_ net563 _05415_ vssd1 vssd1 vccd1 vccd1 _05535_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_141_3280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout266_A _06557_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08544_ net1063 _04484_ _04485_ vssd1 vssd1 vccd1 vccd1 _04486_ sky130_fd_sc_hd__or3_1
XANTENNA__06846__A net1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12075__A2 net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09222__A _04503_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08475_ net431 net424 _04415_ vssd1 vssd1 vccd1 vccd1 _04417_ sky130_fd_sc_hd__or3_2
XFILLER_0_49_268 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout433_A net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12059__S net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1175_A net1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07426_ net1086 team_03_WB.instance_to_wrap.core.register_file.registers_state\[948\]
+ net889 vssd1 vssd1 vccd1 vccd1 _03368_ sky130_fd_sc_hd__or3_1
XFILLER_0_174_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11190__C net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07239__C1 net1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07357_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[572\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[540\]
+ net759 vssd1 vssd1 vccd1 vccd1 _03299_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout600_A _06299_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12583__A net1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1342_A net1346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_2389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08987__C1 net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07677__A net1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07288_ net1202 team_03_WB.instance_to_wrap.core.register_file.registers_state\[73\]
+ net788 team_03_WB.instance_to_wrap.core.register_file.registers_state\[105\] net734
+ vssd1 vssd1 vccd1 vccd1 _03230_ sky130_fd_sc_hd__o221a_1
Xclkbuf_leaf_80_wb_clk_i clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_80_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_115_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09027_ net1223 _04967_ _04968_ vssd1 vssd1 vccd1 vccd1 _04969_ sky130_fd_sc_hd__o21a_1
XFILLER_0_62_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_1931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1130_X net1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11338__A1 net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_1942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1228_X net1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold250 team_03_WB.instance_to_wrap.ADR_I\[16\] vssd1 vssd1 vccd1 vccd1 net1743 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_148_3412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_148_3423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold261 team_03_WB.instance_to_wrap.CPU_DAT_I\[11\] vssd1 vssd1 vccd1 vccd1 net1754
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold272 team_03_WB.instance_to_wrap.ADR_I\[24\] vssd1 vssd1 vccd1 vccd1 net1765 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_113_2692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11349__D net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold283 net199 vssd1 vssd1 vccd1 vccd1 net1776 sky130_fd_sc_hd__dlygate4sd3_1
Xhold294 team_03_WB.instance_to_wrap.core.register_file.registers_state\[680\] vssd1
+ vssd1 vccd1 vccd1 net1787 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08754__A2 net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10561__A2 net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout730 net733 vssd1 vssd1 vccd1 vccd1 net730 sky130_fd_sc_hd__clkbuf_4
Xfanout741 net742 vssd1 vssd1 vccd1 vccd1 net741 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_165_3770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09929_ _03277_ net662 vssd1 vssd1 vccd1 vccd1 _05869_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_130_Right_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout752 net754 vssd1 vssd1 vccd1 vccd1 net752 sky130_fd_sc_hd__buf_4
XANTENNA__10550__B net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout763 net765 vssd1 vssd1 vccd1 vccd1 net763 sky130_fd_sc_hd__clkbuf_4
Xfanout774 net777 vssd1 vssd1 vccd1 vccd1 net774 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout855_X net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09703__A1 net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout785 net786 vssd1 vssd1 vccd1 vccd1 net785 sky130_fd_sc_hd__clkbuf_4
Xfanout796 net798 vssd1 vssd1 vccd1 vccd1 net796 sky130_fd_sc_hd__buf_4
X_12940_ net1333 vssd1 vssd1 vccd1 vccd1 _00704_ sky130_fd_sc_hd__inv_2
XANTENNA__08062__S0 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11365__C net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_161_3678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07714__B1 _02869_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_161_3689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08911__C1 net1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12871_ net1400 vssd1 vssd1 vccd1 vccd1 _00635_ sky130_fd_sc_hd__inv_2
X_14610_ clknet_leaf_121_wb_clk_i _02374_ _00975_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[964\]
+ sky130_fd_sc_hd__dfstp_1
X_11822_ net648 _06652_ net454 net323 net1825 vssd1 vssd1 vccd1 vccd1 _01717_ sky130_fd_sc_hd__a32o_1
XFILLER_0_29_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10077__A1 _04475_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_566 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11274__B1 net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14541_ clknet_leaf_188_wb_clk_i _02305_ _00906_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[895\]
+ sky130_fd_sc_hd__dfrtp_1
X_11753_ _06578_ net461 net332 net2360 vssd1 vssd1 vccd1 vccd1 _01784_ sky130_fd_sc_hd__a22o_1
X_10704_ _05933_ _06310_ vssd1 vssd1 vccd1 vccd1 _06341_ sky130_fd_sc_hd__nor2_1
XANTENNA__10709__C net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14472_ clknet_leaf_12_wb_clk_i _02236_ _00837_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[826\]
+ sky130_fd_sc_hd__dfrtp_1
X_11684_ _06726_ net382 net338 net1970 vssd1 vssd1 vccd1 vccd1 _01850_ sky130_fd_sc_hd__a22o_1
XFILLER_0_126_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10635_ team_03_WB.instance_to_wrap.core.decoder.inst\[26\] net2783 net844 vssd1
+ vssd1 vccd1 vccd1 _02493_ sky130_fd_sc_hd__mux2_1
X_13423_ net1420 vssd1 vssd1 vccd1 vccd1 _01187_ sky130_fd_sc_hd__inv_2
XFILLER_0_102_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09427__C_N _05126_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_153_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_260 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_411 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11601__S net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload109 clknet_leaf_157_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload109/Y sky130_fd_sc_hd__clkinv_1
X_13354_ net1308 vssd1 vssd1 vccd1 vccd1 _01118_ sky130_fd_sc_hd__inv_2
XFILLER_0_23_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10566_ net1735 net532 net599 _05876_ vssd1 vssd1 vccd1 vccd1 _02557_ sky130_fd_sc_hd__a22o_1
XFILLER_0_122_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_682 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12305_ net1267 vssd1 vssd1 vccd1 vccd1 _00069_ sky130_fd_sc_hd__inv_2
X_13285_ net1345 vssd1 vssd1 vccd1 vccd1 _01049_ sky130_fd_sc_hd__inv_2
X_10497_ net1739 net1030 net907 net1611 vssd1 vssd1 vccd1 vccd1 _02612_ sky130_fd_sc_hd__a22o_1
XFILLER_0_121_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15024_ clknet_leaf_95_wb_clk_i _02744_ _01389_ vssd1 vssd1 vccd1 vccd1 net180 sky130_fd_sc_hd__dfrtp_1
X_12236_ net1796 vssd1 vssd1 vccd1 vccd1 _01421_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__08910__S net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12167_ net1507 vssd1 vssd1 vccd1 vccd1 _02386_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_120_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10552__A2 _06293_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11118_ net834 net266 vssd1 vssd1 vccd1 vccd1 _06633_ sky130_fd_sc_hd__and2_1
XANTENNA__09307__A _04565_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12098_ _06795_ net477 net442 net2499 vssd1 vssd1 vccd1 vccd1 _01449_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_30_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11049_ net659 net705 _06527_ net829 vssd1 vssd1 vccd1 vccd1 _06602_ sky130_fd_sc_hd__and4_1
XANTENNA__11275__C net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07705__B1 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput7 DAT_I[14] vssd1 vssd1 vccd1 vccd1 net7 sky130_fd_sc_hd__buf_1
XANTENNA__07181__A1 net1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11572__A net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14808_ clknet_leaf_103_wb_clk_i net1615 _01173_ vssd1 vssd1 vccd1 vccd1 net147 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_864 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11291__B net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14739_ clknet_leaf_48_wb_clk_i _02503_ _01104_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10188__A _03460_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_156_240 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08260_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[946\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[914\]
+ net951 vssd1 vssd1 vccd1 vccd1 _04202_ sky130_fd_sc_hd__mux2_1
XFILLER_0_157_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07484__A2 net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_145_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07211_ net1170 team_03_WB.instance_to_wrap.core.register_file.registers_state\[722\]
+ net756 team_03_WB.instance_to_wrap.core.register_file.registers_state\[754\] net740
+ vssd1 vssd1 vccd1 vccd1 _03153_ sky130_fd_sc_hd__o221a_1
XFILLER_0_27_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08191_ net1217 _04131_ _04132_ vssd1 vssd1 vccd1 vccd1 _04133_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_116_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11568__B2 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11511__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07142_ net1104 team_03_WB.instance_to_wrap.core.register_file.registers_state\[160\]
+ net902 vssd1 vssd1 vccd1 vccd1 _03084_ sky130_fd_sc_hd__or3_1
XANTENNA__07236__A2 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_742 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07641__C1 net1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07073_ _03011_ _03014_ net818 vssd1 vssd1 vccd1 vccd1 _03015_ sky130_fd_sc_hd__o21a_1
XFILLER_0_125_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07784__X _03726_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_2286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08197__B1 net995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_1004 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10543__A2 net1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11740__A1 net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07975_ net1203 team_03_WB.instance_to_wrap.core.register_file.registers_state\[464\]
+ vssd1 vssd1 vccd1 vccd1 _03917_ sky130_fd_sc_hd__or2_1
XANTENNA__08121__A net1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_143_3320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout383_A net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09714_ _05073_ _05586_ _05655_ vssd1 vssd1 vccd1 vccd1 _05656_ sky130_fd_sc_hd__a21bo_1
X_06926_ net1193 team_03_WB.instance_to_wrap.core.register_file.registers_state\[484\]
+ net886 _02867_ vssd1 vssd1 vccd1 vccd1 _02868_ sky130_fd_sc_hd__a31o_1
XANTENNA__07960__A net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09161__A2 net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09645_ _05552_ _05586_ net573 vssd1 vssd1 vccd1 vccd1 _05587_ sky130_fd_sc_hd__mux2_2
X_06857_ team_03_WB.instance_to_wrap.core.control_logic.instruction\[3\] team_03_WB.instance_to_wrap.core.control_logic.instruction\[2\]
+ team_03_WB.instance_to_wrap.core.control_logic.instruction\[1\] team_03_WB.instance_to_wrap.core.control_logic.instruction\[0\]
+ vssd1 vssd1 vccd1 vccd1 _02799_ sky130_fd_sc_hd__and4b_4
XANTENNA_fanout550_A net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07172__A1 net1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout269_X net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout648_A net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09576_ net581 _05504_ _05505_ _05516_ vssd1 vssd1 vccd1 vccd1 _05518_ sky130_fd_sc_hd__a31o_1
XFILLER_0_78_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_69_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10059__A1 net28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08527_ net1227 team_03_WB.instance_to_wrap.core.register_file.registers_state\[351\]
+ net952 team_03_WB.instance_to_wrap.core.register_file.registers_state\[383\] net1070
+ vssd1 vssd1 vccd1 vccd1 _04469_ sky130_fd_sc_hd__o221a_1
XANTENNA__11256__B1 net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1080_X net1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout815_A net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1178_X net1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07959__X _03901_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08458_ net871 _04396_ _04399_ _04393_ vssd1 vssd1 vccd1 vccd1 _04400_ sky130_fd_sc_hd__a31o_1
XFILLER_0_92_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08672__A1 net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07409_ _03341_ _03350_ net717 _03333_ vssd1 vssd1 vccd1 vccd1 _03351_ sky130_fd_sc_hd__a2bb2o_4
XTAP_TAPCELL_ROW_137_3179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout603_X net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08389_ net1245 team_03_WB.instance_to_wrap.core.register_file.registers_state\[89\]
+ net989 team_03_WB.instance_to_wrap.core.register_file.registers_state\[121\] net931
+ vssd1 vssd1 vccd1 vccd1 _04331_ sky130_fd_sc_hd__o221a_1
XFILLER_0_151_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10420_ team_03_WB.instance_to_wrap.core.pc.current_pc\[11\] _06139_ vssd1 vssd1
+ vccd1 vccd1 _06242_ sky130_fd_sc_hd__xor2_1
XANTENNA__13202__A net1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09621__B1 _05562_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_230 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_2732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_2743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10351_ team_03_WB.instance_to_wrap.core.pc.current_pc\[24\] _06185_ net680 vssd1
+ vssd1 vccd1 vccd1 _02658_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_167_3810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13070_ net1310 vssd1 vssd1 vccd1 vccd1 _00834_ sky130_fd_sc_hd__inv_2
X_10282_ _03313_ _05972_ vssd1 vssd1 vccd1 vccd1 _06124_ sky130_fd_sc_hd__nand2_1
XANTENNA__08730__S net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout972_X net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1116 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08188__B1 net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12021_ net618 _06582_ net451 net359 net2061 vssd1 vssd1 vccd1 vccd1 _01524_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_163_3718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10534__A2 net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11731__A1 net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07935__B1 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_163_3729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09127__A net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07573__C net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08031__A net1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout560 _03063_ vssd1 vssd1 vccd1 vccd1 net560 sky130_fd_sc_hd__buf_2
Xfanout571 net572 vssd1 vssd1 vccd1 vccd1 net571 sky130_fd_sc_hd__clkbuf_2
Xfanout582 _02950_ vssd1 vssd1 vccd1 vccd1 net582 sky130_fd_sc_hd__buf_4
X_13972_ clknet_leaf_133_wb_clk_i _01736_ _00337_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[326\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11495__A0 _06616_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12923_ net1361 vssd1 vssd1 vccd1 vccd1 _00687_ sky130_fd_sc_hd__inv_2
XFILLER_0_38_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12854_ net1258 vssd1 vssd1 vccd1 vccd1 _00618_ sky130_fd_sc_hd__inv_2
XFILLER_0_38_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12039__A2 net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11805_ net2602 _06631_ net330 vssd1 vssd1 vccd1 vccd1 _01733_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12785_ net1274 vssd1 vssd1 vccd1 vccd1 _00549_ sky130_fd_sc_hd__inv_2
XFILLER_0_173_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14524_ clknet_leaf_150_wb_clk_i _02288_ _00889_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[878\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_139_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11736_ net597 net265 net469 _06808_ net2189 vssd1 vssd1 vccd1 vccd1 _01800_ sky130_fd_sc_hd__a32o_1
XANTENNA__08905__S net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_25_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14455_ clknet_leaf_111_wb_clk_i _02219_ _00820_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[809\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07871__C1 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11667_ net2446 _06519_ net343 vssd1 vssd1 vccd1 vccd1 _01866_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11331__S net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13112__A net1380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13406_ net1424 vssd1 vssd1 vccd1 vccd1 _01170_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10618_ net2231 team_03_WB.instance_to_wrap.CPU_DAT_O\[11\] net842 vssd1 vssd1 vccd1
+ vccd1 _02510_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08415__A1 net1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_1020 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11598_ net296 net2403 net450 vssd1 vssd1 vccd1 vccd1 _01931_ sky130_fd_sc_hd__mux2_1
X_14386_ clknet_leaf_164_wb_clk_i _02150_ _00751_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[740\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10549_ net1142 team_03_WB.instance_to_wrap.core.d_hit _02837_ vssd1 vssd1 vccd1
+ vccd1 _06292_ sky130_fd_sc_hd__nor3_4
X_13337_ net1334 vssd1 vssd1 vccd1 vccd1 _01101_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11970__A1 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13268_ net1308 vssd1 vssd1 vccd1 vccd1 _01032_ sky130_fd_sc_hd__inv_2
X_15007_ clknet_leaf_52_wb_clk_i net55 _01372_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11567__A net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12219_ net1626 vssd1 vssd1 vccd1 vccd1 _01438_ sky130_fd_sc_hd__clkbuf_1
X_13199_ net1339 vssd1 vssd1 vccd1 vccd1 _00963_ sky130_fd_sc_hd__inv_2
XANTENNA__07077__S1 net1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10525__A2 net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11722__A1 _06454_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10902__C net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07760_ net1098 team_03_WB.instance_to_wrap.core.register_file.registers_state\[652\]
+ vssd1 vssd1 vccd1 vccd1 _03702_ sky130_fd_sc_hd__and2_1
XFILLER_0_47_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09679__B1 net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07691_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[830\] net767
+ net1041 vssd1 vssd1 vccd1 vccd1 _03633_ sky130_fd_sc_hd__o21a_1
XANTENNA__12398__A net1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09430_ net550 _04863_ _05042_ vssd1 vssd1 vccd1 vccd1 _05372_ sky130_fd_sc_hd__o21ba_1
XANTENNA__11506__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09361_ _05294_ _05298_ _05293_ vssd1 vssd1 vccd1 vccd1 _05303_ sky130_fd_sc_hd__o21a_1
XANTENNA__11238__B1 net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09203__C _05144_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_19_wb_clk_i clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_19_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_08312_ net1242 team_03_WB.instance_to_wrap.core.register_file.registers_state\[600\]
+ net985 team_03_WB.instance_to_wrap.core.register_file.registers_state\[632\] net928
+ vssd1 vssd1 vccd1 vccd1 _04254_ sky130_fd_sc_hd__o221a_1
X_09292_ _04893_ _05219_ _05215_ _04953_ vssd1 vssd1 vccd1 vccd1 _05234_ sky130_fd_sc_hd__a211o_1
XFILLER_0_145_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08243_ net1226 team_03_WB.instance_to_wrap.core.register_file.registers_state\[210\]
+ net950 team_03_WB.instance_to_wrap.core.register_file.registers_state\[242\] net934
+ vssd1 vssd1 vccd1 vccd1 _04185_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_43_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_644 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_172_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_2326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08174_ net1061 _04112_ _04115_ net1211 vssd1 vssd1 vccd1 vccd1 _04116_ sky130_fd_sc_hd__a211o_1
XANTENNA_clkbuf_leaf_13_wb_clk_i_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_2337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08116__A net1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07020__A net1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11410__A0 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07125_ net1198 team_03_WB.instance_to_wrap.core.register_file.registers_state\[544\]
+ net885 vssd1 vssd1 vccd1 vccd1 _03067_ sky130_fd_sc_hd__and3_1
XFILLER_0_160_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_132_3076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_3087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11961__A1 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1138_A net1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07056_ _02996_ _02997_ vssd1 vssd1 vccd1 vccd1 _02998_ sky130_fd_sc_hd__and2_1
Xoutput130 net130 vssd1 vssd1 vccd1 vccd1 ADR_O[5] sky130_fd_sc_hd__clkbuf_4
Xoutput141 net141 vssd1 vssd1 vccd1 vccd1 DAT_O[14] sky130_fd_sc_hd__buf_2
XANTENNA_fanout598_A net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput152 net152 vssd1 vssd1 vccd1 vccd1 DAT_O[24] sky130_fd_sc_hd__buf_2
XANTENNA__11477__A net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput163 net163 vssd1 vssd1 vccd1 vccd1 DAT_O[5] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_110_2640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput174 net174 vssd1 vssd1 vccd1 vccd1 gpio_oeb[0] sky130_fd_sc_hd__buf_2
XANTENNA__12072__S net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11908__C _06463_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10516__A2 net1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput185 net185 vssd1 vssd1 vccd1 vccd1 gpio_oeb[20] sky130_fd_sc_hd__buf_2
XANTENNA_fanout1305_A net1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11713__A1 _06413_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput196 net196 vssd1 vssd1 vccd1 vccd1 gpio_oeb[31] sky130_fd_sc_hd__clkbuf_4
XANTENNA__11196__B net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout765_A net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout386_X net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07958_ net721 _03899_ _03883_ _03882_ vssd1 vssd1 vccd1 vccd1 _03900_ sky130_fd_sc_hd__o2bb2a_4
X_06909_ net1196 net883 vssd1 vssd1 vccd1 vccd1 _02851_ sky130_fd_sc_hd__nand2_4
XANTENNA__10819__A3 net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout932_A _04088_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07889_ net1091 team_03_WB.instance_to_wrap.core.register_file.registers_state\[207\]
+ net794 team_03_WB.instance_to_wrap.core.register_file.registers_state\[239\] net729
+ vssd1 vssd1 vccd1 vccd1 _03831_ sky130_fd_sc_hd__a221o_1
XFILLER_0_98_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08342__B1 net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1295_X net1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11416__S net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_959 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_2591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09628_ _05102_ _05104_ net564 vssd1 vssd1 vccd1 vccd1 _05570_ sky130_fd_sc_hd__a21o_1
XFILLER_0_69_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11643__C net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_167_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11229__A0 _06536_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_52_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09559_ _05302_ _05305_ _05187_ vssd1 vssd1 vccd1 vccd1 _05501_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout720_X net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_514 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout818_X net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_368 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12570_ net1379 vssd1 vssd1 vccd1 vccd1 _00334_ sky130_fd_sc_hd__inv_2
XANTENNA__07448__A2 net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08645__A1 net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08952__C _04893_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_156_3577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_156_3588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11521_ _06381_ net650 _06634_ _06394_ vssd1 vssd1 vccd1 vccd1 _06779_ sky130_fd_sc_hd__or4b_4
XFILLER_0_80_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_22_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14240_ clknet_leaf_191_wb_clk_i _02004_ _00605_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[594\]
+ sky130_fd_sc_hd__dfrtp_1
X_11452_ net651 _06577_ vssd1 vssd1 vccd1 vccd1 _06765_ sky130_fd_sc_hd__nor2_1
XFILLER_0_33_241 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10403_ _06227_ _06228_ team_03_WB.instance_to_wrap.core.pc.current_pc\[15\] net680
+ vssd1 vssd1 vccd1 vccd1 _02649_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__10204__A1 net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11401__A0 _06413_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14171_ clknet_leaf_122_wb_clk_i _01935_ _00536_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[525\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11383_ net713 _06527_ net697 vssd1 vssd1 vccd1 vccd1 _06744_ sky130_fd_sc_hd__and3_1
XANTENNA__09070__A1 net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12771__A net1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06959__A1 net1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11952__A1 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input61_A gpio_in[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10334_ net283 _06171_ vssd1 vssd1 vccd1 vccd1 _06172_ sky130_fd_sc_hd__nand2_1
XFILLER_0_150_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13122_ net1352 vssd1 vssd1 vccd1 vccd1 _00886_ sky130_fd_sc_hd__inv_2
XFILLER_0_108_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13053_ net1383 vssd1 vssd1 vccd1 vccd1 _00817_ sky130_fd_sc_hd__inv_2
XANTENNA__11387__A net1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10265_ _06089_ _06103_ _06106_ vssd1 vssd1 vccd1 vccd1 _06107_ sky130_fd_sc_hd__o21bai_2
XFILLER_0_30_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12004_ net263 _06756_ net467 net445 net2016 vssd1 vssd1 vccd1 vccd1 _01540_ sky130_fd_sc_hd__a32o_1
Xfanout1300 net1301 vssd1 vssd1 vccd1 vccd1 net1300 sky130_fd_sc_hd__buf_4
Xfanout1311 net1312 vssd1 vssd1 vccd1 vccd1 net1311 sky130_fd_sc_hd__buf_4
Xfanout1322 net1324 vssd1 vssd1 vccd1 vccd1 net1322 sky130_fd_sc_hd__buf_4
X_10196_ _04679_ _05950_ vssd1 vssd1 vccd1 vccd1 _06038_ sky130_fd_sc_hd__nand2_1
Xfanout1333 net1335 vssd1 vssd1 vccd1 vccd1 net1333 sky130_fd_sc_hd__buf_4
XANTENNA__07384__A1 net1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1344 net1346 vssd1 vssd1 vccd1 vccd1 net1344 sky130_fd_sc_hd__buf_2
XANTENNA__11180__A2 net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1355 net1357 vssd1 vssd1 vccd1 vccd1 net1355 sky130_fd_sc_hd__buf_4
Xfanout1366 net1367 vssd1 vssd1 vccd1 vccd1 net1366 sky130_fd_sc_hd__buf_4
XANTENNA_clkbuf_leaf_91_wb_clk_i_A clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout1377 net1381 vssd1 vssd1 vccd1 vccd1 net1377 sky130_fd_sc_hd__buf_4
XFILLER_0_17_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08696__A net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1388 net1389 vssd1 vssd1 vccd1 vccd1 net1388 sky130_fd_sc_hd__buf_4
Xfanout390 _06778_ vssd1 vssd1 vccd1 vccd1 net390 sky130_fd_sc_hd__buf_8
Xfanout1399 net1401 vssd1 vssd1 vccd1 vccd1 net1399 sky130_fd_sc_hd__buf_4
X_13955_ clknet_leaf_31_wb_clk_i _01719_ _00320_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[309\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_17_68 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07136__A1 net1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06928__B net1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11326__S net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12906_ net1280 vssd1 vssd1 vccd1 vccd1 _00670_ sky130_fd_sc_hd__inv_2
XFILLER_0_158_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13886_ clknet_leaf_120_wb_clk_i _01650_ _00251_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[240\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12837_ net1349 vssd1 vssd1 vccd1 vccd1 _00601_ sky130_fd_sc_hd__inv_2
XANTENNA__12946__A net1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08636__A1 net1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1052 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08097__C1 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12768_ net1402 vssd1 vssd1 vccd1 vccd1 _00532_ sky130_fd_sc_hd__inv_2
XFILLER_0_33_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14507_ clknet_leaf_45_wb_clk_i _02271_ _00872_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[861\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_44_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11640__B1 net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11719_ net1831 net301 net335 vssd1 vssd1 vccd1 vccd1 _01817_ sky130_fd_sc_hd__mux2_1
XFILLER_0_127_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_906 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12699_ net1361 vssd1 vssd1 vccd1 vccd1 _00463_ sky130_fd_sc_hd__inv_2
XFILLER_0_140_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_142_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14438_ clknet_leaf_72_wb_clk_i _02202_ _00803_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[792\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput10 DAT_I[17] vssd1 vssd1 vccd1 vccd1 net10 sky130_fd_sc_hd__buf_1
Xinput21 DAT_I[27] vssd1 vssd1 vccd1 vccd1 net21 sky130_fd_sc_hd__buf_1
XFILLER_0_141_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput32 DAT_I[8] vssd1 vssd1 vccd1 vccd1 net32 sky130_fd_sc_hd__clkbuf_1
Xinput43 gpio_in[18] vssd1 vssd1 vccd1 vccd1 net43 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11996__S net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput54 gpio_in[29] vssd1 vssd1 vccd1 vccd1 net54 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_142_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput65 gpio_in[9] vssd1 vssd1 vccd1 vccd1 net65 sky130_fd_sc_hd__clkbuf_1
X_14369_ clknet_leaf_180_wb_clk_i _02133_ _00734_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[723\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold805 team_03_WB.instance_to_wrap.core.register_file.registers_state\[253\] vssd1
+ vssd1 vccd1 vccd1 net2298 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold816 team_03_WB.instance_to_wrap.core.register_file.registers_state\[526\] vssd1
+ vssd1 vccd1 vccd1 net2309 sky130_fd_sc_hd__dlygate4sd3_1
Xinput76 wbs_adr_i[18] vssd1 vssd1 vccd1 vccd1 net76 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_959 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11943__A1 net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput87 wbs_adr_i[28] vssd1 vssd1 vccd1 vccd1 net87 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_141_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_137_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_137_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xhold827 team_03_WB.instance_to_wrap.core.register_file.registers_state\[618\] vssd1
+ vssd1 vccd1 vccd1 net2320 sky130_fd_sc_hd__dlygate4sd3_1
Xinput98 wbs_adr_i[9] vssd1 vssd1 vccd1 vccd1 net98 sky130_fd_sc_hd__clkbuf_1
Xhold838 team_03_WB.instance_to_wrap.core.register_file.registers_state\[79\] vssd1
+ vssd1 vccd1 vccd1 net2331 sky130_fd_sc_hd__dlygate4sd3_1
Xhold849 team_03_WB.instance_to_wrap.core.register_file.registers_state\[798\] vssd1
+ vssd1 vccd1 vccd1 net2342 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_2223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_1051 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_2234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11297__A net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08930_ net1046 team_03_WB.instance_to_wrap.core.register_file.registers_state\[331\]
+ net997 team_03_WB.instance_to_wrap.core.register_file.registers_state\[363\] net1214
+ vssd1 vssd1 vccd1 vccd1 _04872_ sky130_fd_sc_hd__a221o_1
XFILLER_0_23_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_wire354_X net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09364__A2 _05281_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08861_ net1056 team_03_WB.instance_to_wrap.core.register_file.registers_state\[960\]
+ net1009 team_03_WB.instance_to_wrap.core.register_file.registers_state\[992\] net1078
+ vssd1 vssd1 vccd1 vccd1 _04803_ sky130_fd_sc_hd__a221o_1
XANTENNA__07375__A1 net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08572__B1 net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07812_ _03749_ _03753_ _03752_ net1119 vssd1 vssd1 vccd1 vccd1 _03754_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__07914__A3 net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08792_ net925 _04732_ _04733_ vssd1 vssd1 vccd1 vccd1 _04734_ sky130_fd_sc_hd__a21o_1
XFILLER_0_93_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07743_ net1098 net898 team_03_WB.instance_to_wrap.core.register_file.registers_state\[140\]
+ vssd1 vssd1 vccd1 vccd1 _03685_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_88_2174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07127__A1 net1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_2185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07127__B2 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_96 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07674_ net1178 team_03_WB.instance_to_wrap.core.register_file.registers_state\[478\]
+ net771 team_03_WB.instance_to_wrap.core.register_file.registers_state\[510\] net1151
+ vssd1 vssd1 vccd1 vccd1 _03616_ sky130_fd_sc_hd__o221a_1
XFILLER_0_95_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09413_ net573 _04832_ vssd1 vssd1 vccd1 vccd1 _05355_ sky130_fd_sc_hd__nor2_1
XANTENNA__07015__A net1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12856__A net1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout346_A _06804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1088_A net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_165_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09344_ _03170_ _03989_ _05149_ net607 vssd1 vssd1 vccd1 vccd1 _05286_ sky130_fd_sc_hd__a31o_1
XANTENNA__08627__A1 net1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08545__S net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06854__A net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10434__A1 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09230__A _04532_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09275_ _04954_ _05215_ vssd1 vssd1 vccd1 vccd1 _05217_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_8_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07835__C1 net1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11631__B1 net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_163 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12067__S net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_134_3127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout513_A net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_136_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_28_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1255_A net1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08226_ net1233 team_03_WB.instance_to_wrap.core.register_file.registers_state\[849\]
+ net961 team_03_WB.instance_to_wrap.core.register_file.registers_state\[881\] net1217
+ vssd1 vssd1 vccd1 vccd1 _04168_ sky130_fd_sc_hd__o221a_1
XANTENNA__10095__B _05453_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_160_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_758 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_151_3474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08157_ net1230 team_03_WB.instance_to_wrap.core.register_file.registers_state\[468\]
+ net961 team_03_WB.instance_to_wrap.core.register_file.registers_state\[500\] net1210
+ vssd1 vssd1 vccd1 vccd1 _04099_ sky130_fd_sc_hd__o221a_1
XFILLER_0_71_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09052__A1 net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout301_X net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_151_3485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1422_A net1436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1043_X net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10737__A2 net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07108_ net1100 team_03_WB.instance_to_wrap.core.register_file.registers_state\[65\]
+ net799 team_03_WB.instance_to_wrap.core.register_file.registers_state\[97\] net747
+ vssd1 vssd1 vccd1 vccd1 _03050_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_31_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08088_ net1152 net1019 net684 vssd1 vssd1 vccd1 vccd1 _04030_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_28_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout882_A net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_266 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07039_ net815 _02979_ _02980_ vssd1 vssd1 vccd1 vccd1 _02981_ sky130_fd_sc_hd__and3_1
XFILLER_0_12_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_140_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1210_X net1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10050_ net6 net1038 net910 net1715 vssd1 vssd1 vccd1 vccd1 _02681_ sky130_fd_sc_hd__o22a_1
XANTENNA__08012__C1 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08789__S1 net1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11698__B1 net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout670_X net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout768_X net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout935_X net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07118__B2 net1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13740_ clknet_leaf_19_wb_clk_i _01504_ _00105_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[94\]
+ sky130_fd_sc_hd__dfrtp_1
X_10952_ net689 _05768_ vssd1 vssd1 vccd1 vccd1 _06535_ sky130_fd_sc_hd__nand2_1
XANTENNA__08410__S0 net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11373__C net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_175_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_74_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_158_3617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_158_3628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11870__A0 _06536_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13671_ clknet_leaf_109_wb_clk_i _01435_ _00036_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_123_2897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10883_ net838 _06478_ vssd1 vssd1 vccd1 vccd1 _06479_ sky130_fd_sc_hd__nor2_4
XFILLER_0_128_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_168_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08079__C1 net1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12622_ net1305 vssd1 vssd1 vccd1 vccd1 _00386_ sky130_fd_sc_hd__inv_2
XFILLER_0_94_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08618__A1 net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12553_ net1260 vssd1 vssd1 vccd1 vccd1 _00317_ sky130_fd_sc_hd__inv_2
XANTENNA__11622__B1 net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08094__A2 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10976__A2 _05142_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11504_ _06622_ net2439 net391 vssd1 vssd1 vccd1 vccd1 _02002_ sky130_fd_sc_hd__mux2_1
X_12484_ net1376 vssd1 vssd1 vccd1 vccd1 _00248_ sky130_fd_sc_hd__inv_2
XFILLER_0_34_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14223_ clknet_leaf_136_wb_clk_i _01987_ _00588_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[577\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11435_ net1250 _06449_ net650 net701 vssd1 vssd1 vccd1 vccd1 _06757_ sky130_fd_sc_hd__or4_1
XFILLER_0_34_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07054__B1 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07595__A net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14154_ clknet_leaf_2_wb_clk_i _01918_ _00519_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[508\]
+ sky130_fd_sc_hd__dfrtp_1
X_11366_ net501 net630 _06735_ net401 net1969 vssd1 vssd1 vccd1 vccd1 _02097_ sky130_fd_sc_hd__a32o_1
XANTENNA__08043__X _03985_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10317_ team_03_WB.instance_to_wrap.core.pc.current_pc\[30\] _06152_ vssd1 vssd1
+ vccd1 vccd1 _06158_ sky130_fd_sc_hd__or2_1
X_13105_ net1268 vssd1 vssd1 vccd1 vccd1 _00869_ sky130_fd_sc_hd__inv_2
X_11297_ net715 _06557_ net830 vssd1 vssd1 vccd1 vccd1 _06716_ sky130_fd_sc_hd__and3_1
XFILLER_0_81_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14085_ clknet_leaf_15_wb_clk_i _01849_ _00450_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[439\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_120_986 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10248_ _04294_ team_03_WB.instance_to_wrap.core.pc.current_pc\[21\] net673 vssd1
+ vssd1 vccd1 vccd1 _06090_ sky130_fd_sc_hd__mux2_1
X_13036_ net1314 vssd1 vssd1 vccd1 vccd1 _00800_ sky130_fd_sc_hd__inv_2
XANTENNA__11689__B1 net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11267__D net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11153__A2 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1130 _02785_ vssd1 vssd1 vccd1 vccd1 net1130 sky130_fd_sc_hd__buf_4
XFILLER_0_119_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1141 _02784_ vssd1 vssd1 vccd1 vccd1 net1141 sky130_fd_sc_hd__buf_6
XFILLER_0_28_67 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10179_ _06020_ vssd1 vssd1 vccd1 vccd1 _06021_ sky130_fd_sc_hd__inv_2
Xfanout1152 net1159 vssd1 vssd1 vccd1 vccd1 net1152 sky130_fd_sc_hd__clkbuf_8
Xfanout1163 net1169 vssd1 vssd1 vccd1 vccd1 net1163 sky130_fd_sc_hd__buf_4
XANTENNA__10900__A2 _05659_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1174 net1180 vssd1 vssd1 vccd1 vccd1 net1174 sky130_fd_sc_hd__buf_2
Xfanout1185 net1190 vssd1 vssd1 vccd1 vccd1 net1185 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09315__A _02938_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14929__Q team_03_WB.instance_to_wrap.CPU_DAT_O\[16\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__07761__C net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1196 net1199 vssd1 vssd1 vccd1 vccd1 net1196 sky130_fd_sc_hd__buf_4
X_14987_ clknet_leaf_66_wb_clk_i net35 _01352_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_135_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13938_ clknet_leaf_117_wb_clk_i _01702_ _00303_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[292\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11283__C net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11861__A0 net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09969__B net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13869_ clknet_leaf_189_wb_clk_i _01633_ _00234_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[223\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_83_2082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08609__A1 net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07390_ _03328_ _03329_ _03330_ _03331_ net817 vssd1 vssd1 vccd1 vccd1 _03332_ sky130_fd_sc_hd__a221o_1
XFILLER_0_173_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_366 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_675 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11613__B1 net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10196__A _04679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_40_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_151_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09060_ net1047 team_03_WB.instance_to_wrap.core.register_file.registers_state\[687\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[655\] net998 net939
+ vssd1 vssd1 vccd1 vccd1 _05002_ sky130_fd_sc_hd__o221a_1
XFILLER_0_127_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08490__C1 net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_154_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08011_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[945\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[913\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[817\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[785\]
+ net765 net1125 vssd1 vssd1 vccd1 vccd1 _03953_ sky130_fd_sc_hd__mux4_1
XFILLER_0_25_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_712 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09034__A1 net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_66 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold602 team_03_WB.instance_to_wrap.core.register_file.registers_state\[342\] vssd1
+ vssd1 vccd1 vccd1 net2095 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold613 team_03_WB.instance_to_wrap.core.register_file.registers_state\[414\] vssd1
+ vssd1 vccd1 vccd1 net2106 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold624 team_03_WB.instance_to_wrap.core.register_file.registers_state\[122\] vssd1
+ vssd1 vccd1 vccd1 net2117 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08242__C1 net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold635 team_03_WB.instance_to_wrap.core.register_file.registers_state\[132\] vssd1
+ vssd1 vccd1 vccd1 net2128 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold646 team_03_WB.instance_to_wrap.core.register_file.registers_state\[259\] vssd1
+ vssd1 vccd1 vccd1 net2139 sky130_fd_sc_hd__dlygate4sd3_1
Xhold657 team_03_WB.instance_to_wrap.core.register_file.registers_state\[124\] vssd1
+ vssd1 vccd1 vccd1 net2150 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08793__B1 net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11392__A2 net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold668 team_03_WB.instance_to_wrap.core.register_file.registers_state\[418\] vssd1
+ vssd1 vccd1 vccd1 net2161 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold679 team_03_WB.instance_to_wrap.core.register_file.registers_state\[106\] vssd1
+ vssd1 vccd1 vccd1 net2172 sky130_fd_sc_hd__dlygate4sd3_1
X_09962_ _05885_ net1706 net291 vssd1 vssd1 vccd1 vccd1 _02746_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_38_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08913_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[812\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[780\]
+ net979 vssd1 vssd1 vccd1 vccd1 _04855_ sky130_fd_sc_hd__mux2_1
X_09893_ _04031_ _04323_ net538 vssd1 vssd1 vccd1 vccd1 _05835_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07348__A1 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout296_A _06513_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08844_ net865 _04784_ _04785_ vssd1 vssd1 vccd1 vccd1 _04786_ sky130_fd_sc_hd__and3_1
XANTENNA__07443__S1 net1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1052 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06849__A team_03_WB.instance_to_wrap.core.decoder.inst\[13\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1003_A net1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14839__Q net103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08775_ _04715_ _04716_ net857 vssd1 vssd1 vccd1 vccd1 _04717_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout463_A net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_34_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_34_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_170_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07726_ _03665_ _03667_ net1166 vssd1 vssd1 vccd1 vccd1 _03668_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_68_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10655__A1 team_03_WB.instance_to_wrap.CPU_DAT_O\[6\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11852__A0 net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07657_ net1139 _03589_ _03593_ _03596_ _03598_ vssd1 vssd1 vccd1 vccd1 _03599_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_0_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout630_A net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_817 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07520__A1 net1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout728_A net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout349_X net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_2447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07588_ net1205 team_03_WB.instance_to_wrap.core.register_file.registers_state\[57\]
+ net886 vssd1 vssd1 vccd1 vccd1 _03530_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_101_2458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10818__B _05541_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10407__A1 net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11604__A0 net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_153_3514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09327_ _05265_ _05267_ _05249_ _05253_ vssd1 vssd1 vccd1 vccd1 _05269_ sky130_fd_sc_hd__a211o_1
XFILLER_0_47_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_153_3525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout516_X net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1160_X net1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_703 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07284__B1 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09258_ _03866_ _05199_ vssd1 vssd1 vccd1 vccd1 _05200_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_7_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_170_3861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_170_3872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08209_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[49\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[17\]
+ net960 vssd1 vssd1 vccd1 vccd1 _04151_ sky130_fd_sc_hd__mux2_1
X_09189_ net434 net429 _04565_ net545 vssd1 vssd1 vccd1 vccd1 _05131_ sky130_fd_sc_hd__o31a_1
XFILLER_0_133_566 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11907__A1 net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13210__A net1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11220_ _06456_ _06503_ vssd1 vssd1 vccd1 vccd1 _06682_ sky130_fd_sc_hd__nor2_1
XANTENNA__07036__B1 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_542 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07587__A1 _03528_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_238 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout885_X net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08784__B1 net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11151_ net493 net647 _06652_ net412 net1723 vssd1 vssd1 vccd1 vccd1 _02229_ sky130_fd_sc_hd__a32o_1
XFILLER_0_101_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10591__B1 net1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10102_ net304 net303 vssd1 vssd1 vccd1 vccd1 _05946_ sky130_fd_sc_hd__nand2_1
X_11082_ net833 _06442_ vssd1 vssd1 vccd1 vccd1 _06619_ sky130_fd_sc_hd__and2_2
XANTENNA__07339__A1 net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11135__A2 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14910_ clknet_leaf_55_wb_clk_i _00004_ _01275_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.ru.state\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_10033_ net25 net1039 _05906_ net2780 vssd1 vssd1 vccd1 vccd1 _02698_ sky130_fd_sc_hd__a22o_1
XFILLER_0_41_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09135__A net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14841_ clknet_leaf_87_wb_clk_i _02605_ _01206_ vssd1 vssd1 vccd1 vccd1 net125 sky130_fd_sc_hd__dfrtp_2
XANTENNA_input24_A DAT_I[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12096__B1 net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14772_ clknet_leaf_103_wb_clk_i _02536_ _01137_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_I\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_11984_ net300 net2456 net446 vssd1 vssd1 vccd1 vccd1 _01560_ sky130_fd_sc_hd__mux2_1
XFILLER_0_169_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11843__A0 net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13723_ clknet_leaf_145_wb_clk_i _01487_ _00088_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[77\]
+ sky130_fd_sc_hd__dfrtp_1
X_10935_ net314 _05846_ net316 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[7\]
+ vssd1 vssd1 vccd1 vccd1 _06521_ sky130_fd_sc_hd__o31a_1
XFILLER_0_129_817 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07511__A1 net1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11604__S net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13654_ clknet_leaf_153_wb_clk_i _01418_ _00019_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10866_ net493 _06454_ net596 net518 net2014 vssd1 vssd1 vccd1 vccd1 _02326_ sky130_fd_sc_hd__a32o_1
XFILLER_0_112_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12605_ net1389 vssd1 vssd1 vccd1 vccd1 _00369_ sky130_fd_sc_hd__inv_2
XFILLER_0_94_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13585_ net1404 vssd1 vssd1 vccd1 vccd1 _01349_ sky130_fd_sc_hd__inv_2
XFILLER_0_171_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10797_ net687 _05429_ vssd1 vssd1 vccd1 vccd1 _06406_ sky130_fd_sc_hd__and2_1
XFILLER_0_143_308 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07275__B1 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_147_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12536_ net1375 vssd1 vssd1 vccd1 vccd1 _00300_ sky130_fd_sc_hd__inv_2
XANTENNA__08913__S net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_151_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12467_ net1255 vssd1 vssd1 vccd1 vccd1 _00231_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_144_Right_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13120__A net1402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14206_ clknet_leaf_118_wb_clk_i _01970_ _00571_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[560\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_151_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09567__A2 _04235_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12020__B1 net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11418_ net298 net2671 net398 vssd1 vssd1 vccd1 vccd1 _02063_ sky130_fd_sc_hd__mux2_1
XANTENNA__08224__C1 net1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12398_ net1270 vssd1 vssd1 vccd1 vccd1 _00162_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11374__A2 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08775__B1 net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14137_ clknet_leaf_156_wb_clk_i _01901_ _00502_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[491\]
+ sky130_fd_sc_hd__dfrtp_1
X_11349_ net1247 net837 _06438_ net668 vssd1 vssd1 vccd1 vccd1 _06727_ sky130_fd_sc_hd__and4_1
XANTENNA__10582__B1 net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14068_ clknet_leaf_133_wb_clk_i _01832_ _00433_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[422\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08527__B1 net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13019_ net1359 vssd1 vssd1 vccd1 vccd1 _00783_ sky130_fd_sc_hd__inv_2
X_06890_ team_03_WB.instance_to_wrap.core.decoder.inst\[12\] _02820_ vssd1 vssd1 vccd1
+ vccd1 _02832_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_33_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_21 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07117__X _03059_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12087__B1 net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08560_ net875 _04496_ _04501_ vssd1 vssd1 vccd1 vccd1 _04502_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_18_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10637__A1 team_03_WB.instance_to_wrap.CPU_DAT_O\[24\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_07511_ net1204 team_03_WB.instance_to_wrap.core.register_file.registers_state\[487\]
+ net885 _03452_ vssd1 vssd1 vccd1 vccd1 _03453_ sky130_fd_sc_hd__a31o_1
X_08491_ net945 _04431_ _04432_ vssd1 vssd1 vccd1 vccd1 _04433_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_18_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11834__B1 net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11514__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07442_ net1176 team_03_WB.instance_to_wrap.core.register_file.registers_state\[468\]
+ net764 team_03_WB.instance_to_wrap.core.register_file.registers_state\[500\] net1150
+ vssd1 vssd1 vccd1 vccd1 _03384_ sky130_fd_sc_hd__o221a_1
XFILLER_0_162_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07373_ net1084 net889 team_03_WB.instance_to_wrap.core.register_file.registers_state\[31\]
+ vssd1 vssd1 vccd1 vccd1 _03315_ sky130_fd_sc_hd__o21a_1
XFILLER_0_162_606 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08689__S0 net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09112_ net1066 _05052_ _05053_ vssd1 vssd1 vccd1 vccd1 _05054_ sky130_fd_sc_hd__a21o_1
Xclkbuf_leaf_152_wb_clk_i clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_152_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08463__C1 net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11062__B2 net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09043_ net433 net427 net590 vssd1 vssd1 vccd1 vccd1 _04985_ sky130_fd_sc_hd__nor3_1
XFILLER_0_115_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_167_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout309_A _05846_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13030__A net1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold410 _02624_ vssd1 vssd1 vccd1 vccd1 net1903 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_111_Right_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12011__B1 net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold421 team_03_WB.instance_to_wrap.core.register_file.registers_state\[289\] vssd1
+ vssd1 vccd1 vccd1 net1914 sky130_fd_sc_hd__dlygate4sd3_1
Xhold432 team_03_WB.instance_to_wrap.CPU_DAT_I\[27\] vssd1 vssd1 vccd1 vccd1 net1925
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07569__A1 net1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold443 team_03_WB.instance_to_wrap.core.register_file.registers_state\[55\] vssd1
+ vssd1 vccd1 vccd1 net1936 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold454 team_03_WB.instance_to_wrap.core.register_file.registers_state\[36\] vssd1
+ vssd1 vccd1 vccd1 net1947 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11188__C _06536_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold465 team_03_WB.instance_to_wrap.core.register_file.registers_state\[58\] vssd1
+ vssd1 vccd1 vccd1 net1958 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1120_A net1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_3015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10573__B1 net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold476 team_03_WB.instance_to_wrap.core.register_file.registers_state\[687\] vssd1
+ vssd1 vccd1 vccd1 net1969 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_3026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold487 team_03_WB.instance_to_wrap.core.register_file.registers_state\[701\] vssd1
+ vssd1 vccd1 vccd1 net1980 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1218_A net1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout901 net902 vssd1 vssd1 vccd1 vccd1 net901 sky130_fd_sc_hd__clkbuf_4
Xhold498 team_03_WB.instance_to_wrap.core.register_file.registers_state\[903\] vssd1
+ vssd1 vccd1 vccd1 net1991 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout912 net914 vssd1 vssd1 vccd1 vccd1 net912 sky130_fd_sc_hd__clkbuf_2
X_09945_ _03425_ net662 vssd1 vssd1 vccd1 vccd1 _05877_ sky130_fd_sc_hd__nor2_1
XANTENNA__09881__C _05821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout580_A _02992_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_1892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout923 _04088_ vssd1 vssd1 vccd1 vccd1 net923 sky130_fd_sc_hd__buf_2
Xfanout934 net936 vssd1 vssd1 vccd1 vccd1 net934 sky130_fd_sc_hd__buf_4
XANTENNA_fanout678_A net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout945 net948 vssd1 vssd1 vccd1 vccd1 net945 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout299_X net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout956 net974 vssd1 vssd1 vccd1 vccd1 net956 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_146_3373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09876_ net538 _05816_ net664 vssd1 vssd1 vccd1 vccd1 _05818_ sky130_fd_sc_hd__a21bo_1
Xfanout967 net969 vssd1 vssd1 vccd1 vccd1 net967 sky130_fd_sc_hd__clkbuf_2
Xhold1110 team_03_WB.instance_to_wrap.core.register_file.registers_state\[141\] vssd1
+ vssd1 vccd1 vccd1 net2603 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1006_X net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout978 net994 vssd1 vssd1 vccd1 vccd1 net978 sky130_fd_sc_hd__clkbuf_4
Xhold1121 team_03_WB.instance_to_wrap.core.register_file.registers_state\[154\] vssd1
+ vssd1 vccd1 vccd1 net2614 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout989 net990 vssd1 vssd1 vccd1 vccd1 net989 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_5_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1132 team_03_WB.instance_to_wrap.core.register_file.registers_state\[86\] vssd1
+ vssd1 vccd1 vccd1 net2625 sky130_fd_sc_hd__dlygate4sd3_1
X_08827_ net1208 _04761_ net848 vssd1 vssd1 vccd1 vccd1 _04769_ sky130_fd_sc_hd__a21o_1
Xhold1143 team_03_WB.instance_to_wrap.core.register_file.registers_state\[606\] vssd1
+ vssd1 vccd1 vccd1 net2636 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout845_A _06303_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1154 team_03_WB.instance_to_wrap.core.register_file.registers_state\[861\] vssd1
+ vssd1 vccd1 vccd1 net2647 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout466_X net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1165 team_03_WB.instance_to_wrap.core.register_file.registers_state\[843\] vssd1
+ vssd1 vccd1 vccd1 net2658 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1176 team_03_WB.instance_to_wrap.core.register_file.registers_state\[172\] vssd1
+ vssd1 vccd1 vccd1 net2669 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12078__B1 net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1187 team_03_WB.instance_to_wrap.core.register_file.registers_state\[616\] vssd1
+ vssd1 vccd1 vccd1 net2680 sky130_fd_sc_hd__dlygate4sd3_1
X_08758_ net1221 _04698_ _04699_ vssd1 vssd1 vccd1 vccd1 _04700_ sky130_fd_sc_hd__and3_1
Xhold1198 team_03_WB.instance_to_wrap.core.register_file.registers_state\[585\] vssd1
+ vssd1 vccd1 vccd1 net2691 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_135_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10628__A1 team_03_WB.instance_to_wrap.CPU_DAT_O\[1\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_07709_ net815 _03646_ _03647_ _03650_ vssd1 vssd1 vccd1 vccd1 _03651_ sky130_fd_sc_hd__o22a_1
XANTENNA__11825__B1 net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08689_ _04627_ _04628_ _04629_ _04630_ net862 net924 vssd1 vssd1 vccd1 vccd1 _04631_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout633_X net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_120_2834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_2845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10720_ net522 _06350_ _06351_ net527 net2089 vssd1 vssd1 vccd1 vccd1 _02455_ sky130_fd_sc_hd__a32o_1
XFILLER_0_49_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_172_3901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_172_3912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07203__A net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09246__A1 _03391_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10651_ team_03_WB.instance_to_wrap.core.decoder.inst\[10\] team_03_WB.instance_to_wrap.CPU_DAT_O\[10\]
+ net845 vssd1 vssd1 vccd1 vccd1 _02477_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout800_X net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13370_ net1321 vssd1 vssd1 vccd1 vccd1 _01134_ sky130_fd_sc_hd__inv_2
X_10582_ net1622 net532 net599 _03488_ vssd1 vssd1 vccd1 vccd1 _02541_ sky130_fd_sc_hd__a22o_1
XFILLER_0_134_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08454__C1 net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_987 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_544 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12321_ net1281 vssd1 vssd1 vccd1 vccd1 _00085_ sky130_fd_sc_hd__inv_2
XFILLER_0_35_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_2796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15040_ clknet_leaf_88_wb_clk_i _02760_ _01405_ vssd1 vssd1 vccd1 vccd1 net196 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_160_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09549__A2 _04267_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12252_ net1430 vssd1 vssd1 vccd1 vccd1 _00016_ sky130_fd_sc_hd__inv_2
XFILLER_0_50_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12002__B1 net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08757__B1 net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11356__A2 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11203_ net302 net2487 net488 vssd1 vssd1 vccd1 vccd1 _02205_ sky130_fd_sc_hd__mux2_1
XFILLER_0_142_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12183_ net1814 vssd1 vssd1 vccd1 vccd1 _02370_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__10564__B1 net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07655__S1 net1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1146 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11134_ net1044 net836 net278 net668 vssd1 vssd1 vccd1 vccd1 _06643_ sky130_fd_sc_hd__and4_1
XANTENNA__11395__A net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11065_ _06609_ net2377 net416 vssd1 vssd1 vccd1 vccd1 _02273_ sky130_fd_sc_hd__mux2_1
X_10016_ net98 net97 net69 net68 vssd1 vssd1 vccd1 vccd1 _05894_ sky130_fd_sc_hd__or4_1
XANTENNA_output228_A net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14824_ clknet_leaf_102_wb_clk_i net1712 _01189_ vssd1 vssd1 vccd1 vccd1 net144 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_116_37 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10619__A1 team_03_WB.instance_to_wrap.CPU_DAT_O\[10\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14755_ clknet_leaf_50_wb_clk_i net1829 _01120_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11816__B1 net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11842__B net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09485__A1 net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11967_ net637 _06744_ net470 net365 net2442 vssd1 vssd1 vccd1 vccd1 _01576_ sky130_fd_sc_hd__a32o_1
XANTENNA__09485__B2 net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12084__A3 net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11292__A1 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13706_ clknet_leaf_1_wb_clk_i _01470_ _00071_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[60\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13115__A net1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_2030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_934 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09312__B _05125_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10918_ team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[10\] net305 vssd1
+ vssd1 vccd1 vccd1 _06507_ sky130_fd_sc_hd__nand2_1
XANTENNA__07496__B1 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14686_ clknet_leaf_64_wb_clk_i _02450_ _01051_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.ADR_I\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11831__A3 net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11898_ net644 _06707_ net475 net374 net2065 vssd1 vssd1 vccd1 vccd1 _01643_ sky130_fd_sc_hd__a32o_1
XANTENNA__07113__A net1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13637_ net1426 vssd1 vssd1 vccd1 vccd1 _01401_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_157_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10849_ _06394_ _06447_ vssd1 vssd1 vccd1 vccd1 _06448_ sky130_fd_sc_hd__and2_1
XANTENNA__07248__B1 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_680 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08445__C1 net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_976 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13568_ net1433 vssd1 vssd1 vccd1 vccd1 _01332_ sky130_fd_sc_hd__inv_2
XFILLER_0_54_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08996__B1 net995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12519_ net1368 vssd1 vssd1 vccd1 vccd1 _00283_ sky130_fd_sc_hd__inv_2
XANTENNA__10474__A net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13499_ net1340 vssd1 vssd1 vccd1 vccd1 _01263_ sky130_fd_sc_hd__inv_2
XFILLER_0_41_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11289__B net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1079 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_140_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_3_2_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_2_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_67_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_160_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_35_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11898__A3 net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07783__A net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07991_ _02872_ _03931_ _03932_ _02870_ _03930_ vssd1 vssd1 vccd1 vccd1 _03933_ sky130_fd_sc_hd__o221a_1
XFILLER_0_10_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11509__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07971__A1 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09730_ _05669_ _05670_ net577 vssd1 vssd1 vccd1 vccd1 _05672_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_52_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06942_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[996\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[964\]
+ net776 vssd1 vssd1 vccd1 vccd1 _02884_ sky130_fd_sc_hd__mux2_1
XFILLER_0_158_1023 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_52_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10858__A1 team_03_WB.instance_to_wrap.core.decoder.inst\[10\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09661_ net575 _05527_ _05602_ vssd1 vssd1 vccd1 vccd1 _05603_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_119_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06873_ team_03_WB.instance_to_wrap.core.control_logic.instruction\[6\] team_03_WB.instance_to_wrap.core.control_logic.instruction\[5\]
+ _02807_ vssd1 vssd1 vccd1 vccd1 _02815_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_2_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08612_ net1245 team_03_WB.instance_to_wrap.core.register_file.registers_state\[133\]
+ net992 team_03_WB.instance_to_wrap.core.register_file.registers_state\[165\] net947
+ vssd1 vssd1 vccd1 vccd1 _04554_ sky130_fd_sc_hd__o221a_1
X_09592_ net575 _05533_ vssd1 vssd1 vccd1 vccd1 _05534_ sky130_fd_sc_hd__nor2_1
XFILLER_0_96_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_141_3270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09503__A net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08543_ net1229 team_03_WB.instance_to_wrap.core.register_file.registers_state\[606\]
+ net955 team_03_WB.instance_to_wrap.core.register_file.registers_state\[638\] net1070
+ vssd1 vssd1 vccd1 vccd1 _04485_ sky130_fd_sc_hd__o221a_1
XFILLER_0_148_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08474_ _04080_ _04415_ vssd1 vssd1 vccd1 vccd1 _04416_ sky130_fd_sc_hd__nor2_1
XFILLER_0_65_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11822__A3 net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07023__A net1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07425_ _03364_ _03366_ net1169 vssd1 vssd1 vccd1 vccd1 _03367_ sky130_fd_sc_hd__o21a_1
XFILLER_0_58_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11190__D net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1070_A net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12864__A net1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout426_A _04079_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10087__C _05706_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1168_A net1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07239__B1 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07356_ net1172 team_03_WB.instance_to_wrap.core.register_file.registers_state\[732\]
+ net759 team_03_WB.instance_to_wrap.core.register_file.registers_state\[764\] net739
+ vssd1 vssd1 vccd1 vccd1 _03298_ sky130_fd_sc_hd__o221a_1
XFILLER_0_33_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08987__B1 net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_2379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07287_ _03226_ _03228_ net813 vssd1 vssd1 vccd1 vccd1 _03229_ sky130_fd_sc_hd__a21o_1
XANTENNA__10384__A _06086_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1335_A net1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07169__S net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09026_ net1067 _04965_ _04966_ vssd1 vssd1 vccd1 vccd1 _04968_ sky130_fd_sc_hd__or3_1
XFILLER_0_20_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_1932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_1943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11338__A2 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout795_A _02850_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold240 net210 vssd1 vssd1 vccd1 vccd1 net1733 sky130_fd_sc_hd__dlygate4sd3_1
Xhold251 _02619_ vssd1 vssd1 vccd1 vccd1 net1744 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_148_3413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1123_X net1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_148_3424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold262 _02582_ vssd1 vssd1 vccd1 vccd1 net1755 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11889__A3 net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold273 _02627_ vssd1 vssd1 vccd1 vccd1 net1766 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_113_2693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold284 team_03_WB.instance_to_wrap.core.register_file.registers_state\[6\] vssd1
+ vssd1 vccd1 vccd1 net1777 sky130_fd_sc_hd__dlygate4sd3_1
Xhold295 team_03_WB.instance_to_wrap.core.register_file.registers_state\[898\] vssd1
+ vssd1 vccd1 vccd1 net1788 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout583_X net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout962_A net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07962__A1 net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout720 _02864_ vssd1 vssd1 vccd1 vccd1 net720 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_165_3760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11419__S net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout731 net733 vssd1 vssd1 vccd1 vccd1 net731 sky130_fd_sc_hd__buf_4
X_09928_ _05868_ net1776 net294 vssd1 vssd1 vccd1 vccd1 _02763_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_165_3771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout742 net755 vssd1 vssd1 vccd1 vccd1 net742 sky130_fd_sc_hd__clkbuf_4
Xfanout753 net754 vssd1 vssd1 vccd1 vccd1 net753 sky130_fd_sc_hd__buf_2
Xfanout764 net765 vssd1 vssd1 vccd1 vccd1 net764 sky130_fd_sc_hd__clkbuf_4
Xfanout775 net777 vssd1 vssd1 vccd1 vccd1 net775 sky130_fd_sc_hd__buf_4
Xfanout786 net789 vssd1 vssd1 vccd1 vccd1 net786 sky130_fd_sc_hd__clkbuf_4
X_15103__1483 vssd1 vssd1 vccd1 vccd1 _15103__1483/HI net1483 sky130_fd_sc_hd__conb_1
X_09859_ _05730_ net319 _05800_ _05757_ vssd1 vssd1 vccd1 vccd1 _05801_ sky130_fd_sc_hd__or4b_1
Xfanout797 net798 vssd1 vssd1 vccd1 vccd1 net797 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout750_X net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07175__C1 net1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11365__D net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08062__S1 net1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout848_X net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_161_3679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12870_ net1293 vssd1 vssd1 vccd1 vccd1 _00634_ sky130_fd_sc_hd__inv_2
X_11821_ net648 _06651_ net455 net323 net1775 vssd1 vssd1 vccd1 vccd1 _01718_ sky130_fd_sc_hd__a32o_1
XFILLER_0_157_208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_843 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07478__B1 net1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11274__A1 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14540_ clknet_leaf_22_wb_clk_i _02304_ _00905_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[894\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11381__C net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11752_ _06576_ net458 net332 net2304 vssd1 vssd1 vccd1 vccd1 _01785_ sky130_fd_sc_hd__a22o_1
XFILLER_0_68_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11813__A3 net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10703_ net523 _06339_ _06340_ net528 net1633 vssd1 vssd1 vccd1 vccd1 _02461_ sky130_fd_sc_hd__a32o_1
XFILLER_0_166_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14471_ clknet_leaf_110_wb_clk_i _02235_ _00836_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[825\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10846__X _06446_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11683_ _06725_ net386 net341 net2066 vssd1 vssd1 vccd1 vccd1 _01851_ sky130_fd_sc_hd__a22o_1
XANTENNA__12774__A net1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input91_A wbs_adr_i[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13422_ net1427 vssd1 vssd1 vccd1 vccd1 _01186_ sky130_fd_sc_hd__inv_2
X_10634_ team_03_WB.instance_to_wrap.core.decoder.inst\[27\] net1650 net847 vssd1
+ vssd1 vccd1 vccd1 _02494_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_820 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08427__C1 net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11026__B2 net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13353_ net1325 vssd1 vssd1 vccd1 vccd1 _01117_ sky130_fd_sc_hd__inv_2
XFILLER_0_10_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_423 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10565_ net1595 net533 net600 _05875_ vssd1 vssd1 vccd1 vccd1 _02558_ sky130_fd_sc_hd__a22o_1
XFILLER_0_107_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12304_ net1411 vssd1 vssd1 vccd1 vccd1 _00068_ sky130_fd_sc_hd__inv_2
XFILLER_0_134_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07650__B1 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13284_ net1345 vssd1 vssd1 vccd1 vccd1 _01048_ sky130_fd_sc_hd__inv_2
XFILLER_0_133_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10496_ net104 net1030 net907 net1654 vssd1 vssd1 vccd1 vccd1 _02613_ sky130_fd_sc_hd__a22o_1
XFILLER_0_121_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15023_ clknet_leaf_84_wb_clk_i _02743_ _01388_ vssd1 vssd1 vccd1 vccd1 net179 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11131__C_N net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12235_ net1568 vssd1 vssd1 vccd1 vccd1 _01422_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__10537__B1 net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12166_ net1543 vssd1 vssd1 vccd1 vccd1 _02387_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__11329__S net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11117_ _06632_ net2549 net418 vssd1 vssd1 vccd1 vccd1 _02243_ sky130_fd_sc_hd__mux2_1
X_12097_ _06794_ net464 net441 net1893 vssd1 vssd1 vccd1 vccd1 _01450_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_30_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11048_ net2585 net423 _06601_ net516 vssd1 vssd1 vccd1 vccd1 _02281_ sky130_fd_sc_hd__a22o_1
XANTENNA__07705__A1 net1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput8 DAT_I[15] vssd1 vssd1 vccd1 vccd1 net8 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09170__A3 _04922_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14937__Q team_03_WB.instance_to_wrap.CPU_DAT_O\[24\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11572__B net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14807_ clknet_leaf_104_wb_clk_i net1819 _01172_ vssd1 vssd1 vccd1 vccd1 net136 sky130_fd_sc_hd__dfrtp_1
X_12999_ net1370 vssd1 vssd1 vccd1 vccd1 _00763_ sky130_fd_sc_hd__inv_2
XFILLER_0_98_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14738_ clknet_leaf_32_wb_clk_i _02502_ _01103_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11291__C net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08666__C1 team_03_WB.instance_to_wrap.core.decoder.inst\[17\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11999__S net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14669_ clknet_leaf_189_wb_clk_i _02433_ _01034_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1023\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_129_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07210_ _03146_ _03151_ net821 vssd1 vssd1 vccd1 vccd1 _03152_ sky130_fd_sc_hd__mux2_1
X_08190_ net1061 _04129_ _04130_ vssd1 vssd1 vccd1 vccd1 _04132_ sky130_fd_sc_hd__or3_1
XANTENNA__08418__C1 net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_336 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_907 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11568__A2 net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07141_ net1197 net885 team_03_WB.instance_to_wrap.core.register_file.registers_state\[0\]
+ vssd1 vssd1 vccd1 vccd1 _03083_ sky130_fd_sc_hd__a21o_1
XANTENNA__08969__B1 net1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09091__C1 net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07072_ net815 _03012_ _03013_ vssd1 vssd1 vccd1 vccd1 _03014_ sky130_fd_sc_hd__and3_1
XFILLER_0_124_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_144_Left_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_2287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10528__B1 net1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10932__A net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08197__A1 net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_1840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07974_ net1111 team_03_WB.instance_to_wrap.core.register_file.registers_state\[368\]
+ net901 _03915_ net1135 vssd1 vssd1 vccd1 vccd1 _03916_ sky130_fd_sc_hd__o311a_1
XTAP_TAPCELL_ROW_143_3310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_3321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09932__S net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09713_ _05551_ _05654_ _05653_ _05652_ vssd1 vssd1 vccd1 vccd1 _05655_ sky130_fd_sc_hd__o211a_1
X_06925_ net1106 team_03_WB.instance_to_wrap.core.register_file.registers_state\[452\]
+ vssd1 vssd1 vccd1 vccd1 _02867_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout376_A _06812_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09644_ _04269_ _04326_ _04448_ _04386_ net553 net563 vssd1 vssd1 vccd1 vccd1 _05586_
+ sky130_fd_sc_hd__mux4_2
XANTENNA__09161__A3 _04532_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07960__B _03901_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06856_ net1383 vssd1 vssd1 vccd1 vccd1 _00011_ sky130_fd_sc_hd__inv_2
XFILLER_0_97_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_153_Left_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09575_ net581 _05504_ _05505_ _05516_ vssd1 vssd1 vccd1 vccd1 _05517_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_96_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout543_A _03106_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_42_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08526_ net859 _04464_ _04467_ vssd1 vssd1 vccd1 vccd1 _04468_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_72_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11256__A1 net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_731 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08657__C1 net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_775 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08457_ net1062 _04397_ _04398_ net1210 vssd1 vssd1 vccd1 vccd1 _04399_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout710_A net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout331_X net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_740 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout808_A net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1073_X net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07408_ net717 _03349_ vssd1 vssd1 vccd1 vccd1 _03350_ sky130_fd_sc_hd__or2_1
XANTENNA__07880__B1 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08283__S net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08388_ net947 _04328_ _04329_ vssd1 vssd1 vccd1 vccd1 _04330_ sky130_fd_sc_hd__o21a_1
XFILLER_0_46_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07339_ net1083 net888 team_03_WB.instance_to_wrap.core.register_file.registers_state\[28\]
+ vssd1 vssd1 vccd1 vccd1 _03281_ sky130_fd_sc_hd__o21a_1
XANTENNA__09621__A1 net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1240_X net1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_162_Left_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11003__A net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1338_X net1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_2733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10350_ _06184_ _06183_ net284 vssd1 vssd1 vccd1 vccd1 _06185_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_115_2744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout798_X net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_167_3800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09009_ net871 _04949_ _04950_ vssd1 vssd1 vccd1 vccd1 _04951_ sky130_fd_sc_hd__or3b_1
XFILLER_0_42_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_167_3811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10281_ _05975_ _06111_ _06120_ _06122_ vssd1 vssd1 vccd1 vccd1 _06123_ sky130_fd_sc_hd__a31o_1
XANTENNA__10519__B1 net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12020_ net623 _06581_ net457 net359 net2135 vssd1 vssd1 vccd1 vccd1 _01525_ sky130_fd_sc_hd__a32o_1
XFILLER_0_104_1128 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout965_X net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_163_3719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07935__A1 net1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11731__A2 _06505_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout550 net552 vssd1 vssd1 vccd1 vccd1 net550 sky130_fd_sc_hd__buf_2
XANTENNA_clkbuf_leaf_81_wb_clk_i_A clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout561 net562 vssd1 vssd1 vccd1 vccd1 net561 sky130_fd_sc_hd__buf_2
Xfanout572 _03024_ vssd1 vssd1 vccd1 vccd1 net572 sky130_fd_sc_hd__clkbuf_4
Xfanout583 _02892_ vssd1 vssd1 vccd1 vccd1 net583 sky130_fd_sc_hd__clkbuf_4
X_13971_ clknet_leaf_103_wb_clk_i _01735_ _00336_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[325\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09688__A1 net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout594 net595 vssd1 vssd1 vccd1 vccd1 net594 sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_171_Left_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07699__A0 _03638_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12922_ net1373 vssd1 vssd1 vccd1 vccd1 _00686_ sky130_fd_sc_hd__inv_2
XANTENNA__09152__A3 _04444_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12853_ net1272 vssd1 vssd1 vccd1 vccd1 _00617_ sky130_fd_sc_hd__inv_2
XFILLER_0_69_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11804_ net2527 net264 net329 vssd1 vssd1 vccd1 vccd1 _01734_ sky130_fd_sc_hd__mux2_1
X_12784_ net1411 vssd1 vssd1 vccd1 vccd1 _00548_ sky130_fd_sc_hd__inv_2
XFILLER_0_138_230 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14523_ clknet_leaf_124_wb_clk_i _02287_ _00888_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[877\]
+ sky130_fd_sc_hd__dfrtp_1
X_11735_ net1888 net295 net337 vssd1 vssd1 vccd1 vccd1 _01801_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_548 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07598__A net1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input94_X net94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14454_ clknet_leaf_152_wb_clk_i _02218_ _00819_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[808\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_436 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07871__B1 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11666_ net2000 _06628_ net344 vssd1 vssd1 vccd1 vccd1 _01867_ sky130_fd_sc_hd__mux2_1
X_13405_ net1407 vssd1 vssd1 vccd1 vccd1 _01169_ sky130_fd_sc_hd__inv_2
X_10617_ net1710 team_03_WB.instance_to_wrap.CPU_DAT_O\[12\] net842 vssd1 vssd1 vccd1
+ vccd1 _02511_ sky130_fd_sc_hd__mux2_1
X_14385_ clknet_leaf_139_wb_clk_i _02149_ _00750_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[739\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10758__B1 net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11597_ net270 net2513 net447 vssd1 vssd1 vccd1 vccd1 _01932_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13336_ net1333 vssd1 vssd1 vccd1 vccd1 _01100_ sky130_fd_sc_hd__inv_2
X_10548_ _06287_ _06290_ _06291_ team_03_WB.instance_to_wrap.BUSY_O vssd1 vssd1 vccd1
+ vccd1 _02567_ sky130_fd_sc_hd__o22a_1
XFILLER_0_150_940 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13267_ net1265 vssd1 vssd1 vccd1 vccd1 _01031_ sky130_fd_sc_hd__inv_2
X_10479_ net1634 net1028 net906 net1633 vssd1 vssd1 vccd1 vccd1 _02630_ sky130_fd_sc_hd__a22o_1
X_15006_ clknet_leaf_7_wb_clk_i net54 _01371_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[25\]
+ sky130_fd_sc_hd__dfrtp_4
X_12218_ net1557 vssd1 vssd1 vccd1 vccd1 _01439_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11567__B net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13198_ net1303 vssd1 vssd1 vccd1 vccd1 _00962_ sky130_fd_sc_hd__inv_2
XANTENNA__11722__A2 net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10671__C_N _05563_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10902__D net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12149_ net1573 vssd1 vssd1 vccd1 vccd1 _02404_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__09605__X _05547_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09143__A3 net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07690_ _03630_ _03631_ net1162 vssd1 vssd1 vccd1 vccd1 _03632_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_155_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07272__S net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11238__A1 net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09360_ _05278_ _05281_ _05301_ vssd1 vssd1 vccd1 vccd1 _05302_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_47_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08639__C1 net1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08892__A net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_824 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09300__B1 net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08311_ net1242 team_03_WB.instance_to_wrap.core.register_file.registers_state\[728\]
+ net985 team_03_WB.instance_to_wrap.core.register_file.registers_state\[760\] net939
+ vssd1 vssd1 vccd1 vccd1 _04253_ sky130_fd_sc_hd__o221a_1
XFILLER_0_157_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09291_ _05227_ _05232_ vssd1 vssd1 vccd1 vccd1 _05233_ sky130_fd_sc_hd__nand2_1
XANTENNA__07311__C1 net1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08654__A2 net1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_126_wb_clk_i_A clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_75_879 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_157_594 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08242_ net1226 team_03_WB.instance_to_wrap.core.register_file.registers_state\[82\]
+ net950 team_03_WB.instance_to_wrap.core.register_file.registers_state\[114\] net916
+ vssd1 vssd1 vccd1 vccd1 _04184_ sky130_fd_sc_hd__o221a_1
XANTENNA__07862__B1 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_656 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_59_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_59_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_16_935 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_144_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10138__S net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08173_ net1230 team_03_WB.instance_to_wrap.core.register_file.registers_state\[852\]
+ net958 team_03_WB.instance_to_wrap.core.register_file.registers_state\[884\] net1217
+ vssd1 vssd1 vccd1 vccd1 _04115_ sky130_fd_sc_hd__o221a_1
XANTENNA__09064__C1 net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_2327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_166_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07124_ net614 _03065_ vssd1 vssd1 vccd1 vccd1 _03066_ sky130_fd_sc_hd__or2_1
XANTENNA__07614__B1 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_3077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_132_3088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07055_ net1095 team_03_WB.instance_to_wrap.core.register_file.registers_state\[962\]
+ net796 team_03_WB.instance_to_wrap.core.register_file.registers_state\[994\] net1131
+ vssd1 vssd1 vccd1 vccd1 _02997_ sky130_fd_sc_hd__a221o_1
XANTENNA__07090__A1 net1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_815 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput120 net120 vssd1 vssd1 vccd1 vccd1 ADR_O[25] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_113_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput131 net131 vssd1 vssd1 vccd1 vccd1 ADR_O[6] sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout1033_A net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_9_wb_clk_i_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xoutput142 net142 vssd1 vssd1 vccd1 vccd1 DAT_O[15] sky130_fd_sc_hd__buf_2
XFILLER_0_88_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput153 net153 vssd1 vssd1 vccd1 vccd1 DAT_O[25] sky130_fd_sc_hd__buf_2
XANTENNA__09228__A _04532_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_2630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11477__B net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput164 net164 vssd1 vssd1 vccd1 vccd1 DAT_O[6] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_110_2641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput175 net175 vssd1 vssd1 vccd1 vccd1 gpio_oeb[10] sky130_fd_sc_hd__clkbuf_4
XANTENNA__07378__C1 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout493_A net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11174__B1 net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput186 net186 vssd1 vssd1 vccd1 vccd1 gpio_oeb[21] sky130_fd_sc_hd__buf_2
Xoutput197 net197 vssd1 vssd1 vccd1 vccd1 gpio_oeb[32] sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout1200_A net1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11196__C net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08590__A1 net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07957_ net1116 _03897_ _03898_ _03894_ vssd1 vssd1 vccd1 vccd1 _03899_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout660_A _05950_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout281_X net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout758_A net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout379_X net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06908_ net1096 net896 vssd1 vssd1 vccd1 vccd1 _02850_ sky130_fd_sc_hd__nor2_1
X_07888_ net1186 team_03_WB.instance_to_wrap.core.register_file.registers_state\[111\]
+ net877 _03829_ vssd1 vssd1 vccd1 vccd1 _03830_ sky130_fd_sc_hd__a31o_1
XANTENNA__08342__A1 net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_165_wb_clk_i_A clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09627_ net575 _05568_ _05566_ vssd1 vssd1 vccd1 vccd1 _05569_ sky130_fd_sc_hd__o21ai_2
X_06839_ team_03_WB.instance_to_wrap.core.decoder.inst\[31\] vssd1 vssd1 vccd1 vccd1
+ _02782_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_108_2592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1190_X net1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout925_A net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09558_ _05479_ _05499_ vssd1 vssd1 vccd1 vccd1 _05500_ sky130_fd_sc_hd__nor2_1
XFILLER_0_38_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08509_ net934 _04449_ _04450_ net854 vssd1 vssd1 vccd1 vccd1 _04451_ sky130_fd_sc_hd__o211a_1
XFILLER_0_77_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09489_ _05332_ _05430_ _05324_ vssd1 vssd1 vccd1 vccd1 _05431_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout713_X net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11520_ _06633_ net2572 net391 vssd1 vssd1 vccd1 vccd1 _01986_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_156_3578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_22_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_907 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07849__C net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08307__A net1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11451_ net2341 net392 _06764_ net497 vssd1 vssd1 vccd1 vccd1 _02041_ sky130_fd_sc_hd__a22o_1
XFILLER_0_34_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_163_586 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10402_ net284 _06142_ _06224_ net680 vssd1 vssd1 vccd1 vccd1 _06228_ sky130_fd_sc_hd__o31a_1
XFILLER_0_150_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10204__A2 _05950_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14170_ clknet_leaf_147_wb_clk_i _01934_ _00535_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[524\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_33_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11382_ net516 net642 _06743_ net403 net2040 vssd1 vssd1 vccd1 vccd1 _02089_ sky130_fd_sc_hd__a32o_1
X_13121_ net1260 vssd1 vssd1 vccd1 vccd1 _00885_ sky130_fd_sc_hd__inv_2
XANTENNA__07081__A1 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10333_ _06118_ _06170_ vssd1 vssd1 vccd1 vccd1 _06171_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07357__S net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09138__A net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13052_ net1413 vssd1 vssd1 vccd1 vccd1 _00816_ sky130_fd_sc_hd__inv_2
XANTENNA_input54_A gpio_in[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11387__B net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10264_ _06092_ _06102_ _06104_ _06105_ vssd1 vssd1 vccd1 vccd1 _06106_ sky130_fd_sc_hd__a31o_1
X_12003_ net268 net2543 net445 vssd1 vssd1 vccd1 vccd1 _01541_ sky130_fd_sc_hd__mux2_1
XANTENNA__11704__A2 net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1301 net1302 vssd1 vssd1 vccd1 vccd1 net1301 sky130_fd_sc_hd__clkbuf_4
X_10195_ _06035_ _06036_ vssd1 vssd1 vccd1 vccd1 _06037_ sky130_fd_sc_hd__nor2_1
Xfanout1312 net1330 vssd1 vssd1 vccd1 vccd1 net1312 sky130_fd_sc_hd__clkbuf_4
Xfanout1323 net1324 vssd1 vssd1 vccd1 vccd1 net1323 sky130_fd_sc_hd__buf_2
Xfanout1334 net1335 vssd1 vssd1 vccd1 vccd1 net1334 sky130_fd_sc_hd__buf_2
Xfanout1345 net1346 vssd1 vssd1 vccd1 vccd1 net1345 sky130_fd_sc_hd__buf_4
Xfanout1356 net1357 vssd1 vssd1 vccd1 vccd1 net1356 sky130_fd_sc_hd__buf_4
Xfanout1367 net1370 vssd1 vssd1 vccd1 vccd1 net1367 sky130_fd_sc_hd__buf_2
Xfanout1378 net1381 vssd1 vssd1 vccd1 vccd1 net1378 sky130_fd_sc_hd__buf_2
Xfanout380 net387 vssd1 vssd1 vccd1 vccd1 net380 sky130_fd_sc_hd__buf_2
Xfanout1389 net1393 vssd1 vssd1 vccd1 vccd1 net1389 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11607__S net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout391 _06778_ vssd1 vssd1 vccd1 vccd1 net391 sky130_fd_sc_hd__buf_4
X_13954_ clknet_leaf_174_wb_clk_i _01718_ _00319_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[308\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09530__B1 net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12905_ net1257 vssd1 vssd1 vccd1 vccd1 _00669_ sky130_fd_sc_hd__inv_2
X_13885_ clknet_leaf_24_wb_clk_i _01649_ _00250_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[239\]
+ sky130_fd_sc_hd__dfrtp_1
X_12836_ net1382 vssd1 vssd1 vccd1 vccd1 _00600_ sky130_fd_sc_hd__inv_2
XANTENNA__08916__S net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08097__B1 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12767_ net1348 vssd1 vssd1 vccd1 vccd1 _00531_ sky130_fd_sc_hd__inv_2
XANTENNA__10979__A0 net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09833__A1 net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14506_ clknet_leaf_7_wb_clk_i _02270_ _00871_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[860\]
+ sky130_fd_sc_hd__dfrtp_1
X_11718_ net2080 net276 net335 vssd1 vssd1 vccd1 vccd1 _01818_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12698_ net1379 vssd1 vssd1 vccd1 vccd1 _00462_ sky130_fd_sc_hd__inv_2
XFILLER_0_72_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14437_ clknet_leaf_39_wb_clk_i _02201_ _00802_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[791\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput11 DAT_I[18] vssd1 vssd1 vccd1 vccd1 net11 sky130_fd_sc_hd__clkbuf_1
X_11649_ net2756 _06615_ net342 vssd1 vssd1 vccd1 vccd1 _01884_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09046__C1 net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput22 DAT_I[28] vssd1 vssd1 vccd1 vccd1 net22 sky130_fd_sc_hd__buf_1
XFILLER_0_114_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_140_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput33 DAT_I[9] vssd1 vssd1 vccd1 vccd1 net33 sky130_fd_sc_hd__clkbuf_1
Xinput44 gpio_in[19] vssd1 vssd1 vccd1 vccd1 net44 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_141_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput55 gpio_in[30] vssd1 vssd1 vccd1 vccd1 net55 sky130_fd_sc_hd__clkbuf_1
X_14368_ clknet_leaf_191_wb_clk_i _02132_ _00733_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[722\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput66 wb_rst_i vssd1 vssd1 vccd1 vccd1 net66 sky130_fd_sc_hd__clkbuf_1
Xinput77 wbs_adr_i[19] vssd1 vssd1 vccd1 vccd1 net77 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold806 team_03_WB.instance_to_wrap.core.register_file.registers_state\[353\] vssd1
+ vssd1 vccd1 vccd1 net2299 sky130_fd_sc_hd__dlygate4sd3_1
Xhold817 team_03_WB.instance_to_wrap.core.register_file.registers_state\[26\] vssd1
+ vssd1 vccd1 vccd1 net2310 sky130_fd_sc_hd__dlygate4sd3_1
Xinput88 wbs_adr_i[29] vssd1 vssd1 vccd1 vccd1 net88 sky130_fd_sc_hd__buf_1
XANTENNA__09698__A1_N _02804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13319_ net1318 vssd1 vssd1 vccd1 vccd1 _01083_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold828 team_03_WB.instance_to_wrap.core.register_file.registers_state\[43\] vssd1
+ vssd1 vccd1 vccd1 net2321 sky130_fd_sc_hd__dlygate4sd3_1
Xhold839 team_03_WB.instance_to_wrap.core.register_file.registers_state\[627\] vssd1
+ vssd1 vccd1 vccd1 net2332 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput99 wbs_cyc_i vssd1 vssd1 vccd1 vccd1 net99 sky130_fd_sc_hd__clkbuf_2
X_14299_ clknet_leaf_121_wb_clk_i _02063_ _00664_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[653\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_90_2224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_2235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11297__B _06557_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_177_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_177_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_08860_ net1056 team_03_WB.instance_to_wrap.core.register_file.registers_state\[832\]
+ net1010 team_03_WB.instance_to_wrap.core.register_file.registers_state\[864\] net1216
+ vssd1 vssd1 vccd1 vccd1 _04802_ sky130_fd_sc_hd__a221o_1
XANTENNA__07375__A2 net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08572__A1 net1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07811_ net1131 _03751_ net1164 vssd1 vssd1 vccd1 vccd1 _03753_ sky130_fd_sc_hd__o21ai_1
Xclkbuf_leaf_106_wb_clk_i clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_106_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_08791_ net1050 team_03_WB.instance_to_wrap.core.register_file.registers_state\[674\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[642\] net1002 net943
+ vssd1 vssd1 vccd1 vccd1 _04733_ sky130_fd_sc_hd__o221a_1
XFILLER_0_74_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11517__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07742_ net1098 _02795_ net897 vssd1 vssd1 vccd1 vccd1 _03684_ sky130_fd_sc_hd__or3_1
XANTENNA__11459__B2 net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_2175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_2186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08324__B2 net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07673_ net1178 team_03_WB.instance_to_wrap.core.register_file.registers_state\[350\]
+ net771 team_03_WB.instance_to_wrap.core.register_file.registers_state\[382\] net1126
+ vssd1 vssd1 vccd1 vccd1 _03615_ sky130_fd_sc_hd__o221a_1
XFILLER_0_149_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08875__A2 _04770_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09412_ _05350_ _05353_ net564 vssd1 vssd1 vccd1 vccd1 _05354_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08088__B1 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09343_ _05283_ _05284_ vssd1 vssd1 vccd1 vccd1 _05285_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_158_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_158_Right_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout339_A _06806_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_62_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09274_ _04953_ _05215_ vssd1 vssd1 vccd1 vccd1 _05216_ sky130_fd_sc_hd__nor2_1
XFILLER_0_118_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07835__B1 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_134_3117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07669__C net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_145_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_134_3128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_326 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08225_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[817\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[785\]
+ net962 vssd1 vssd1 vccd1 vccd1 _04167_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12872__A net1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1150_A net1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout506_A net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1248_A net1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09588__B1 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08156_ net1230 team_03_WB.instance_to_wrap.core.register_file.registers_state\[340\]
+ net961 team_03_WB.instance_to_wrap.core.register_file.registers_state\[372\] net1071
+ vssd1 vssd1 vccd1 vccd1 _04098_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_151_3475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10198__A1 team_03_WB.instance_to_wrap.core.pc.current_pc\[4\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11488__A net1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07107_ _03046_ _03048_ net1118 _03044_ vssd1 vssd1 vccd1 vccd1 _03049_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_160_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08087_ net722 _03999_ _04007_ _04028_ vssd1 vssd1 vccd1 vccd1 _04029_ sky130_fd_sc_hd__o31a_2
XANTENNA_fanout1036_X net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07038_ net1099 team_03_WB.instance_to_wrap.core.register_file.registers_state\[195\]
+ net801 team_03_WB.instance_to_wrap.core.register_file.registers_state\[227\] net731
+ vssd1 vssd1 vccd1 vccd1 _02980_ sky130_fd_sc_hd__a221o_1
XFILLER_0_30_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11147__B1 net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout496_X net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08012__B1 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1203_X net1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input1_X net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout663_X net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08989_ _04927_ _04930_ net867 vssd1 vssd1 vccd1 vccd1 _04931_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07771__C1 net1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13208__A net1380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08315__A1 net1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_2990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09899__Y _05841_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10951_ team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[4\] net308 net689 vssd1
+ vssd1 vccd1 vccd1 _06534_ sky130_fd_sc_hd__a21o_1
XFILLER_0_98_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout830_X net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08410__S1 net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout928_X net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_158_3618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_158_3629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13670_ clknet_leaf_75_wb_clk_i _01434_ _00035_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_10882_ net692 _06475_ _06476_ _06474_ vssd1 vssd1 vccd1 vccd1 _06478_ sky130_fd_sc_hd__a31o_4
XTAP_TAPCELL_ROW_123_2898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12621_ net1331 vssd1 vssd1 vccd1 vccd1 _00385_ sky130_fd_sc_hd__inv_2
XFILLER_0_38_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09815__A1 _02954_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_125_Right_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07826__B1 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12552_ net1299 vssd1 vssd1 vccd1 vccd1 _00316_ sky130_fd_sc_hd__inv_2
XFILLER_0_65_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11503_ _06479_ net2546 net388 vssd1 vssd1 vccd1 vccd1 _02003_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10830__C1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12483_ net1371 vssd1 vssd1 vccd1 vccd1 _00247_ sky130_fd_sc_hd__inv_2
X_14222_ clknet_leaf_131_wb_clk_i _01986_ _00587_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[576\]
+ sky130_fd_sc_hd__dfrtp_1
X_11434_ _06557_ net2352 net398 vssd1 vssd1 vccd1 vccd1 _02050_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11386__B1 net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14153_ clknet_leaf_75_wb_clk_i _01917_ _00518_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[507\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11365_ net1250 net839 net299 net669 vssd1 vssd1 vccd1 vccd1 _06735_ sky130_fd_sc_hd__and4_1
Xclkbuf_leaf_4_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_4_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_81_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13104_ net1412 vssd1 vssd1 vccd1 vccd1 _00868_ sky130_fd_sc_hd__inv_2
X_10316_ net282 _06128_ _06156_ vssd1 vssd1 vccd1 vccd1 _06157_ sky130_fd_sc_hd__and3_1
X_14084_ clknet_leaf_36_wb_clk_i _01848_ _00449_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[438\]
+ sky130_fd_sc_hd__dfrtp_1
X_11296_ net509 net636 _06715_ net410 net2181 vssd1 vssd1 vccd1 vccd1 _02147_ sky130_fd_sc_hd__a32o_1
XFILLER_0_120_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13035_ net1288 vssd1 vssd1 vccd1 vccd1 _00799_ sky130_fd_sc_hd__inv_2
X_10247_ _05986_ _05991_ _06086_ _05988_ _05983_ vssd1 vssd1 vccd1 vccd1 _06089_ sky130_fd_sc_hd__o311ai_4
XFILLER_0_119_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08554__A1 net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1120 net1122 vssd1 vssd1 vccd1 vccd1 net1120 sky130_fd_sc_hd__buf_6
XANTENNA__09751__B1 net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1131 net1132 vssd1 vssd1 vccd1 vccd1 net1131 sky130_fd_sc_hd__buf_4
Xfanout1142 _02765_ vssd1 vssd1 vccd1 vccd1 net1142 sky130_fd_sc_hd__clkbuf_4
X_10178_ _03242_ _06018_ _06019_ vssd1 vssd1 vccd1 vccd1 _06020_ sky130_fd_sc_hd__and3_1
XANTENNA__10361__A1 net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1153 net1159 vssd1 vssd1 vccd1 vccd1 net1153 sky130_fd_sc_hd__buf_2
XFILLER_0_28_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1164 net1166 vssd1 vssd1 vccd1 vccd1 net1164 sky130_fd_sc_hd__buf_4
Xfanout1175 net1179 vssd1 vssd1 vccd1 vccd1 net1175 sky130_fd_sc_hd__clkbuf_4
Xfanout1186 net1188 vssd1 vssd1 vccd1 vccd1 net1186 sky130_fd_sc_hd__buf_2
XANTENNA__09729__S1 net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1197 net1198 vssd1 vssd1 vccd1 vccd1 net1197 sky130_fd_sc_hd__clkbuf_4
X_14986_ clknet_leaf_66_wb_clk_i net65 _01351_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12102__A2 net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13937_ clknet_leaf_143_wb_clk_i _01701_ _00302_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[291\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_407 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13868_ clknet_leaf_19_wb_clk_i _01632_ _00233_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[222\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_83_2072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_818 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_2083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12819_ net1271 vssd1 vssd1 vccd1 vccd1 _00583_ sky130_fd_sc_hd__inv_2
XFILLER_0_57_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13799_ clknet_leaf_108_wb_clk_i _01563_ _00164_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[153\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07817__A0 _03756_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_451 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07122__Y _03064_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09282__A2 _05146_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10196__B _05950_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_873 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11800__S net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08010_ net1125 _03950_ _03951_ net1115 _03949_ vssd1 vssd1 vccd1 vccd1 _03952_ sky130_fd_sc_hd__a311o_1
XFILLER_0_25_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10924__B net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold603 team_03_WB.instance_to_wrap.core.register_file.registers_state\[284\] vssd1
+ vssd1 vccd1 vccd1 net2096 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07045__A1 net1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_770 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold614 team_03_WB.instance_to_wrap.core.register_file.registers_state\[405\] vssd1
+ vssd1 vccd1 vccd1 net2107 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold625 team_03_WB.instance_to_wrap.core.register_file.registers_state\[270\] vssd1
+ vssd1 vccd1 vccd1 net2118 sky130_fd_sc_hd__dlygate4sd3_1
Xhold636 team_03_WB.instance_to_wrap.core.register_file.registers_state\[345\] vssd1
+ vssd1 vccd1 vccd1 net2129 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08793__A1 net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold647 team_03_WB.instance_to_wrap.core.register_file.registers_state\[249\] vssd1
+ vssd1 vccd1 vccd1 net2140 sky130_fd_sc_hd__dlygate4sd3_1
Xhold658 team_03_WB.instance_to_wrap.core.register_file.registers_state\[634\] vssd1
+ vssd1 vccd1 vccd1 net2151 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09961_ _03678_ net661 vssd1 vssd1 vccd1 vccd1 _05885_ sky130_fd_sc_hd__nor2_2
XFILLER_0_0_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold669 team_03_WB.instance_to_wrap.core.register_file.registers_state\[239\] vssd1
+ vssd1 vccd1 vccd1 net2162 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08912_ net1208 _04850_ _04853_ vssd1 vssd1 vccd1 vccd1 _04854_ sky130_fd_sc_hd__or3_1
XFILLER_0_110_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09892_ _05182_ _05502_ _05503_ net594 vssd1 vssd1 vccd1 vccd1 _05834_ sky130_fd_sc_hd__a211o_1
XANTENNA__10888__C1 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08843_ net1056 team_03_WB.instance_to_wrap.core.register_file.registers_state\[192\]
+ net1009 team_03_WB.instance_to_wrap.core.register_file.registers_state\[224\] net930
+ vssd1 vssd1 vccd1 vccd1 _04785_ sky130_fd_sc_hd__a221o_1
XANTENNA__07899__A3 net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout289_A net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10151__S net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08774_ net1240 team_03_WB.instance_to_wrap.core.register_file.registers_state\[130\]
+ net977 team_03_WB.instance_to_wrap.core.register_file.registers_state\[162\] net943
+ vssd1 vssd1 vccd1 vccd1 _04716_ sky130_fd_sc_hd__o221a_1
XANTENNA__09940__S net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07725_ net1097 team_03_WB.instance_to_wrap.core.register_file.registers_state\[653\]
+ net732 _03666_ vssd1 vssd1 vccd1 vccd1 _03667_ sky130_fd_sc_hd__a211o_1
XANTENNA__10939__X _06524_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_2540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout456_A net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07505__C1 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1198_A net1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07656_ net1119 _03597_ net1139 vssd1 vssd1 vccd1 vccd1 _03598_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_95_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_74_wb_clk_i clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_74_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_165_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_101_2448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07587_ _03526_ _03528_ net610 vssd1 vssd1 vccd1 vccd1 _03529_ sky130_fd_sc_hd__mux2_2
XANTENNA_fanout623_A net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_2459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1365_A net1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09326_ _05265_ _05267_ _05253_ vssd1 vssd1 vccd1 vccd1 _05268_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_48_676 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_153_3515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_153_3526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07284__A1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[9\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09895__B _04323_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09257_ _04072_ _05147_ net608 vssd1 vssd1 vccd1 vccd1 _05199_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_106_715 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10674__X _06316_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08481__B1 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout411_X net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1153_X net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout509_X net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_170_3862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08208_ _04120_ net354 net548 vssd1 vssd1 vccd1 vccd1 _04150_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_170_3873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_331 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09188_ _05128_ _05129_ vssd1 vssd1 vccd1 vccd1 _05130_ sky130_fd_sc_hd__nor2_1
XANTENNA__08144__X _04086_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout992_A net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11368__B1 net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_578 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08139_ net1081 net1015 vssd1 vssd1 vccd1 vccd1 _04081_ sky130_fd_sc_hd__nor2_1
XFILLER_0_31_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_79_1996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10040__B1 net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11011__A net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11150_ net704 _06468_ net696 vssd1 vssd1 vccd1 vccd1 _06652_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout780_X net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10591__A1 _06293_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout878_X net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10101_ _05921_ _05922_ _05941_ _05944_ _05920_ vssd1 vssd1 vccd1 vccd1 _05945_ sky130_fd_sc_hd__a221o_4
XFILLER_0_101_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11081_ _06618_ net2493 net417 vssd1 vssd1 vccd1 vccd1 _02265_ sky130_fd_sc_hd__mux2_1
XANTENNA__07339__A2 net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10032_ net26 net1036 net909 net2228 vssd1 vssd1 vccd1 vccd1 _02699_ sky130_fd_sc_hd__o22a_1
XANTENNA__11540__B1 net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07744__C1 net1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14840_ clknet_leaf_87_wb_clk_i _02604_ _01205_ vssd1 vssd1 vccd1 vccd1 net114 sky130_fd_sc_hd__dfrtp_1
XANTENNA__09135__B _05076_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14771_ clknet_leaf_104_wb_clk_i _02535_ _01136_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_I\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input17_A DAT_I[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11983_ net301 net2613 net446 vssd1 vssd1 vccd1 vccd1 _01561_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_919 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08839__A2 net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_932 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08395__S0 net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13722_ clknet_leaf_141_wb_clk_i _01486_ _00087_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[76\]
+ sky130_fd_sc_hd__dfrtp_1
X_10934_ net688 _05730_ _06399_ vssd1 vssd1 vccd1 vccd1 _06520_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_14_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13653_ clknet_leaf_127_wb_clk_i _01417_ _00018_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_156_626 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10865_ net656 net704 _06463_ vssd1 vssd1 vccd1 vccd1 _06464_ sky130_fd_sc_hd__and3_1
XFILLER_0_39_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12604_ net1414 vssd1 vssd1 vccd1 vccd1 _00368_ sky130_fd_sc_hd__inv_2
XFILLER_0_27_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13584_ net1345 vssd1 vssd1 vccd1 vccd1 _01348_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10796_ net281 net2618 net518 vssd1 vssd1 vccd1 vccd1 _02337_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07275__A1 net1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12535_ net1385 vssd1 vssd1 vccd1 vccd1 _00299_ sky130_fd_sc_hd__inv_2
XFILLER_0_81_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12466_ net1395 vssd1 vssd1 vccd1 vccd1 _00230_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10744__B net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14205_ clknet_leaf_26_wb_clk_i _01969_ _00570_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[559\]
+ sky130_fd_sc_hd__dfrtp_1
X_11417_ _06491_ net2435 net398 vssd1 vssd1 vccd1 vccd1 _02064_ sky130_fd_sc_hd__mux2_1
XANTENNA__10236__S net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12397_ net1331 vssd1 vssd1 vccd1 vccd1 _00161_ sky130_fd_sc_hd__inv_2
X_14136_ clknet_leaf_185_wb_clk_i _01900_ _00501_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[490\]
+ sky130_fd_sc_hd__dfrtp_1
X_11348_ net512 net640 _06726_ net400 net1896 vssd1 vssd1 vccd1 vccd1 _02106_ sky130_fd_sc_hd__a32o_1
XFILLER_0_120_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10582__B2 _03488_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14067_ clknet_leaf_106_wb_clk_i _01831_ _00432_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[421\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10760__A _05784_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11279_ net714 net296 net830 vssd1 vssd1 vccd1 vccd1 _06707_ sky130_fd_sc_hd__and3_1
XANTENNA__08527__A1 net1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09724__B1 net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13018_ net1372 vssd1 vssd1 vccd1 vccd1 _00782_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11531__B1 net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11067__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_33 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_85_2123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12087__A1 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14969_ clknet_leaf_92_wb_clk_i _02721_ _01334_ vssd1 vssd1 vccd1 vccd1 net221 sky130_fd_sc_hd__dfrtp_1
X_07510_ net1109 team_03_WB.instance_to_wrap.core.register_file.registers_state\[455\]
+ vssd1 vssd1 vccd1 vccd1 _03452_ sky130_fd_sc_hd__and2_1
X_08490_ net1243 team_03_WB.instance_to_wrap.core.register_file.registers_state\[187\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[155\] net987 net921
+ vssd1 vssd1 vccd1 vccd1 _04432_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_18_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08376__S net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_604 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07441_ net1179 team_03_WB.instance_to_wrap.core.register_file.registers_state\[340\]
+ net764 team_03_WB.instance_to_wrap.core.register_file.registers_state\[372\] net1125
+ vssd1 vssd1 vccd1 vccd1 _03383_ sky130_fd_sc_hd__o221a_1
XFILLER_0_174_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07372_ _03312_ _03313_ net610 vssd1 vssd1 vccd1 vccd1 _03314_ sky130_fd_sc_hd__mux2_2
XFILLER_0_17_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11598__A0 net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08689__S1 net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09111_ net1222 _05050_ _05051_ vssd1 vssd1 vccd1 vccd1 _05053_ sky130_fd_sc_hd__and3_1
XANTENNA__07266__A1 net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11062__A2 net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13311__A net1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09042_ net848 _04970_ _04983_ vssd1 vssd1 vccd1 vccd1 _04984_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_72_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08405__A net1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_192_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_192_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xhold400 team_03_WB.instance_to_wrap.core.register_file.registers_state\[40\] vssd1
+ vssd1 vccd1 vccd1 net1893 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12011__A1 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold411 team_03_WB.instance_to_wrap.core.register_file.registers_state\[310\] vssd1
+ vssd1 vccd1 vccd1 net1904 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold422 team_03_WB.instance_to_wrap.core.register_file.registers_state\[802\] vssd1
+ vssd1 vccd1 vccd1 net1915 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08766__A1 net1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07569__A2 net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold433 team_03_WB.instance_to_wrap.core.register_file.registers_state\[560\] vssd1
+ vssd1 vccd1 vccd1 net1926 sky130_fd_sc_hd__dlygate4sd3_1
Xhold444 team_03_WB.instance_to_wrap.core.register_file.registers_state\[165\] vssd1
+ vssd1 vccd1 vccd1 net1937 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_121_wb_clk_i clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_121_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_57_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold455 team_03_WB.instance_to_wrap.core.register_file.registers_state\[559\] vssd1
+ vssd1 vccd1 vccd1 net1948 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11188__D net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold466 team_03_WB.instance_to_wrap.core.register_file.registers_state\[826\] vssd1
+ vssd1 vccd1 vccd1 net1959 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10573__B2 net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_3016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07974__C1 net1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold477 team_03_WB.instance_to_wrap.core.register_file.registers_state\[440\] vssd1
+ vssd1 vccd1 vccd1 net1970 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11770__B1 net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_3027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09944_ _05876_ net1753 net294 vssd1 vssd1 vccd1 vccd1 _02755_ sky130_fd_sc_hd__mux2_1
Xfanout902 net903 vssd1 vssd1 vccd1 vccd1 net902 sky130_fd_sc_hd__clkbuf_4
Xhold488 net186 vssd1 vssd1 vccd1 vccd1 net1981 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout913 net914 vssd1 vssd1 vccd1 vccd1 net913 sky130_fd_sc_hd__buf_1
XANTENNA__10670__A _05583_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold499 team_03_WB.instance_to_wrap.core.register_file.registers_state\[442\] vssd1
+ vssd1 vccd1 vccd1 net1992 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1113_A _02787_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout924 net932 vssd1 vssd1 vccd1 vccd1 net924 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_74_1893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout935 net936 vssd1 vssd1 vccd1 vccd1 net935 sky130_fd_sc_hd__clkbuf_4
Xfanout946 net948 vssd1 vssd1 vccd1 vccd1 net946 sky130_fd_sc_hd__buf_4
X_09875_ _03604_ _04820_ _05069_ _03601_ net1021 vssd1 vssd1 vccd1 vccd1 _05817_ sky130_fd_sc_hd__a32o_1
XANTENNA__08140__A net1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input9_A DAT_I[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout957 net958 vssd1 vssd1 vccd1 vccd1 net957 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_146_3363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout968 net969 vssd1 vssd1 vccd1 vccd1 net968 sky130_fd_sc_hd__clkbuf_4
Xhold1100 team_03_WB.instance_to_wrap.core.register_file.registers_state\[223\] vssd1
+ vssd1 vccd1 vccd1 net2593 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_146_3374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_hold1221_A team_03_WB.instance_to_wrap.CPU_DAT_O\[6\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout979 net981 vssd1 vssd1 vccd1 vccd1 net979 sky130_fd_sc_hd__clkbuf_4
Xhold1111 team_03_WB.instance_to_wrap.core.register_file.registers_state\[121\] vssd1
+ vssd1 vccd1 vccd1 net2604 sky130_fd_sc_hd__dlygate4sd3_1
X_08826_ net1224 _04763_ _04764_ _04767_ net1081 vssd1 vssd1 vccd1 vccd1 _04768_ sky130_fd_sc_hd__o311a_1
Xhold1122 team_03_WB.instance_to_wrap.core.register_file.registers_state\[75\] vssd1
+ vssd1 vccd1 vccd1 net2615 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1133 team_03_WB.instance_to_wrap.core.register_file.registers_state\[153\] vssd1
+ vssd1 vccd1 vccd1 net2626 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1144 team_03_WB.instance_to_wrap.core.register_file.registers_state\[733\] vssd1
+ vssd1 vccd1 vccd1 net2637 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1155 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[22\] vssd1 vssd1
+ vccd1 vccd1 net2648 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07741__A2 net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1166 team_03_WB.instance_to_wrap.core.register_file.registers_state\[831\] vssd1
+ vssd1 vccd1 vccd1 net2659 sky130_fd_sc_hd__dlygate4sd3_1
X_08757_ net1052 team_03_WB.instance_to_wrap.core.register_file.registers_state\[707\]
+ net1004 team_03_WB.instance_to_wrap.core.register_file.registers_state\[739\] net926
+ vssd1 vssd1 vccd1 vccd1 _04699_ sky130_fd_sc_hd__a221o_1
Xhold1177 team_03_WB.instance_to_wrap.core.register_file.registers_state\[594\] vssd1
+ vssd1 vccd1 vccd1 net2670 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1188 team_03_WB.instance_to_wrap.core.register_file.registers_state\[515\] vssd1
+ vssd1 vccd1 vccd1 net2681 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout740_A net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout361_X net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1199 team_03_WB.instance_to_wrap.core.register_file.registers_state\[92\] vssd1
+ vssd1 vccd1 vccd1 net2692 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_239 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout459_X net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout838_A net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07708_ net747 _03648_ _03649_ net809 vssd1 vssd1 vccd1 vccd1 _03650_ sky130_fd_sc_hd__a31o_1
XFILLER_0_135_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11825__A1 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08688_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[872\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[840\]
+ net975 vssd1 vssd1 vccd1 vccd1 _04630_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_120_2835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08151__C1 net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_2846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07639_ net1192 team_03_WB.instance_to_wrap.core.register_file.registers_state\[494\]
+ net881 _03580_ vssd1 vssd1 vccd1 vccd1 _03581_ sky130_fd_sc_hd__a31o_1
XFILLER_0_95_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1270_X net1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout626_X net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_172_3902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11006__A net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_172_3913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10650_ team_03_WB.instance_to_wrap.core.decoder.inst\[11\] team_03_WB.instance_to_wrap.CPU_DAT_O\[11\]
+ net847 vssd1 vssd1 vccd1 vccd1 _02478_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09309_ net609 _05126_ vssd1 vssd1 vccd1 vccd1 _05251_ sky130_fd_sc_hd__nor2_1
XFILLER_0_134_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10581_ net1661 net532 net599 _03458_ vssd1 vssd1 vccd1 vccd1 _02542_ sky130_fd_sc_hd__a22o_1
XFILLER_0_63_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_999 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12320_ net1399 vssd1 vssd1 vccd1 vccd1 _00084_ sky130_fd_sc_hd__inv_2
XFILLER_0_145_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_556 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout995_X net995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_2797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_39_Left_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12002__A1 net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12251_ net1362 vssd1 vssd1 vccd1 vccd1 _00015_ sky130_fd_sc_hd__inv_2
XFILLER_0_32_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11379__C net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10013__A0 _03103_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08757__A1 net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11202_ net279 net2396 net486 vssd1 vssd1 vccd1 vccd1 _02206_ sky130_fd_sc_hd__mux2_1
X_12182_ net1604 vssd1 vssd1 vccd1 vccd1 _02371_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__11761__B1 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11133_ net2158 net415 _06642_ net512 vssd1 vssd1 vccd1 vccd1 _02237_ sky130_fd_sc_hd__a22o_1
XFILLER_0_43_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08509__A1 net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11064_ net1248 _06449_ net629 _06463_ vssd1 vssd1 vccd1 vccd1 _06610_ sky130_fd_sc_hd__or4_4
XANTENNA__11395__B net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10015_ net78 net67 net92 net89 vssd1 vssd1 vccd1 vccd1 _05893_ sky130_fd_sc_hd__or4_1
XANTENNA__08390__C1 net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_48_Left_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07732__A2 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14823_ clknet_leaf_102_wb_clk_i net1685 _01188_ vssd1 vssd1 vccd1 vccd1 net143 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_116_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14754_ clknet_leaf_47_wb_clk_i _02518_ _01119_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08196__S net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11966_ net642 _06743_ net477 net366 net1792 vssd1 vssd1 vccd1 vccd1 _01577_ sky130_fd_sc_hd__a32o_1
XFILLER_0_168_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_157_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10917_ net691 _05686_ net585 vssd1 vssd1 vccd1 vccd1 _06506_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_129_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13705_ clknet_leaf_77_wb_clk_i _01469_ _00070_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[59\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_80_2020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07496__A1 net1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14685_ clknet_leaf_65_wb_clk_i _02449_ _01050_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.ADR_I\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11292__A2 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11897_ net624 _06706_ net452 net371 net2184 vssd1 vssd1 vccd1 vccd1 _01644_ sky130_fd_sc_hd__a32o_1
XFILLER_0_132_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13636_ net1405 vssd1 vssd1 vccd1 vccd1 _01400_ sky130_fd_sc_hd__inv_2
XFILLER_0_156_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_37 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10848_ _06381_ _06390_ vssd1 vssd1 vccd1 vccd1 _06447_ sky130_fd_sc_hd__nor2_1
XFILLER_0_116_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09920__C_N _05583_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13567_ net1420 vssd1 vssd1 vccd1 vccd1 _01331_ sky130_fd_sc_hd__inv_2
X_10779_ net1042 _02808_ _06388_ vssd1 vssd1 vccd1 vccd1 _06389_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_137_692 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08996__A1 net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07799__A2 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_57_Left_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_180 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08540__S0 net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12518_ net1300 vssd1 vssd1 vccd1 vccd1 _00282_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13498_ net1340 vssd1 vssd1 vccd1 vccd1 _01262_ sky130_fd_sc_hd__inv_2
XFILLER_0_70_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12449_ net1281 vssd1 vssd1 vccd1 vccd1 _00213_ sky130_fd_sc_hd__inv_2
XANTENNA__12970__A net1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11289__C _06536_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_1128 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11752__B1 net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07956__C1 net1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14119_ clknet_leaf_113_wb_clk_i _01883_ _00484_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[473\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07783__B _03724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15099_ net1482 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[4] sky130_fd_sc_hd__buf_2
XANTENNA__07420__B2 net1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07990_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[944\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[912\]
+ net782 vssd1 vssd1 vccd1 vccd1 _03932_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06941_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[932\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[900\]
+ net776 vssd1 vssd1 vccd1 vccd1 _02883_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_52_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_52_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_66_Left_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09660_ net575 _05601_ vssd1 vssd1 vccd1 vccd1 _05602_ sky130_fd_sc_hd__nand2_1
XFILLER_0_59_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06872_ _02811_ _02813_ vssd1 vssd1 vccd1 vccd1 _02814_ sky130_fd_sc_hd__nor2_2
XANTENNA__07184__B1 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08611_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[5\] net1011
+ net931 _04552_ vssd1 vssd1 vccd1 vccd1 _04553_ sky130_fd_sc_hd__o211a_1
XANTENNA__07723__A2 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09591_ _05393_ _05418_ net569 vssd1 vssd1 vccd1 vccd1 _05533_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_141_3271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_32_wb_clk_i_A clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_08542_ net1229 team_03_WB.instance_to_wrap.core.register_file.registers_state\[734\]
+ net956 team_03_WB.instance_to_wrap.core.register_file.registers_state\[766\] net1210
+ vssd1 vssd1 vccd1 vccd1 _04484_ sky130_fd_sc_hd__o221a_1
XANTENNA__07304__A net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08473_ net850 _04414_ _04401_ vssd1 vssd1 vccd1 vccd1 _04415_ sky130_fd_sc_hd__o21a_4
XFILLER_0_159_283 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10491__B1 net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07424_ net1086 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1012\]
+ net889 _03365_ net1150 vssd1 vssd1 vccd1 vccd1 _03366_ sky130_fd_sc_hd__o311a_1
XFILLER_0_174_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07239__A1 net1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_75_Left_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07355_ net1172 team_03_WB.instance_to_wrap.core.register_file.registers_state\[604\]
+ net759 team_03_WB.instance_to_wrap.core.register_file.registers_state\[636\] net725
+ vssd1 vssd1 vccd1 vccd1 _03297_ sky130_fd_sc_hd__o221a_1
XFILLER_0_116_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1063_A net1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout419_A _06610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08987__A1 net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_476 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13041__A net1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07286_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[137\] net788
+ net735 _03227_ vssd1 vssd1 vccd1 vccd1 _03228_ sky130_fd_sc_hd__a211o_1
XANTENNA__11991__A0 net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_143_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09025_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[432\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[400\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[304\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[272\]
+ net984 net1079 vssd1 vssd1 vccd1 vccd1 _04967_ sky130_fd_sc_hd__mux4_1
XFILLER_0_103_515 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1230_A net1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09936__A0 _05872_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1328_A net1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_1933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_1944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold230 team_03_WB.instance_to_wrap.core.register_file.registers_state\[819\] vssd1
+ vssd1 vccd1 vccd1 net1723 sky130_fd_sc_hd__dlygate4sd3_1
Xhold241 net190 vssd1 vssd1 vccd1 vccd1 net1734 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_148_3414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold252 team_03_WB.instance_to_wrap.core.register_file.registers_state\[395\] vssd1
+ vssd1 vccd1 vccd1 net1745 sky130_fd_sc_hd__dlygate4sd3_1
Xhold263 team_03_WB.instance_to_wrap.core.register_file.registers_state\[46\] vssd1
+ vssd1 vccd1 vccd1 net1756 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout788_A net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold274 net213 vssd1 vssd1 vccd1 vccd1 net1767 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10604__S net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_2694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold285 team_03_WB.instance_to_wrap.core.register_file.registers_state\[966\] vssd1
+ vssd1 vccd1 vccd1 net1778 sky130_fd_sc_hd__dlygate4sd3_1
Xhold296 team_03_WB.instance_to_wrap.core.register_file.registers_state\[572\] vssd1
+ vssd1 vccd1 vccd1 net1789 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout710 net711 vssd1 vssd1 vccd1 vccd1 net710 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout1116_X net1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout721 _02863_ vssd1 vssd1 vccd1 vccd1 net721 sky130_fd_sc_hd__buf_6
XANTENNA__07962__A2 _03900_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout732 net733 vssd1 vssd1 vccd1 vccd1 net732 sky130_fd_sc_hd__buf_2
X_09927_ _03638_ net663 vssd1 vssd1 vccd1 vccd1 _05868_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_165_3761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_71_wb_clk_i_A clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_165_3772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout743 net745 vssd1 vssd1 vccd1 vccd1 net743 sky130_fd_sc_hd__buf_4
Xfanout754 net755 vssd1 vssd1 vccd1 vccd1 net754 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout955_A net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout765 net773 vssd1 vssd1 vccd1 vccd1 net765 sky130_fd_sc_hd__buf_2
Xfanout776 net777 vssd1 vssd1 vccd1 vccd1 net776 sky130_fd_sc_hd__buf_2
X_09858_ _05768_ _05784_ _05798_ vssd1 vssd1 vccd1 vccd1 _05800_ sky130_fd_sc_hd__or3_1
Xfanout787 net788 vssd1 vssd1 vccd1 vccd1 net787 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_102_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06877__X _02819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout798 net805 vssd1 vssd1 vccd1 vccd1 net798 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08911__A1 net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07714__A2 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08372__C1 net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08809_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[417\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[385\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[289\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[257\]
+ net981 net1076 vssd1 vssd1 vccd1 vccd1 _04751_ sky130_fd_sc_hd__mux4_1
X_09789_ _05250_ _05269_ _05246_ vssd1 vssd1 vccd1 vccd1 _05731_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout743_X net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11820_ net650 _06650_ net461 net324 net1868 vssd1 vssd1 vccd1 vccd1 _01719_ sky130_fd_sc_hd__a32o_1
XFILLER_0_96_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout910_X net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11751_ _06574_ net463 net332 net2285 vssd1 vssd1 vccd1 vccd1 _01786_ sky130_fd_sc_hd__a22o_1
XANTENNA__11274__A2 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_732 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10702_ _06311_ _06337_ net603 vssd1 vssd1 vccd1 vccd1 _06340_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_139_968 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10482__B1 net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14470_ clknet_leaf_72_wb_clk_i _02234_ _00835_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[824\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_154_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11682_ _06724_ net381 net338 net1992 vssd1 vssd1 vccd1 vccd1 _01852_ sky130_fd_sc_hd__a22o_1
XFILLER_0_37_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13421_ net1415 vssd1 vssd1 vccd1 vccd1 _01185_ sky130_fd_sc_hd__inv_2
X_10633_ team_03_WB.instance_to_wrap.core.decoder.inst\[28\] net2391 net844 vssd1
+ vssd1 vccd1 vccd1 _02495_ sky130_fd_sc_hd__mux2_1
XANTENNA__08427__B1 net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11026__A2 net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_990 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13352_ net1318 vssd1 vssd1 vccd1 vccd1 _01116_ sky130_fd_sc_hd__inv_2
Xmax_cap1016 net1017 vssd1 vssd1 vccd1 vccd1 net1016 sky130_fd_sc_hd__dlymetal6s2s_1
X_10564_ net1716 net531 net598 _05874_ vssd1 vssd1 vccd1 vccd1 _02559_ sky130_fd_sc_hd__a22o_1
XANTENNA_input84_A wbs_adr_i[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11982__A0 _06434_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12303_ net1394 vssd1 vssd1 vccd1 vccd1 _00067_ sky130_fd_sc_hd__inv_2
XFILLER_0_162_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13283_ net1345 vssd1 vssd1 vccd1 vccd1 _01047_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_20_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10495_ net105 net1030 net907 net1673 vssd1 vssd1 vccd1 vccd1 _02614_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_20_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12790__A net1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15022_ clknet_leaf_92_wb_clk_i _02742_ _01387_ vssd1 vssd1 vccd1 vccd1 net178 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_133_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12234_ net1625 vssd1 vssd1 vccd1 vccd1 _01423_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__07884__A net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_833 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11734__B1 _06808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_378 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12165_ net1576 vssd1 vssd1 vccd1 vccd1 _02388_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_9_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11116_ net835 _06550_ vssd1 vssd1 vccd1 vccd1 _06632_ sky130_fd_sc_hd__and2_1
XANTENNA__07953__A2 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12096_ _06793_ net478 net442 net1884 vssd1 vssd1 vccd1 vccd1 _01451_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_30_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11047_ net643 _06600_ vssd1 vssd1 vccd1 vccd1 _06601_ sky130_fd_sc_hd__nor2_1
XFILLER_0_127_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08363__C1 net1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput9 DAT_I[16] vssd1 vssd1 vccd1 vccd1 net9 sky130_fd_sc_hd__clkbuf_1
XANTENNA__09604__A _05545_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06913__B1 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14806_ clknet_leaf_56_wb_clk_i _02570_ _01171_ vssd1 vssd1 vccd1 vccd1 net171 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11572__C net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12998_ net1294 vssd1 vssd1 vccd1 vccd1 _00762_ sky130_fd_sc_hd__inv_2
X_14737_ clknet_leaf_33_wb_clk_i _02501_ _01102_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08666__B1 net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11949_ net640 _06726_ net475 net363 net1835 vssd1 vssd1 vccd1 vccd1 _01594_ sky130_fd_sc_hd__a32o_1
XFILLER_0_143_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_116_wb_clk_i_A clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_28_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_89 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14668_ clknet_leaf_15_wb_clk_i _02432_ _01033_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1022\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_156_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_966 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13619_ net1431 vssd1 vssd1 vccd1 vccd1 _01383_ sky130_fd_sc_hd__inv_2
XFILLER_0_171_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14599_ clknet_leaf_110_wb_clk_i _02363_ _00964_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[953\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_116_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07140_ net1104 team_03_WB.instance_to_wrap.core.register_file.registers_state\[32\]
+ net901 vssd1 vssd1 vccd1 vccd1 _03082_ sky130_fd_sc_hd__or3_1
XFILLER_0_15_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11973__B1 net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07071_ net1097 team_03_WB.instance_to_wrap.core.register_file.registers_state\[194\]
+ net797 team_03_WB.instance_to_wrap.core.register_file.registers_state\[226\] net733
+ vssd1 vssd1 vccd1 vccd1 _03013_ sky130_fd_sc_hd__a221o_1
XANTENNA__07641__B2 net1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_2277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10528__A1 net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10932__B _06517_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_2288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11725__B1 _06808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10424__S net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_71_1830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11740__A3 net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_1841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07973_ net1203 team_03_WB.instance_to_wrap.core.register_file.registers_state\[336\]
+ vssd1 vssd1 vccd1 vccd1 _03915_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_143_3311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09712_ net583 _04775_ vssd1 vssd1 vccd1 vccd1 _05654_ sky130_fd_sc_hd__or2_1
XANTENNA__08121__C net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06924_ net1106 team_03_WB.instance_to_wrap.core.register_file.registers_state\[324\]
+ net1157 vssd1 vssd1 vccd1 vccd1 _02866_ sky130_fd_sc_hd__a21o_1
XANTENNA__07157__B1 _02872_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09643_ _05185_ _05501_ _05192_ vssd1 vssd1 vccd1 vccd1 _05585_ sky130_fd_sc_hd__a21oi_1
X_06855_ team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[29\] vssd1 vssd1 vccd1
+ vccd1 _02798_ sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_155_wb_clk_i_A clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout271_A _06491_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout369_A _06814_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_1032 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09574_ net352 _05508_ _05515_ vssd1 vssd1 vccd1 vccd1 _05516_ sky130_fd_sc_hd__a21o_1
XFILLER_0_167_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07034__A net1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08525_ net854 _04465_ _04466_ vssd1 vssd1 vccd1 vccd1 _04467_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_69_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11256__A2 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08657__B1 net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout536_A net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12875__A net1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1180_A net1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_743 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_120 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1278_A net1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08456_ net1228 team_03_WB.instance_to_wrap.core.register_file.registers_state\[860\]
+ net953 team_03_WB.instance_to_wrap.core.register_file.registers_state\[892\] net1218
+ vssd1 vssd1 vccd1 vccd1 _04398_ sky130_fd_sc_hd__o221a_1
XANTENNA__07969__A net1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08564__S net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_148_787 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07407_ net1146 _03347_ _03348_ net1160 _03346_ vssd1 vssd1 vccd1 vccd1 _03349_ sky130_fd_sc_hd__o311a_1
XFILLER_0_92_346 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07880__A1 team_03_WB.instance_to_wrap.core.decoder.inst\[27\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08387_ net1245 team_03_WB.instance_to_wrap.core.register_file.registers_state\[185\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[153\] net992 net931
+ vssd1 vssd1 vccd1 vccd1 _04329_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout324_X net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout703_A net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1066_X net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07338_ _03277_ _03279_ net610 vssd1 vssd1 vccd1 vccd1 _03280_ sky130_fd_sc_hd__mux2_2
XFILLER_0_144_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_150_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11964__B1 net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_2734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11003__B net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07269_ net1205 team_03_WB.instance_to_wrap.core.register_file.registers_state\[969\]
+ vssd1 vssd1 vccd1 vccd1 _03211_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_115_2745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1233_X net1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_788 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09008_ net917 _04947_ _04948_ net860 vssd1 vssd1 vccd1 vccd1 _04950_ sky130_fd_sc_hd__a211o_1
XFILLER_0_103_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_167_3801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10280_ _03822_ _06117_ _06121_ vssd1 vssd1 vccd1 vccd1 _06122_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_131_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_167_3812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout693_X net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout860_X net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout540 _04815_ vssd1 vssd1 vccd1 vccd1 net540 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout958_X net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout551 net552 vssd1 vssd1 vccd1 vccd1 net551 sky130_fd_sc_hd__clkbuf_2
Xfanout562 _03063_ vssd1 vssd1 vccd1 vccd1 net562 sky130_fd_sc_hd__clkbuf_4
Xfanout573 net577 vssd1 vssd1 vccd1 vccd1 net573 sky130_fd_sc_hd__clkbuf_4
X_13970_ clknet_leaf_165_wb_clk_i _01734_ _00335_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[324\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout584 _02891_ vssd1 vssd1 vccd1 vccd1 net584 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07148__B1 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout595 _02951_ vssd1 vssd1 vccd1 vccd1 net595 sky130_fd_sc_hd__buf_4
XANTENNA__07699__A1 _03640_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12921_ net1359 vssd1 vssd1 vccd1 vccd1 _00685_ sky130_fd_sc_hd__inv_2
XANTENNA__08896__B1 net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12852_ net1306 vssd1 vssd1 vccd1 vccd1 _00616_ sky130_fd_sc_hd__inv_2
XFILLER_0_69_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11803_ net2509 _06630_ net330 vssd1 vssd1 vccd1 vccd1 _01735_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_1127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12783_ net1394 vssd1 vssd1 vccd1 vccd1 _00547_ sky130_fd_sc_hd__inv_2
XANTENNA__10857__X _06456_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08982__B net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11734_ net596 _06519_ net464 _06808_ net1807 vssd1 vssd1 vccd1 vccd1 _01802_ sky130_fd_sc_hd__a32o_1
X_14522_ clknet_leaf_142_wb_clk_i _02286_ _00887_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[876\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_68_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07320__B1 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_154_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11665_ net2103 _06627_ net342 vssd1 vssd1 vccd1 vccd1 _01868_ sky130_fd_sc_hd__mux2_1
X_14453_ clknet_leaf_107_wb_clk_i _02217_ _00818_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[807\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07871__A1 net1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13404_ net1321 vssd1 vssd1 vccd1 vccd1 _01168_ sky130_fd_sc_hd__inv_2
X_10616_ net1668 team_03_WB.instance_to_wrap.CPU_DAT_O\[13\] net843 vssd1 vssd1 vccd1
+ vccd1 _02512_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14384_ clknet_leaf_155_wb_clk_i _02148_ _00749_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[738\]
+ sky130_fd_sc_hd__dfrtp_1
X_11596_ _06504_ net2223 net447 vssd1 vssd1 vccd1 vccd1 _01933_ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_1056 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_418 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11955__B1 net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13335_ net1308 vssd1 vssd1 vccd1 vccd1 _01099_ sky130_fd_sc_hd__inv_2
XFILLER_0_109_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10547_ team_03_WB.instance_to_wrap.wb.curr_state\[0\] _06284_ _06289_ vssd1 vssd1
+ vccd1 vccd1 _06291_ sky130_fd_sc_hd__o21a_1
XFILLER_0_122_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_479 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_952 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13266_ net1398 vssd1 vssd1 vccd1 vccd1 _01030_ sky130_fd_sc_hd__inv_2
XANTENNA__11970__A3 net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10478_ net123 net1027 net905 net1640 vssd1 vssd1 vccd1 vccd1 _02631_ sky130_fd_sc_hd__a22o_1
XANTENNA__10752__B net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08503__A _04444_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_985 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11707__B1 net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15005_ clknet_leaf_51_wb_clk_i net53 _01370_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_12217_ net1607 vssd1 vssd1 vccd1 vccd1 _01440_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__11567__C net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13197_ net1294 vssd1 vssd1 vccd1 vccd1 _00961_ sky130_fd_sc_hd__inv_2
XANTENNA__07387__B1 net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11183__B2 net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12148_ net1581 vssd1 vssd1 vccd1 vccd1 _02405_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_10_Right_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12079_ net626 _06643_ net460 net440 net1958 vssd1 vssd1 vccd1 vccd1 _01468_ sky130_fd_sc_hd__a32o_1
XANTENNA__08649__S net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07139__B1 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_139_Right_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11075__S net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11238__A2 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10767__X _06378_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08892__B net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_47_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09300__A1 net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08310_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[952\] net973
+ vssd1 vssd1 vccd1 vccd1 _04252_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_47_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11803__S net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09290_ _05228_ _05230_ vssd1 vssd1 vccd1 vccd1 _05232_ sky130_fd_sc_hd__nand2_1
XANTENNA__07311__B1 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08241_ net934 _04181_ _04182_ vssd1 vssd1 vccd1 vccd1 _04183_ sky130_fd_sc_hd__o21a_1
XFILLER_0_118_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_459 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11104__A net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_136_3170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08172_ net1061 _04111_ _04113_ net1071 vssd1 vssd1 vccd1 vccd1 _04114_ sky130_fd_sc_hd__a211o_1
XFILLER_0_16_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09064__B1 net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_95_2328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_1107 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11946__B1 net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07123_ net1189 net1016 _02835_ net1252 vssd1 vssd1 vccd1 vccd1 _03065_ sky130_fd_sc_hd__a22oi_4
XANTENNA__07614__A1 net1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07020__C net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10943__A net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_3078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_939 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_852 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_3089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_99_wb_clk_i clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_99_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_07054_ net1095 team_03_WB.instance_to_wrap.core.register_file.registers_state\[834\]
+ net796 team_03_WB.instance_to_wrap.core.register_file.registers_state\[866\] net1154
+ vssd1 vssd1 vccd1 vccd1 _02996_ sky130_fd_sc_hd__a221o_1
Xoutput110 net110 vssd1 vssd1 vccd1 vccd1 ADR_O[16] sky130_fd_sc_hd__clkbuf_4
XANTENNA__11961__A3 net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput121 net121 vssd1 vssd1 vccd1 vccd1 ADR_O[26] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_101_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput132 net132 vssd1 vssd1 vccd1 vccd1 ADR_O[7] sky130_fd_sc_hd__clkbuf_4
Xoutput143 net143 vssd1 vssd1 vccd1 vccd1 DAT_O[16] sky130_fd_sc_hd__buf_2
XFILLER_0_112_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_28_wb_clk_i clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_28_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xoutput154 net154 vssd1 vssd1 vccd1 vccd1 DAT_O[26] sky130_fd_sc_hd__clkbuf_4
Xoutput165 net165 vssd1 vssd1 vccd1 vccd1 DAT_O[7] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_110_2631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11174__A1 net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11477__C _06527_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1026_A _06286_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_2642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07378__B1 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput176 net176 vssd1 vssd1 vccd1 vccd1 gpio_oeb[11] sky130_fd_sc_hd__buf_2
XFILLER_0_11_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07917__A2 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput187 net187 vssd1 vssd1 vccd1 vccd1 gpio_oeb[22] sky130_fd_sc_hd__buf_2
Xoutput198 net198 vssd1 vssd1 vccd1 vccd1 gpio_oeb[33] sky130_fd_sc_hd__clkbuf_4
XANTENNA__11196__D net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout486_A _06680_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07956_ net729 _03886_ _03887_ net1147 vssd1 vssd1 vccd1 vccd1 _03898_ sky130_fd_sc_hd__a211o_1
XANTENNA__09244__A _04119_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06907_ net1164 net882 vssd1 vssd1 vccd1 vccd1 _02849_ sky130_fd_sc_hd__nand2_1
X_07887_ net1090 team_03_WB.instance_to_wrap.core.register_file.registers_state\[79\]
+ vssd1 vssd1 vccd1 vccd1 _03829_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout653_A net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_106_Right_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1395_A net1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09626_ _03024_ _05483_ _05567_ vssd1 vssd1 vccd1 vccd1 _05568_ sky130_fd_sc_hd__a21oi_2
X_06838_ team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[8\] vssd1 vssd1 vccd1
+ vccd1 _02781_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_108_2593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09557_ net594 _05430_ _05480_ _05498_ vssd1 vssd1 vccd1 vccd1 _05499_ sky130_fd_sc_hd__o31a_1
XANTENNA_fanout441_X net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1183_X net1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout539_X net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout918_A net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11713__S net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08508_ net1045 team_03_WB.instance_to_wrap.core.register_file.registers_state\[671\]
+ net995 team_03_WB.instance_to_wrap.core.register_file.registers_state\[703\] net916
+ vssd1 vssd1 vccd1 vccd1 _04450_ sky130_fd_sc_hd__a221o_1
XFILLER_0_37_1090 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09488_ _05306_ _05307_ _05311_ _05329_ vssd1 vssd1 vccd1 vccd1 _05430_ sky130_fd_sc_hd__o31a_1
XFILLER_0_109_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10988__B2 net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_156_3568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08439_ net867 _04380_ _04375_ net851 vssd1 vssd1 vccd1 vccd1 _04381_ sky130_fd_sc_hd__o211a_1
XANTENNA__10329__S net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_156_3579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout706_X net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11450_ net626 _06575_ vssd1 vssd1 vccd1 vccd1 _06764_ sky130_fd_sc_hd__and2_1
XFILLER_0_151_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_163_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10401_ net284 _06226_ vssd1 vssd1 vccd1 vccd1 _06227_ sky130_fd_sc_hd__nand2_1
XANTENNA__09150__S0 net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08802__B1 net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11381_ net715 net295 net699 vssd1 vssd1 vccd1 vccd1 _06743_ sky130_fd_sc_hd__and3_1
XFILLER_0_150_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13120_ net1402 vssd1 vssd1 vccd1 vccd1 _00884_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_12_Left_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10332_ _05975_ _06111_ _06116_ _06114_ vssd1 vssd1 vccd1 vccd1 _06170_ sky130_fd_sc_hd__a31o_1
XANTENNA__09419__A _04820_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11952__A3 net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_484 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13051_ net1364 vssd1 vssd1 vccd1 vccd1 _00815_ sky130_fd_sc_hd__inv_2
X_10263_ _06097_ _06100_ _06096_ vssd1 vssd1 vccd1 vccd1 _06105_ sky130_fd_sc_hd__a21bo_1
XANTENNA__11387__C _06536_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12002_ net264 _06756_ net474 net444 net2128 vssd1 vssd1 vccd1 vccd1 _01542_ sky130_fd_sc_hd__a32o_1
Xfanout1302 net1438 vssd1 vssd1 vccd1 vccd1 net1302 sky130_fd_sc_hd__buf_2
XANTENNA__08030__A1 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10194_ _04565_ net676 _06033_ _02893_ vssd1 vssd1 vccd1 vccd1 _06036_ sky130_fd_sc_hd__o211a_1
XANTENNA_input47_A gpio_in[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1313 net1315 vssd1 vssd1 vccd1 vccd1 net1313 sky130_fd_sc_hd__buf_4
XFILLER_0_79_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1324 net1330 vssd1 vssd1 vccd1 vccd1 net1324 sky130_fd_sc_hd__buf_2
Xfanout1335 net1339 vssd1 vssd1 vccd1 vccd1 net1335 sky130_fd_sc_hd__buf_2
Xfanout1346 net1438 vssd1 vssd1 vccd1 vccd1 net1346 sky130_fd_sc_hd__clkbuf_4
Xfanout1357 net1358 vssd1 vssd1 vccd1 vccd1 net1357 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_17_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout370 _06814_ vssd1 vssd1 vccd1 vccd1 net370 sky130_fd_sc_hd__buf_4
Xfanout1368 net1369 vssd1 vssd1 vccd1 vccd1 net1368 sky130_fd_sc_hd__buf_4
Xfanout1379 net1380 vssd1 vssd1 vccd1 vccd1 net1379 sky130_fd_sc_hd__buf_4
Xfanout381 net387 vssd1 vssd1 vccd1 vccd1 net381 sky130_fd_sc_hd__buf_4
Xfanout392 net395 vssd1 vssd1 vccd1 vccd1 net392 sky130_fd_sc_hd__buf_6
X_13953_ clknet_leaf_184_wb_clk_i _01717_ _00318_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[307\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09530__A1 net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_21_Left_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12904_ net1299 vssd1 vssd1 vccd1 vccd1 _00668_ sky130_fd_sc_hd__inv_2
X_13884_ clknet_leaf_149_wb_clk_i _01648_ _00249_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[238\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08993__A net1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_326 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12835_ net1371 vssd1 vssd1 vccd1 vccd1 _00599_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_1106 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10428__B1 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08097__A1 net1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12766_ net1409 vssd1 vssd1 vccd1 vccd1 _00530_ sky130_fd_sc_hd__inv_2
XFILLER_0_68_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14505_ clknet_leaf_75_wb_clk_i _02269_ _00870_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[859\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07402__A net1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11717_ net2006 net277 net336 vssd1 vssd1 vccd1 vccd1 _01819_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12697_ net1357 vssd1 vssd1 vccd1 vccd1 _00461_ sky130_fd_sc_hd__inv_2
XANTENNA__11640__A2 net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11648_ net2271 _06614_ net344 vssd1 vssd1 vccd1 vccd1 _01885_ sky130_fd_sc_hd__mux2_1
X_14436_ clknet_leaf_23_wb_clk_i _02200_ _00801_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[790\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_64_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput12 DAT_I[19] vssd1 vssd1 vccd1 vccd1 net12 sky130_fd_sc_hd__buf_1
Xinput23 DAT_I[29] vssd1 vssd1 vccd1 vccd1 net23 sky130_fd_sc_hd__buf_1
Xinput34 gpio_in[0] vssd1 vssd1 vccd1 vccd1 net34 sky130_fd_sc_hd__clkbuf_1
Xinput45 gpio_in[20] vssd1 vssd1 vccd1 vccd1 net45 sky130_fd_sc_hd__clkbuf_1
XANTENNA__10763__A _05798_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14367_ clknet_leaf_172_wb_clk_i _02131_ _00732_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[721\]
+ sky130_fd_sc_hd__dfrtp_1
X_11579_ net279 net2417 net447 vssd1 vssd1 vccd1 vccd1 _01950_ sky130_fd_sc_hd__mux2_1
Xinput56 gpio_in[31] vssd1 vssd1 vccd1 vccd1 net56 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput67 wbs_adr_i[0] vssd1 vssd1 vccd1 vccd1 net67 sky130_fd_sc_hd__buf_1
Xhold807 team_03_WB.instance_to_wrap.core.register_file.registers_state\[574\] vssd1
+ vssd1 vccd1 vccd1 net2300 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput78 wbs_adr_i[1] vssd1 vssd1 vccd1 vccd1 net78 sky130_fd_sc_hd__clkbuf_1
X_13318_ net1342 vssd1 vssd1 vccd1 vccd1 _01082_ sky130_fd_sc_hd__inv_2
Xhold818 team_03_WB.instance_to_wrap.core.register_file.registers_state\[769\] vssd1
+ vssd1 vccd1 vccd1 net2311 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11943__A3 net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput89 wbs_adr_i[2] vssd1 vssd1 vccd1 vccd1 net89 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_126_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold829 team_03_WB.instance_to_wrap.core.register_file.registers_state\[716\] vssd1
+ vssd1 vccd1 vccd1 net2322 sky130_fd_sc_hd__dlygate4sd3_1
X_14298_ clknet_leaf_146_wb_clk_i _02062_ _00663_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[652\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07775__C net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_90_2225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13249_ net1260 vssd1 vssd1 vccd1 vccd1 _01013_ sky130_fd_sc_hd__inv_2
XANTENNA__11297__C net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11156__B2 net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08557__C1 net1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08021__A1 net1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07810_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[427\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[395\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[299\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[267\]
+ net775 net1126 vssd1 vssd1 vccd1 vccd1 _03752_ sky130_fd_sc_hd__mux4_1
X_08790_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[546\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[514\]
+ net977 vssd1 vssd1 vccd1 vccd1 _04732_ sky130_fd_sc_hd__mux2_1
XANTENNA__12105__B1 net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08309__C1 net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07780__B1 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07741_ net1194 net883 _02796_ vssd1 vssd1 vccd1 vccd1 _03683_ sky130_fd_sc_hd__a21o_1
XANTENNA__11459__A2 net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_2176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_2187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_146_wb_clk_i clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_146_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_07672_ net811 _03609_ _03610_ _03613_ vssd1 vssd1 vccd1 vccd1 _03614_ sky130_fd_sc_hd__o22a_1
XFILLER_0_79_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09411_ _05351_ _05352_ net554 vssd1 vssd1 vccd1 vccd1 _05353_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07015__C net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09342_ _04207_ _05282_ vssd1 vssd1 vccd1 vccd1 _05284_ sky130_fd_sc_hd__nand2_1
XANTENNA__08088__A1 net1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_3210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_2490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09273_ _03790_ _05214_ vssd1 vssd1 vccd1 vccd1 _05215_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_30_1127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07835__A1 net1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11631__A2 net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_134_3118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09938__S net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_134_3129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08224_ net1061 _04165_ _04164_ net1071 vssd1 vssd1 vccd1 vccd1 _04166_ sky130_fd_sc_hd__a211o_1
XFILLER_0_62_338 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08155_ team_03_WB.instance_to_wrap.core.decoder.inst\[19\] _02820_ vssd1 vssd1 vccd1
+ vccd1 _04097_ sky130_fd_sc_hd__nand2_4
XFILLER_0_126_790 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout401_A _06718_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_160_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1143_A net1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_151_3476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10198__A2 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11121__X _06635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07106_ net1165 _03047_ vssd1 vssd1 vccd1 vccd1 _03048_ sky130_fd_sc_hd__nand2_1
X_08086_ net1147 _04017_ _04027_ vssd1 vssd1 vccd1 vccd1 _04028_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_140_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07037_ net1099 team_03_WB.instance_to_wrap.core.register_file.registers_state\[67\]
+ net801 team_03_WB.instance_to_wrap.core.register_file.registers_state\[99\] net748
+ vssd1 vssd1 vccd1 vccd1 _02979_ sky130_fd_sc_hd__a221o_1
XANTENNA__11147__A1 net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1029_X net1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1408_A net1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08012__A1 net1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11698__A2 net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout770_A net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout391_X net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout489_X net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout868_A net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09760__A1 _04777_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10612__S net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08289__S net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08988_ net859 _04928_ _04929_ vssd1 vssd1 vccd1 vccd1 _04930_ sky130_fd_sc_hd__and3_1
XFILLER_0_138_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07939_ net1128 _03877_ _03878_ net1116 vssd1 vssd1 vccd1 vccd1 _03881_ sky130_fd_sc_hd__a211oi_1
XANTENNA_fanout656_X net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_127_2980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11009__A net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1398_X net1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10950_ team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[4\] net306 vssd1 vssd1
+ vccd1 vccd1 _06533_ sky130_fd_sc_hd__and2_1
XFILLER_0_138_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_127_2991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09609_ net568 _04535_ vssd1 vssd1 vccd1 vccd1 _05551_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_27_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_158_3619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10881_ net692 _06475_ _06476_ _06474_ vssd1 vssd1 vccd1 vccd1 _06477_ sky130_fd_sc_hd__a31oi_4
XFILLER_0_39_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout823_X net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_123_2899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input101_A wbs_stb_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08079__A1 net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12620_ net1312 vssd1 vssd1 vccd1 vccd1 _00384_ sky130_fd_sc_hd__inv_2
XFILLER_0_149_860 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09276__B1 net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09815__A2 _05587_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11083__A0 _06619_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12551_ net1368 vssd1 vssd1 vccd1 vccd1 _00315_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11622__A2 net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11502_ _06621_ net2670 net388 vssd1 vssd1 vccd1 vccd1 _02004_ sky130_fd_sc_hd__mux2_1
X_12482_ net1359 vssd1 vssd1 vccd1 vccd1 _00246_ sky130_fd_sc_hd__inv_2
XFILLER_0_164_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_738 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_145_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09123__S0 net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14221_ clknet_leaf_183_wb_clk_i _01985_ _00586_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[575\]
+ sky130_fd_sc_hd__dfrtp_1
X_11433_ net267 net2662 net398 vssd1 vssd1 vccd1 vccd1 _02051_ sky130_fd_sc_hd__mux2_1
XANTENNA__11386__A1 net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_202 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08787__C1 net1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14152_ clknet_leaf_8_wb_clk_i _01916_ _00517_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[506\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_151_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11398__B _06751_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11364_ net511 net641 _06734_ net403 net2555 vssd1 vssd1 vccd1 vccd1 _02098_ sky130_fd_sc_hd__a32o_1
XFILLER_0_105_996 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10315_ _05969_ _06127_ _05970_ _05964_ vssd1 vssd1 vccd1 vccd1 _06156_ sky130_fd_sc_hd__a211o_1
XFILLER_0_132_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13103_ net1338 vssd1 vssd1 vccd1 vccd1 _00867_ sky130_fd_sc_hd__inv_2
X_14083_ clknet_leaf_31_wb_clk_i _01847_ _00448_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[437\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_104_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10870__X _06468_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11295_ net712 _06550_ net829 vssd1 vssd1 vccd1 vccd1 _06715_ sky130_fd_sc_hd__and3_1
XFILLER_0_21_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08988__A net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09436__X _05378_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13034_ net1279 vssd1 vssd1 vccd1 vccd1 _00798_ sky130_fd_sc_hd__inv_2
X_10246_ _05987_ _06087_ vssd1 vssd1 vccd1 vccd1 _06088_ sky130_fd_sc_hd__nor2_1
XFILLER_0_119_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11689__A2 net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1110 net1111 vssd1 vssd1 vccd1 vccd1 net1110 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09751__A1 _04816_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11167__C_N net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1121 net1122 vssd1 vssd1 vccd1 vccd1 net1121 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07211__C1 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1132 net1137 vssd1 vssd1 vccd1 vccd1 net1132 sky130_fd_sc_hd__clkbuf_4
X_10177_ _04922_ net675 vssd1 vssd1 vccd1 vccd1 _06019_ sky130_fd_sc_hd__or2_1
XANTENNA__08199__S net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1143 net1144 vssd1 vssd1 vccd1 vccd1 net1143 sky130_fd_sc_hd__buf_2
XANTENNA__10361__A2 net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1154 net1157 vssd1 vssd1 vccd1 vccd1 net1154 sky130_fd_sc_hd__buf_4
Xfanout1165 net1166 vssd1 vssd1 vccd1 vccd1 net1165 sky130_fd_sc_hd__buf_4
Xfanout1176 net1179 vssd1 vssd1 vccd1 vccd1 net1176 sky130_fd_sc_hd__clkbuf_4
X_14985_ clknet_leaf_66_wb_clk_i net64 _01350_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[4\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1187 net1188 vssd1 vssd1 vccd1 vccd1 net1187 sky130_fd_sc_hd__clkbuf_4
Xfanout1198 net1199 vssd1 vssd1 vccd1 vccd1 net1198 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10649__A0 team_03_WB.instance_to_wrap.core.decoder.inst\[12\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13936_ clknet_leaf_160_wb_clk_i _01700_ _00301_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[290\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_77_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08711__C1 net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09612__A net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13867_ clknet_leaf_41_wb_clk_i _01631_ _00232_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[221\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_2073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_83_2084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12818_ net1397 vssd1 vssd1 vccd1 vccd1 _00582_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13798_ clknet_leaf_73_wb_clk_i _01562_ _00163_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[152\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07817__A1 _03758_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_463 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12749_ net1332 vssd1 vssd1 vccd1 vccd1 _00513_ sky130_fd_sc_hd__inv_2
XANTENNA__11613__A2 net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10821__B1 net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09019__B1 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_142_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08490__A1 net1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08490__B2 net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09114__S0 net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_844 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14419_ clknet_leaf_97_wb_clk_i _02183_ _00784_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[773\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_13_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_511 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10924__C _05845_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07278__S net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08242__A1 net1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold604 team_03_WB.instance_to_wrap.core.register_file.registers_state\[226\] vssd1
+ vssd1 vccd1 vccd1 net2097 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold615 team_03_WB.instance_to_wrap.core.register_file.registers_state\[698\] vssd1
+ vssd1 vccd1 vccd1 net2108 sky130_fd_sc_hd__dlygate4sd3_1
Xwire590 _04984_ vssd1 vssd1 vccd1 vccd1 net590 sky130_fd_sc_hd__buf_4
Xhold626 team_03_WB.instance_to_wrap.core.register_file.registers_state\[543\] vssd1
+ vssd1 vccd1 vccd1 net2119 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold637 team_03_WB.instance_to_wrap.core.register_file.registers_state\[287\] vssd1
+ vssd1 vccd1 vccd1 net2130 sky130_fd_sc_hd__dlygate4sd3_1
Xhold648 team_03_WB.instance_to_wrap.core.register_file.registers_state\[849\] vssd1
+ vssd1 vccd1 vccd1 net2141 sky130_fd_sc_hd__dlygate4sd3_1
Xhold659 team_03_WB.instance_to_wrap.core.register_file.registers_state\[610\] vssd1
+ vssd1 vccd1 vccd1 net2152 sky130_fd_sc_hd__dlygate4sd3_1
X_09960_ _05884_ net1689 net291 vssd1 vssd1 vccd1 vccd1 _02747_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_38_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08911_ net942 _04852_ _04851_ net1065 vssd1 vssd1 vccd1 vccd1 _04853_ sky130_fd_sc_hd__o211a_1
X_09891_ _05825_ _05826_ _05832_ vssd1 vssd1 vccd1 vccd1 _05833_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_0_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07202__C1 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09742__B2 _04777_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08842_ net1056 team_03_WB.instance_to_wrap.core.register_file.registers_state\[64\]
+ net1009 team_03_WB.instance_to_wrap.core.register_file.registers_state\[96\] net946
+ vssd1 vssd1 vccd1 vccd1 _04784_ sky130_fd_sc_hd__a221o_1
XFILLER_0_100_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08773_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[2\] net1002
+ net925 _04714_ vssd1 vssd1 vccd1 vccd1 _04715_ sky130_fd_sc_hd__o211a_1
XFILLER_0_26_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07724_ net1193 team_03_WB.instance_to_wrap.core.register_file.registers_state\[685\]
+ net882 vssd1 vssd1 vccd1 vccd1 _03666_ sky130_fd_sc_hd__and3_1
XFILLER_0_79_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_105_2530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07505__B1 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_105_2541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07655_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[942\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[910\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[814\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[782\]
+ net774 net1131 vssd1 vssd1 vccd1 vccd1 _03597_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_0_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10668__A _05541_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1093_A _02787_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_216 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout449_A _06801_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07586_ net684 _03527_ vssd1 vssd1 vccd1 vccd1 _03528_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_101_2449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09325_ _05253_ _05266_ vssd1 vssd1 vccd1 vccd1 _05267_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_153_3516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1260_A net1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout616_A net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_11_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1358_A net1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10812__A0 _06418_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09256_ _05196_ _05197_ vssd1 vssd1 vccd1 vccd1 _05198_ sky130_fd_sc_hd__or2_1
XFILLER_0_62_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07284__A2 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09895__C net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06881__A team_03_WB.instance_to_wrap.core.decoder.inst\[14\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08207_ net431 net426 _04148_ vssd1 vssd1 vccd1 vccd1 _04149_ sky130_fd_sc_hd__nor3_1
XFILLER_0_91_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_43_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_43_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_170_3863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09187_ net434 net429 _04592_ net552 vssd1 vssd1 vccd1 vccd1 _05129_ sky130_fd_sc_hd__o31a_1
XFILLER_0_44_872 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_170_3874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout404_X net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11368__A1 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1146_X net1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08138_ net435 net430 vssd1 vssd1 vccd1 vccd1 _04080_ sky130_fd_sc_hd__or2_4
XANTENNA__11907__A3 net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08233__A1 net1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_79_1997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout985_A net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10040__A1 net17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11011__B net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07441__C1 net1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08069_ net729 _04008_ _04009_ net1116 vssd1 vssd1 vccd1 vccd1 _04011_ sky130_fd_sc_hd__a31o_1
X_10100_ _02831_ _02926_ _05940_ _05943_ vssd1 vssd1 vccd1 vccd1 _05944_ sky130_fd_sc_hd__o31a_1
XANTENNA__07992__B1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11080_ net832 net301 vssd1 vssd1 vccd1 vccd1 _06618_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout773_X net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10031_ team_03_WB.instance_to_wrap.BUSY_O net1040 team_03_WB.instance_to_wrap.wb.prev_BUSY_O
+ vssd1 vssd1 vccd1 vccd1 _05907_ sky130_fd_sc_hd__or3b_1
XANTENNA__13219__A net1358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11540__A1 net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07744__B1 net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08941__C1 net1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout940_X net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14770_ clknet_leaf_55_wb_clk_i _02534_ _01135_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.WRITE_I
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12096__A2 net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11982_ _06434_ net2553 net444 vssd1 vssd1 vccd1 vccd1 _01562_ sky130_fd_sc_hd__mux2_1
XFILLER_0_169_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08395__S1 net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13721_ clknet_leaf_162_wb_clk_i _01485_ _00086_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[75\]
+ sky130_fd_sc_hd__dfrtp_1
X_10933_ net503 net596 _06519_ net520 net1933 vssd1 vssd1 vccd1 vccd1 _02314_ sky130_fd_sc_hd__a32o_1
XFILLER_0_168_443 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07511__A3 net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10864_ net1252 _02808_ team_03_WB.instance_to_wrap.core.decoder.inst\[8\] vssd1
+ vssd1 vccd1 vccd1 _06463_ sky130_fd_sc_hd__or3b_4
X_13652_ clknet_leaf_133_wb_clk_i _01416_ _00017_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_156_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12603_ net1361 vssd1 vssd1 vccd1 vccd1 _00367_ sky130_fd_sc_hd__inv_2
XFILLER_0_151_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13583_ net1343 vssd1 vssd1 vccd1 vccd1 _01347_ sky130_fd_sc_hd__inv_2
XFILLER_0_137_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10795_ net685 _06398_ net585 _06402_ vssd1 vssd1 vccd1 vccd1 _06405_ sky130_fd_sc_hd__o211a_4
XANTENNA__10803__B1 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07887__A net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12534_ net1262 vssd1 vssd1 vccd1 vccd1 _00298_ sky130_fd_sc_hd__inv_2
XFILLER_0_137_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_164_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07680__C1 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12465_ net1266 vssd1 vssd1 vccd1 vccd1 _00229_ sky130_fd_sc_hd__inv_2
X_14204_ clknet_leaf_153_wb_clk_i _01968_ _00569_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[558\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08224__A1 net1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11416_ net299 net2283 net397 vssd1 vssd1 vccd1 vccd1 _02065_ sky130_fd_sc_hd__mux2_1
XANTENNA__09421__B1 team_03_WB.instance_to_wrap.core.decoder.inst\[31\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12396_ net1331 vssd1 vssd1 vccd1 vccd1 _00160_ sky130_fd_sc_hd__inv_2
XFILLER_0_104_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11347_ net276 net711 net696 vssd1 vssd1 vccd1 vccd1 _06726_ sky130_fd_sc_hd__and3_1
X_14135_ clknet_leaf_113_wb_clk_i _01899_ _00500_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[489\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10582__A2 net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11278_ net490 net621 _06706_ net408 net2160 vssd1 vssd1 vccd1 vccd1 _02156_ sky130_fd_sc_hd__a32o_1
X_14066_ clknet_leaf_117_wb_clk_i _01830_ _00431_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[420\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10760__B net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09724__A1 _04816_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10229_ team_03_WB.instance_to_wrap.core.pc.current_pc\[15\] net674 vssd1 vssd1 vccd1
+ vccd1 _06071_ sky130_fd_sc_hd__nand2_1
XANTENNA__13129__A net1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13017_ net1359 vssd1 vssd1 vccd1 vccd1 _00781_ sky130_fd_sc_hd__inv_2
XANTENNA__07735__B1 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11531__A1 net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[950\] vssd1
+ vssd1 vccd1 vccd1 net1494 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12968__A net1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_85_2113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_22_wb_clk_i_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_14968_ clknet_leaf_95_wb_clk_i _02720_ _01333_ vssd1 vssd1 vccd1 vccd1 net220 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_89 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09342__A _04207_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13919_ clknet_leaf_170_wb_clk_i _01683_ _00284_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[273\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11834__A2 net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14899_ clknet_leaf_59_wb_clk_i _02662_ _01264_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.pc.current_pc\[28\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_18_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11083__S net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07440_ _03378_ _03381_ net821 vssd1 vssd1 vccd1 vccd1 _03382_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_58_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_159_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_8_Right_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_638 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07371_ team_03_WB.instance_to_wrap.core.decoder.inst\[28\] net1019 net684 vssd1
+ vssd1 vccd1 vccd1 _03313_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_146_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_174_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09110_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[430\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[398\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[302\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[270\]
+ net976 net1075 vssd1 vssd1 vccd1 vccd1 _05052_ sky130_fd_sc_hd__mux4_1
XFILLER_0_45_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_174_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_161_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07266__A2 _03205_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08463__A1 net1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09041_ net869 _04981_ _04982_ net853 vssd1 vssd1 vccd1 vccd1 _04983_ sky130_fd_sc_hd__o211a_1
XFILLER_0_142_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_652 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08215__A1 net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold401 team_03_WB.instance_to_wrap.core.register_file.registers_state\[398\] vssd1
+ vssd1 vccd1 vccd1 net1894 sky130_fd_sc_hd__dlygate4sd3_1
Xhold412 team_03_WB.instance_to_wrap.core.register_file.registers_state\[37\] vssd1
+ vssd1 vccd1 vccd1 net1905 sky130_fd_sc_hd__dlygate4sd3_1
Xhold423 team_03_WB.instance_to_wrap.core.register_file.registers_state\[419\] vssd1
+ vssd1 vccd1 vccd1 net1916 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold434 team_03_WB.instance_to_wrap.core.register_file.registers_state\[882\] vssd1
+ vssd1 vccd1 vccd1 net1927 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold445 team_03_WB.instance_to_wrap.core.register_file.registers_state\[394\] vssd1
+ vssd1 vccd1 vccd1 net1938 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_1075 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold456 team_03_WB.instance_to_wrap.core.register_file.registers_state\[401\] vssd1
+ vssd1 vccd1 vccd1 net1949 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10573__A2 net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold467 team_03_WB.instance_to_wrap.core.register_file.registers_state\[57\] vssd1
+ vssd1 vccd1 vccd1 net1960 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11770__A1 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_129_3017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold478 team_03_WB.instance_to_wrap.core.register_file.registers_state\[279\] vssd1
+ vssd1 vccd1 vccd1 net1971 sky130_fd_sc_hd__dlygate4sd3_1
X_09943_ _04029_ net663 vssd1 vssd1 vccd1 vccd1 _05876_ sky130_fd_sc_hd__nor2_4
XTAP_TAPCELL_ROW_129_3028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold489 team_03_WB.instance_to_wrap.core.register_file.registers_state\[564\] vssd1
+ vssd1 vccd1 vccd1 net1982 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_61_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout903 net904 vssd1 vssd1 vccd1 vccd1 net903 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_111_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout914 net915 vssd1 vssd1 vccd1 vccd1 net914 sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_39_Right_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout925 net932 vssd1 vssd1 vccd1 vccd1 net925 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09715__A1 _04777_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13039__A net1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout936 net949 vssd1 vssd1 vccd1 vccd1 net936 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_74_1894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_0_wb_clk_i_X clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout399_A _06752_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09874_ _03604_ _05069_ vssd1 vssd1 vccd1 vccd1 _05816_ sky130_fd_sc_hd__nand2_1
Xfanout947 net948 vssd1 vssd1 vccd1 vccd1 net947 sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_161_wb_clk_i clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_161_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_146_3364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout958 net974 vssd1 vssd1 vccd1 vccd1 net958 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07726__B1 net1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_146_3375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout969 net974 vssd1 vssd1 vccd1 vccd1 net969 sky130_fd_sc_hd__buf_2
Xhold1101 team_03_WB.instance_to_wrap.core.register_file.registers_state\[721\] vssd1
+ vssd1 vccd1 vccd1 net2594 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1106_A net1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1112 team_03_WB.instance_to_wrap.core.register_file.registers_state\[89\] vssd1
+ vssd1 vccd1 vccd1 net2605 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1123 team_03_WB.instance_to_wrap.core.register_file.registers_state\[665\] vssd1
+ vssd1 vccd1 vccd1 net2616 sky130_fd_sc_hd__dlygate4sd3_1
X_08825_ _04765_ _04766_ net1066 vssd1 vssd1 vccd1 vccd1 _04767_ sky130_fd_sc_hd__a21o_1
Xhold1134 team_03_WB.instance_to_wrap.core.register_file.registers_state\[714\] vssd1
+ vssd1 vccd1 vccd1 net2627 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout566_A _03025_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1145 team_03_WB.instance_to_wrap.core.register_file.registers_state\[614\] vssd1
+ vssd1 vccd1 vccd1 net2638 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1156 team_03_WB.instance_to_wrap.core.register_file.registers_state\[633\] vssd1
+ vssd1 vccd1 vccd1 net2649 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1167 net180 vssd1 vssd1 vccd1 vccd1 net2660 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_135_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12078__A2 net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08756_ net1052 team_03_WB.instance_to_wrap.core.register_file.registers_state\[579\]
+ net1004 team_03_WB.instance_to_wrap.core.register_file.registers_state\[611\] net942
+ vssd1 vssd1 vccd1 vccd1 _04698_ sky130_fd_sc_hd__a221o_1
Xhold1178 team_03_WB.instance_to_wrap.core.register_file.registers_state\[653\] vssd1
+ vssd1 vccd1 vccd1 net2671 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_174_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1189 team_03_WB.instance_to_wrap.core.register_file.registers_state\[64\] vssd1
+ vssd1 vccd1 vccd1 net2682 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10089__A1 net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07707_ net1195 team_03_WB.instance_to_wrap.core.register_file.registers_state\[205\]
+ vssd1 vssd1 vccd1 vccd1 _03649_ sky130_fd_sc_hd__or2_1
XANTENNA__11286__B1 net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout733_A net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08687_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[808\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[776\]
+ net975 vssd1 vssd1 vccd1 vccd1 _04629_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout1096_X net1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08151__B1 net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_2836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_2847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07638_ net1095 team_03_WB.instance_to_wrap.core.register_file.registers_state\[462\]
+ vssd1 vssd1 vccd1 vccd1 _03580_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_48_Right_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_172_3903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_172_3914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout521_X net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout900_A net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07569_ net1201 net886 team_03_WB.instance_to_wrap.core.register_file.registers_state\[664\]
+ vssd1 vssd1 vccd1 vccd1 _03511_ sky130_fd_sc_hd__a21o_1
XFILLER_0_49_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1263_X net1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout619_X net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11721__S net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13502__A net1328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09308_ _04565_ _05248_ vssd1 vssd1 vccd1 vccd1 _05250_ sky130_fd_sc_hd__nand2_2
X_10580_ net1725 net534 net601 _05890_ vssd1 vssd1 vccd1 vccd1 _02543_ sky130_fd_sc_hd__a22o_1
XANTENNA__08454__A1 net1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10845__B _05596_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07500__A net1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09239_ _05180_ vssd1 vssd1 vccd1 vccd1 _05181_ sky130_fd_sc_hd__inv_2
XFILLER_0_51_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11022__A net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12250_ net1372 vssd1 vssd1 vccd1 vccd1 _00014_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_118_2798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout890_X net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12002__A2 _06756_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_1007 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11201_ _06413_ net2424 net487 vssd1 vssd1 vccd1 vccd1 _02207_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout988_X net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11210__A0 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12181_ net1548 vssd1 vssd1 vccd1 vccd1 _02372_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_102_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10564__A2 net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11761__A1 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_57_Right_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11132_ net640 _06641_ vssd1 vssd1 vccd1 vccd1 _06642_ sky130_fd_sc_hd__nor2_1
XANTENNA__09427__A _04476_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11676__B net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold990 team_03_WB.instance_to_wrap.core.register_file.registers_state\[578\] vssd1
+ vssd1 vccd1 vccd1 net2483 sky130_fd_sc_hd__dlygate4sd3_1
X_11063_ net832 net281 vssd1 vssd1 vccd1 vccd1 _06609_ sky130_fd_sc_hd__and2_2
XANTENNA__11395__C net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10014_ net94 net93 net96 net95 vssd1 vssd1 vccd1 vccd1 _05892_ sky130_fd_sc_hd__or4_1
XANTENNA__07193__A1 net1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07193__B2 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08390__B1 net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14822_ clknet_leaf_100_wb_clk_i net1747 _01187_ vssd1 vssd1 vccd1 vccd1 net142 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_4_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14753_ clknet_leaf_44_wb_clk_i net1810 _01118_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11816__A2 net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11965_ net632 _06742_ net464 net365 net1842 vssd1 vssd1 vccd1 vccd1 _01578_ sky130_fd_sc_hd__a32o_1
XFILLER_0_99_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_763 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_66_Right_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13704_ clknet_leaf_9_wb_clk_i _01468_ _00069_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[58\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_80_2010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10916_ net495 net596 _06505_ net518 net1977 vssd1 vssd1 vccd1 vccd1 _02317_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_80_2021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14684_ clknet_leaf_66_wb_clk_i _02448_ _01049_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.ADR_I\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08693__A1 net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_106_wb_clk_i_A clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_11896_ net633 _06705_ net466 net373 net2256 vssd1 vssd1 vccd1 vccd1 _01645_ sky130_fd_sc_hd__a32o_1
XFILLER_0_74_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13635_ net1429 vssd1 vssd1 vccd1 vccd1 _01399_ sky130_fd_sc_hd__inv_2
XFILLER_0_128_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10847_ net275 net2411 net518 vssd1 vssd1 vccd1 vccd1 _02327_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_49 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07248__A2 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08445__A1 net1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13566_ net1420 vssd1 vssd1 vccd1 vccd1 _01330_ sky130_fd_sc_hd__inv_2
X_10778_ net1251 net1252 net1018 vssd1 vssd1 vccd1 vccd1 _06388_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_27_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_4_Left_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07653__C1 net1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12517_ net1355 vssd1 vssd1 vccd1 vccd1 _00281_ sky130_fd_sc_hd__inv_2
XANTENNA__08540__S1 net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_488 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13497_ net1342 vssd1 vssd1 vccd1 vccd1 _01261_ sky130_fd_sc_hd__inv_2
XFILLER_0_140_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12448_ net1400 vssd1 vssd1 vccd1 vccd1 _00212_ sky130_fd_sc_hd__inv_2
XANTENNA__11289__D net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_75_Right_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11201__A0 _06413_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_352 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07405__C1 net1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12379_ net1362 vssd1 vssd1 vccd1 vccd1 _00143_ sky130_fd_sc_hd__inv_2
XFILLER_0_22_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07409__X _03351_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14118_ clknet_leaf_28_wb_clk_i _01882_ _00483_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[472\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15098_ net912 vssd1 vssd1 vccd1 vccd1 net258 sky130_fd_sc_hd__clkbuf_1
X_06940_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[804\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[772\]
+ net776 vssd1 vssd1 vccd1 vccd1 _02882_ sky130_fd_sc_hd__mux2_1
X_14049_ clknet_leaf_177_wb_clk_i _01813_ _00414_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[403\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_157_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07708__B1 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_52_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06871_ team_03_WB.instance_to_wrap.core.control_logic.instruction\[3\] team_03_WB.instance_to_wrap.core.control_logic.instruction\[2\]
+ team_03_WB.instance_to_wrap.core.control_logic.instruction\[1\] team_03_WB.instance_to_wrap.core.control_logic.instruction\[0\]
+ vssd1 vssd1 vccd1 vccd1 _02813_ sky130_fd_sc_hd__nand4_4
XFILLER_0_94_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_145_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_59_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_4_4__f_wb_clk_i_A clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11806__S net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08610_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[37\] net992
+ vssd1 vssd1 vccd1 vccd1 _04552_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_2_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09590_ _05420_ _05525_ net568 vssd1 vssd1 vccd1 vccd1 _05532_ sky130_fd_sc_hd__mux2_1
XFILLER_0_173_23 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_84_Right_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_141_3261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_141_3272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08541_ net1220 _04482_ _04481_ vssd1 vssd1 vccd1 vccd1 _04483_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_77_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11268__B1 net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11107__A net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_251 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08472_ _04408_ _04413_ net871 vssd1 vssd1 vccd1 vccd1 _04414_ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09800__A net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07423_ net1176 team_03_WB.instance_to_wrap.core.register_file.registers_state\[980\]
+ vssd1 vssd1 vccd1 vccd1 _03365_ sky130_fd_sc_hd__or2_1
XFILLER_0_9_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_159_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07023__C net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07354_ _03294_ _03295_ net817 vssd1 vssd1 vccd1 vccd1 _03296_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_162_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07285_ net1202 team_03_WB.instance_to_wrap.core.register_file.registers_state\[169\]
+ vssd1 vssd1 vccd1 vccd1 _03227_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout314_A _05387_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_488 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_91 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1056_A net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09024_ net1244 team_03_WB.instance_to_wrap.core.register_file.registers_state\[464\]
+ net989 team_03_WB.instance_to_wrap.core.register_file.registers_state\[496\] net1216
+ vssd1 vssd1 vccd1 vccd1 _04966_ sky130_fd_sc_hd__o221a_1
XPHY_EDGE_ROW_93_Right_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09946__S net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_574 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_1934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold220 team_03_WB.instance_to_wrap.CPU_DAT_I\[4\] vssd1 vssd1 vccd1 vccd1 net1713
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_1945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10681__A net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold231 team_03_WB.instance_to_wrap.core.register_file.registers_state\[314\] vssd1
+ vssd1 vccd1 vccd1 net1724 sky130_fd_sc_hd__dlygate4sd3_1
Xhold242 team_03_WB.instance_to_wrap.CPU_DAT_I\[22\] vssd1 vssd1 vccd1 vccd1 net1735
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_148_3404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1223_A net1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_184_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_148_3415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold253 team_03_WB.instance_to_wrap.CPU_DAT_I\[15\] vssd1 vssd1 vccd1 vccd1 net1746
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09247__A _03428_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_379 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold264 team_03_WB.instance_to_wrap.core.register_file.registers_state\[306\] vssd1
+ vssd1 vccd1 vccd1 net1757 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_113_2695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold275 team_03_WB.instance_to_wrap.core.register_file.registers_state\[686\] vssd1
+ vssd1 vccd1 vccd1 net1768 sky130_fd_sc_hd__dlygate4sd3_1
Xhold286 team_03_WB.instance_to_wrap.CPU_DAT_I\[18\] vssd1 vssd1 vccd1 vccd1 net1779
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout683_A _05915_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout700 _06561_ vssd1 vssd1 vccd1 vccd1 net700 sky130_fd_sc_hd__clkbuf_4
Xhold297 net184 vssd1 vssd1 vccd1 vccd1 net1790 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout711 net716 vssd1 vssd1 vccd1 vccd1 net711 sky130_fd_sc_hd__buf_4
X_09926_ _05861_ net2011 net292 vssd1 vssd1 vccd1 vccd1 _02764_ sky130_fd_sc_hd__mux2_1
Xfanout722 _02863_ vssd1 vssd1 vccd1 vccd1 net722 sky130_fd_sc_hd__buf_4
XFILLER_0_102_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_165_3762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1011_X net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout733 net738 vssd1 vssd1 vccd1 vccd1 net733 sky130_fd_sc_hd__buf_2
Xfanout744 net745 vssd1 vssd1 vccd1 vccd1 net744 sky130_fd_sc_hd__buf_2
Xfanout755 _02852_ vssd1 vssd1 vccd1 vccd1 net755 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout1109_X net1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout766 net770 vssd1 vssd1 vccd1 vccd1 net766 sky130_fd_sc_hd__clkbuf_4
X_09857_ _05784_ _05798_ vssd1 vssd1 vccd1 vccd1 _05799_ sky130_fd_sc_hd__or2_2
XANTENNA_fanout850_A _04096_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout777 _02851_ vssd1 vssd1 vccd1 vccd1 net777 sky130_fd_sc_hd__buf_2
XANTENNA__07175__A1 net1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout471_X net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout788 net789 vssd1 vssd1 vccd1 vccd1 net788 sky130_fd_sc_hd__buf_4
XANTENNA_fanout569_X net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout948_A net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout799 net800 vssd1 vssd1 vccd1 vccd1 net799 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08372__B1 net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15093__1479 vssd1 vssd1 vccd1 vccd1 _15093__1479/HI net1479 sky130_fd_sc_hd__conb_1
XANTENNA__11716__S net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08808_ net1052 team_03_WB.instance_to_wrap.core.register_file.registers_state\[449\]
+ net1005 team_03_WB.instance_to_wrap.core.register_file.registers_state\[481\] net1076
+ vssd1 vssd1 vccd1 vccd1 _04750_ sky130_fd_sc_hd__a221o_1
X_09788_ net582 _05720_ _05729_ vssd1 vssd1 vccd1 vccd1 _05730_ sky130_fd_sc_hd__a21oi_4
XANTENNA__12401__A net1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08739_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[35\] net980
+ vssd1 vssd1 vccd1 vccd1 _04681_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout1380_X net1380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08124__B1 net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout736_X net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11017__A net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07478__A2 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11750_ _06573_ net478 net334 net2013 vssd1 vssd1 vccd1 vccd1 _01787_ sky130_fd_sc_hd__a22o_1
XFILLER_0_138_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_355 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_744 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10701_ _06316_ _06338_ net606 vssd1 vssd1 vccd1 vccd1 _06339_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout903_X net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11681_ _06723_ net385 net339 net1984 vssd1 vssd1 vccd1 vccd1 _01853_ sky130_fd_sc_hd__a22o_1
XFILLER_0_138_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13420_ net1427 vssd1 vssd1 vccd1 vccd1 _01184_ sky130_fd_sc_hd__inv_2
XFILLER_0_138_479 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13232__A net1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10632_ team_03_WB.instance_to_wrap.core.decoder.inst\[29\] net1808 net845 vssd1
+ vssd1 vccd1 vccd1 _02496_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08427__A1 net1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07230__A net1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11431__A0 net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10563_ net1997 net531 net598 _05873_ vssd1 vssd1 vccd1 vccd1 _02560_ sky130_fd_sc_hd__a22o_1
X_13351_ net1318 vssd1 vssd1 vccd1 vccd1 _01115_ sky130_fd_sc_hd__inv_2
Xmax_cap1017 _02817_ vssd1 vssd1 vccd1 vccd1 net1017 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_10_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12302_ net1274 vssd1 vssd1 vccd1 vccd1 _00066_ sky130_fd_sc_hd__inv_2
XFILLER_0_106_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10494_ net106 net1029 net907 net1526 vssd1 vssd1 vccd1 vccd1 _02615_ sky130_fd_sc_hd__a22o_1
X_13282_ net1404 vssd1 vssd1 vccd1 vccd1 _01046_ sky130_fd_sc_hd__inv_2
XANTENNA_input77_A wbs_adr_i[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07650__A2 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15021_ clknet_leaf_100_wb_clk_i _02741_ _01386_ vssd1 vssd1 vccd1 vccd1 net177 sky130_fd_sc_hd__dfrtp_1
X_12233_ net1694 vssd1 vssd1 vccd1 vccd1 _01424_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__08286__S0 net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11734__A1 net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10537__A2 net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12164_ net1559 vssd1 vssd1 vccd1 vccd1 _02389_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_9_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11115_ net263 net2564 net418 vssd1 vssd1 vccd1 vccd1 _02244_ sky130_fd_sc_hd__mux2_1
X_12095_ net620 _06666_ net453 net439 net2111 vssd1 vssd1 vccd1 vccd1 _01452_ sky130_fd_sc_hd__a32o_1
XANTENNA__09591__S net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11498__A0 _06619_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_16 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11046_ net702 net715 net295 vssd1 vssd1 vccd1 vccd1 _06600_ sky130_fd_sc_hd__or3b_1
XANTENNA__07166__A1 team_03_WB.instance_to_wrap.core.decoder.inst\[19\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08363__B1 net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14805_ clknet_leaf_88_wb_clk_i _02569_ _01170_ vssd1 vssd1 vccd1 vccd1 net173 sky130_fd_sc_hd__dfrtp_1
X_12997_ net1354 vssd1 vssd1 vccd1 vccd1 _00761_ sky130_fd_sc_hd__inv_2
XANTENNA__11572__D net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_157_700 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07124__B _03065_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14736_ clknet_leaf_32_wb_clk_i _02500_ _01101_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_169_571 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11948_ net644 _06725_ net478 net366 net1908 vssd1 vssd1 vccd1 vccd1 _01595_ sky130_fd_sc_hd__a32o_1
XANTENNA__08666__A1 net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09863__B1 net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14667_ clknet_leaf_45_wb_clk_i _02431_ _01032_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1021\]
+ sky130_fd_sc_hd__dfstp_1
X_11879_ net619 _06688_ net452 net371 net1909 vssd1 vssd1 vccd1 vccd1 _01662_ sky130_fd_sc_hd__a32o_1
XFILLER_0_7_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_156_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13618_ net1422 vssd1 vssd1 vccd1 vccd1 _01382_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08418__A1 net1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14598_ clknet_leaf_69_wb_clk_i _02362_ _00963_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[952\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_28_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07140__A net1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13549_ net1321 vssd1 vssd1 vccd1 vccd1 _01313_ sky130_fd_sc_hd__inv_2
XFILLER_0_125_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09091__A1 net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11973__A1 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_2370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_814 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07070_ net1105 team_03_WB.instance_to_wrap.core.register_file.registers_state\[66\]
+ net797 team_03_WB.instance_to_wrap.core.register_file.registers_state\[98\] net746
+ vssd1 vssd1 vccd1 vccd1 _03012_ sky130_fd_sc_hd__a221o_1
XANTENNA__08670__S net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_93_2278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10528__A2 net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11725__A1 net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_2289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_390 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_1831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07972_ net813 _03909_ _03910_ _03913_ vssd1 vssd1 vccd1 vccd1 _03914_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_71_1842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_3312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09711_ _03682_ net536 _05041_ _03679_ _02804_ vssd1 vssd1 vccd1 vccd1 _05653_ sky130_fd_sc_hd__o32a_1
X_06923_ net1200 team_03_WB.instance_to_wrap.core.register_file.registers_state\[356\]
+ net886 vssd1 vssd1 vccd1 vccd1 _02865_ sky130_fd_sc_hd__and3_1
XANTENNA__07157__A1 net1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13317__A net1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09642_ _05185_ _05192_ _05501_ vssd1 vssd1 vccd1 vccd1 _05584_ sky130_fd_sc_hd__and3_1
XFILLER_0_93_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06854_ net1 vssd1 vssd1 vccd1 vccd1 _02797_ sky130_fd_sc_hd__inv_2
XANTENNA__10161__B1 _03679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_160_3670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09573_ net321 _05354_ _05384_ _05513_ _05512_ vssd1 vssd1 vccd1 vccd1 _05515_ sky130_fd_sc_hd__a221o_1
XFILLER_0_171_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_171 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1130 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08524_ net1227 team_03_WB.instance_to_wrap.core.register_file.registers_state\[223\]
+ net952 team_03_WB.instance_to_wrap.core.register_file.registers_state\[255\] net934
+ vssd1 vssd1 vccd1 vccd1 _04466_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_69_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10464__A1 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08455_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[828\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[796\]
+ net953 vssd1 vssd1 vccd1 vccd1 _04397_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1173_A net1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout529_A _06309_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13052__A net1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07406_ net1171 team_03_WB.instance_to_wrap.core.register_file.registers_state\[735\]
+ net758 team_03_WB.instance_to_wrap.core.register_file.registers_state\[767\] net1149
+ vssd1 vssd1 vccd1 vccd1 _03348_ sky130_fd_sc_hd__o221a_1
XFILLER_0_163_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08386_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[57\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[25\]
+ net992 vssd1 vssd1 vccd1 vccd1 _04328_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07880__A2 net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07337_ team_03_WB.instance_to_wrap.core.decoder.inst\[29\] net1019 net684 vssd1
+ vssd1 vccd1 vccd1 _03279_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_135_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1340_A net1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout317_X net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11964__A1 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1059_X net1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07985__A net1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07268_ net1202 team_03_WB.instance_to_wrap.core.register_file.registers_state\[841\]
+ vssd1 vssd1 vccd1 vccd1 _03210_ sky130_fd_sc_hd__or2_1
XFILLER_0_104_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_115_2735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11003__C net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_767 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_2746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout898_A net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09007_ _04945_ _04946_ net854 vssd1 vssd1 vccd1 vccd1 _04949_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_14_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_167_3802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10615__S net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07199_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[178\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[146\]
+ net756 vssd1 vssd1 vccd1 vccd1 _03141_ sky130_fd_sc_hd__mux2_1
XANTENNA__10519__A2 net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_167_3813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1226_X net1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11716__A1 net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout530 _06309_ vssd1 vssd1 vccd1 vccd1 net530 sky130_fd_sc_hd__clkbuf_2
Xfanout541 net542 vssd1 vssd1 vccd1 vccd1 net541 sky130_fd_sc_hd__buf_2
XANTENNA__09705__A _05646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09909_ _05454_ _05563_ _05848_ _05850_ vssd1 vssd1 vccd1 vccd1 _05851_ sky130_fd_sc_hd__or4_1
Xfanout552 _03105_ vssd1 vssd1 vccd1 vccd1 net552 sky130_fd_sc_hd__buf_2
Xfanout563 net564 vssd1 vssd1 vccd1 vccd1 net563 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09910__C_N _05429_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout574 net577 vssd1 vssd1 vccd1 vccd1 net574 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout853_X net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07148__A1 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout585 net586 vssd1 vssd1 vccd1 vccd1 net585 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10350__S net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12920_ net1376 vssd1 vssd1 vccd1 vccd1 _00684_ sky130_fd_sc_hd__inv_2
Xfanout596 net597 vssd1 vssd1 vccd1 vccd1 net596 sky130_fd_sc_hd__buf_4
XFILLER_0_77_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12851_ net1265 vssd1 vssd1 vccd1 vccd1 _00615_ sky130_fd_sc_hd__inv_2
Xclkbuf_4_9__f_wb_clk_i clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_9__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_69_812 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11802_ net2453 net265 net329 vssd1 vssd1 vccd1 vccd1 _01736_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_4_3__f_wb_clk_i_X clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_12782_ net1310 vssd1 vssd1 vccd1 vccd1 _00546_ sky130_fd_sc_hd__inv_2
XFILLER_0_150_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_815 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14521_ clknet_leaf_155_wb_clk_i _02285_ _00886_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[875\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07856__C1 net1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11733_ net1874 net296 net337 vssd1 vssd1 vccd1 vccd1 _01803_ sky130_fd_sc_hd__mux2_1
XFILLER_0_166_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14452_ clknet_leaf_134_wb_clk_i _02216_ _00817_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[806\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_25_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11664_ net2269 _06505_ net344 vssd1 vssd1 vccd1 vccd1 _01869_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08056__A net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11404__A0 net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13403_ net1432 vssd1 vssd1 vccd1 vccd1 _01167_ sky130_fd_sc_hd__inv_2
XFILLER_0_52_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10615_ net1551 team_03_WB.instance_to_wrap.CPU_DAT_O\[14\] net842 vssd1 vssd1 vccd1
+ vccd1 _02513_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07608__C1 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14383_ clknet_leaf_136_wb_clk_i _02147_ _00748_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[737\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11595_ net297 net2368 net449 vssd1 vssd1 vccd1 vccd1 _01934_ sky130_fd_sc_hd__mux2_1
XANTENNA__10758__A2 net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11955__A1 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_148_1068 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13334_ net1325 vssd1 vssd1 vccd1 vccd1 _01098_ sky130_fd_sc_hd__inv_2
X_10546_ _06289_ vssd1 vssd1 vccd1 vccd1 _06290_ sky130_fd_sc_hd__inv_2
XFILLER_0_150_964 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13265_ net1269 vssd1 vssd1 vccd1 vccd1 _01029_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_94_Left_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10477_ net124 net1027 net905 net1699 vssd1 vssd1 vccd1 vccd1 _02632_ sky130_fd_sc_hd__a22o_1
X_15004_ clknet_leaf_59_wb_clk_i net52 _01369_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_150_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_839 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12216_ net1651 vssd1 vssd1 vccd1 vccd1 _01441_ sky130_fd_sc_hd__clkbuf_1
X_13196_ net1314 vssd1 vssd1 vccd1 vccd1 _00960_ sky130_fd_sc_hd__inv_2
XANTENNA__11567__D net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11183__A2 net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07119__B _03060_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12147_ net1558 vssd1 vssd1 vccd1 vccd1 _02406_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__10391__B1 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12078_ _06783_ net475 net441 net1839 vssd1 vssd1 vccd1 vccd1 _01469_ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_1051 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11029_ net701 net712 _06495_ vssd1 vssd1 vccd1 vccd1 _06589_ sky130_fd_sc_hd__or3b_1
XFILLER_0_2_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_154_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07135__A net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_300 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11891__B1 net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09621__Y _05563_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08639__A1 net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08665__S net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_47_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09300__A2 _05144_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14719_ clknet_leaf_44_wb_clk_i _02483_ _01084_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.decoder.inst\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07311__A1 net1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08240_ net1226 team_03_WB.instance_to_wrap.core.register_file.registers_state\[178\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[146\] net950 net916
+ vssd1 vssd1 vccd1 vccd1 _04182_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_99_2410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_3160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08171_ net1230 team_03_WB.instance_to_wrap.core.register_file.registers_state\[980\]
+ net958 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1012\] net1217
+ vssd1 vssd1 vccd1 vccd1 _04113_ sky130_fd_sc_hd__o221a_1
XANTENNA__11104__B net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09064__A1 net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_136_3171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08498__S0 net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_146 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_2318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11946__A1 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_2329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07122_ net614 _03059_ _03061_ vssd1 vssd1 vccd1 vccd1 _03064_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_43_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15092__1478 vssd1 vssd1 vccd1 vccd1 _15092__1478/HI net1478 sky130_fd_sc_hd__conb_1
XFILLER_0_127_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08811__A1 net1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10943__B _06527_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10084__A_N _05082_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_3079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07053_ net614 _02994_ vssd1 vssd1 vccd1 vccd1 _02995_ sky130_fd_sc_hd__nor2_1
XFILLER_0_113_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_864 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07090__A3 net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput111 net111 vssd1 vssd1 vccd1 vccd1 ADR_O[17] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_112_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput122 net122 vssd1 vssd1 vccd1 vccd1 ADR_O[27] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_11_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput133 net133 vssd1 vssd1 vccd1 vccd1 ADR_O[8] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_2_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08024__C1 net1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput144 net144 vssd1 vssd1 vccd1 vccd1 DAT_O[17] sky130_fd_sc_hd__buf_2
XFILLER_0_11_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput155 net155 vssd1 vssd1 vccd1 vccd1 DAT_O[27] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_110_2632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07378__A1 net1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11477__D net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_2643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput166 net166 vssd1 vssd1 vccd1 vccd1 DAT_O[8] sky130_fd_sc_hd__buf_2
XANTENNA__11174__A2 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput177 net177 vssd1 vssd1 vccd1 vccd1 gpio_oeb[12] sky130_fd_sc_hd__buf_2
Xoutput188 net188 vssd1 vssd1 vccd1 vccd1 gpio_oeb[23] sky130_fd_sc_hd__buf_2
Xoutput199 net199 vssd1 vssd1 vccd1 vccd1 gpio_oeb[34] sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_162_3710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1019_A net1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_68_wb_clk_i clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_68_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_07955_ net1128 _03896_ _03895_ net1138 vssd1 vssd1 vccd1 vccd1 _03897_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout381_A net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout479_A net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13047__A net1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06906_ net1116 net895 vssd1 vssd1 vccd1 vccd1 _02848_ sky130_fd_sc_hd__nor2_1
X_07886_ net729 _03824_ _03825_ _03826_ _03827_ vssd1 vssd1 vccd1 vccd1 _03828_ sky130_fd_sc_hd__a32o_1
X_09625_ net565 net556 _05137_ vssd1 vssd1 vccd1 vccd1 _05567_ sky130_fd_sc_hd__and3_1
X_06837_ team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[11\] vssd1 vssd1 vccd1
+ vccd1 _02780_ sky130_fd_sc_hd__inv_2
XFILLER_0_69_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11882__B1 net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_2594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout646_A net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout267_X net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1290_A net1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09556_ _05371_ _05485_ _05497_ vssd1 vssd1 vccd1 vccd1 _05498_ sky130_fd_sc_hd__a21oi_2
XANTENNA__06884__A team_03_WB.instance_to_wrap.core.decoder.inst\[30\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10437__A1 _06057_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09260__A net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08507_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[575\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[543\]
+ net959 vssd1 vssd1 vccd1 vccd1 _04449_ sky130_fd_sc_hd__mux2_1
XANTENNA__11634__B1 net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09487_ _05389_ _05390_ _05428_ vssd1 vssd1 vccd1 vccd1 _05429_ sky130_fd_sc_hd__a21o_2
XANTENNA_fanout813_A net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10988__A2 net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1176_X net1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07051__Y _02993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08438_ _04376_ _04377_ _04379_ _04378_ net937 net861 vssd1 vssd1 vccd1 vccd1 _04380_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_156_3569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_22_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09055__A1 net1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout601_X net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08369_ net1236 team_03_WB.instance_to_wrap.core.register_file.registers_state\[726\]
+ net971 team_03_WB.instance_to_wrap.core.register_file.registers_state\[758\] net939
+ vssd1 vssd1 vccd1 vccd1 _04311_ sky130_fd_sc_hd__o221a_1
XFILLER_0_117_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10400_ _06076_ _06225_ vssd1 vssd1 vccd1 vccd1 _06226_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_150_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_460 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07066__B1 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11380_ net503 net632 _06742_ net402 net1787 vssd1 vssd1 vccd1 vccd1 _02090_ sky130_fd_sc_hd__a32o_1
XFILLER_0_150_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10331_ team_03_WB.instance_to_wrap.core.pc.current_pc\[27\] _06150_ vssd1 vssd1
+ vccd1 vccd1 _06169_ sky130_fd_sc_hd__nor2_1
XANTENNA__11030__A net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10262_ _05981_ _06091_ vssd1 vssd1 vccd1 vccd1 _06104_ sky130_fd_sc_hd__nand2_1
X_13050_ net1372 vssd1 vssd1 vccd1 vccd1 _00814_ sky130_fd_sc_hd__inv_2
XFILLER_0_104_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout970_X net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07369__A1 net1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11387__D net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12001_ net269 net2629 net445 vssd1 vssd1 vccd1 vccd1 _01543_ sky130_fd_sc_hd__mux2_1
X_10193_ _06033_ _06034_ _02893_ vssd1 vssd1 vccd1 vccd1 _06035_ sky130_fd_sc_hd__a21oi_1
Xfanout1303 net1305 vssd1 vssd1 vccd1 vccd1 net1303 sky130_fd_sc_hd__buf_4
Xfanout1314 net1315 vssd1 vssd1 vccd1 vccd1 net1314 sky130_fd_sc_hd__buf_4
Xfanout1325 net1326 vssd1 vssd1 vccd1 vccd1 net1325 sky130_fd_sc_hd__buf_4
XFILLER_0_79_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1336 net1338 vssd1 vssd1 vccd1 vccd1 net1336 sky130_fd_sc_hd__buf_4
Xfanout1347 net1349 vssd1 vssd1 vccd1 vccd1 net1347 sky130_fd_sc_hd__buf_4
XANTENNA__08318__B1 net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1358 net1437 vssd1 vssd1 vccd1 vccd1 net1358 sky130_fd_sc_hd__clkbuf_4
Xfanout360 _06817_ vssd1 vssd1 vccd1 vccd1 net360 sky130_fd_sc_hd__buf_4
XFILLER_0_108_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout371 _06813_ vssd1 vssd1 vccd1 vccd1 net371 sky130_fd_sc_hd__buf_6
Xfanout1369 net1370 vssd1 vssd1 vccd1 vccd1 net1369 sky130_fd_sc_hd__buf_4
XFILLER_0_17_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout382 net387 vssd1 vssd1 vccd1 vccd1 net382 sky130_fd_sc_hd__clkbuf_4
X_13952_ clknet_leaf_2_wb_clk_i _01716_ _00317_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[306\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout393 net395 vssd1 vssd1 vccd1 vccd1 net393 sky130_fd_sc_hd__buf_6
XANTENNA__11873__A0 net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12903_ net1363 vssd1 vssd1 vccd1 vccd1 _00667_ sky130_fd_sc_hd__inv_2
X_13883_ clknet_leaf_134_wb_clk_i _01647_ _00248_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[237\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07541__A1 net1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12834_ net1350 vssd1 vssd1 vccd1 vccd1 _00598_ sky130_fd_sc_hd__inv_2
XANTENNA__09818__B1 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08485__S net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_973 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_338 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10428__A1 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11625__B1 net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12765_ net1384 vssd1 vssd1 vccd1 vccd1 _00529_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14504_ clknet_leaf_10_wb_clk_i _02268_ _00869_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[858\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_166_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11716_ net1897 net278 net335 vssd1 vssd1 vccd1 vccd1 _01820_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_166_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12696_ net1379 vssd1 vssd1 vccd1 vccd1 _00460_ sky130_fd_sc_hd__inv_2
XFILLER_0_44_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_140_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14435_ clknet_leaf_33_wb_clk_i _02199_ _00800_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[789\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_42_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11647_ net2763 _06613_ net342 vssd1 vssd1 vccd1 vccd1 _01886_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_42_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09046__A1 net1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput13 DAT_I[1] vssd1 vssd1 vccd1 vccd1 net13 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__12050__A0 _06619_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_739 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput24 DAT_I[2] vssd1 vssd1 vccd1 vccd1 net24 sky130_fd_sc_hd__buf_1
XFILLER_0_3_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput35 gpio_in[10] vssd1 vssd1 vccd1 vccd1 net35 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14366_ clknet_leaf_119_wb_clk_i _02130_ _00731_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[720\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput46 gpio_in[21] vssd1 vssd1 vccd1 vccd1 net46 sky130_fd_sc_hd__clkbuf_1
X_11578_ _06413_ net2705 net448 vssd1 vssd1 vccd1 vccd1 _01951_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10763__B net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput57 gpio_in[32] vssd1 vssd1 vccd1 vccd1 net57 sky130_fd_sc_hd__clkbuf_1
Xinput68 wbs_adr_i[10] vssd1 vssd1 vccd1 vccd1 net68 sky130_fd_sc_hd__clkbuf_1
X_13317_ net1326 vssd1 vssd1 vccd1 vccd1 _01081_ sky130_fd_sc_hd__inv_2
Xhold808 team_03_WB.instance_to_wrap.core.register_file.registers_state\[620\] vssd1
+ vssd1 vccd1 vccd1 net2301 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10529_ net137 net1031 net1023 net1782 vssd1 vssd1 vccd1 vccd1 _02581_ sky130_fd_sc_hd__a22o_1
Xinput79 wbs_adr_i[20] vssd1 vssd1 vccd1 vccd1 net79 sky130_fd_sc_hd__buf_1
Xhold819 team_03_WB.instance_to_wrap.core.register_file.registers_state\[511\] vssd1
+ vssd1 vccd1 vccd1 net2312 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_172_Right_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14297_ clknet_leaf_168_wb_clk_i _02061_ _00662_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[651\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_90_2215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_2226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13248_ net1403 vssd1 vssd1 vccd1 vccd1 _01012_ sky130_fd_sc_hd__inv_2
XFILLER_0_161_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_973 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11156__A2 net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08557__B1 net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11875__A net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13179_ net1365 vssd1 vssd1 vccd1 vccd1 _00943_ sky130_fd_sc_hd__inv_2
XANTENNA__08021__A2 net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07765__D1 net1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11086__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07740_ _03680_ _03681_ vssd1 vssd1 vccd1 vccd1 _03682_ sky130_fd_sc_hd__or2_1
XANTENNA__07207__S1 net1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_88_2177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_2188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07671_ net742 _03611_ _03612_ net806 vssd1 vssd1 vccd1 vccd1 _03613_ sky130_fd_sc_hd__a31o_1
X_09410_ net543 net354 _04209_ vssd1 vssd1 vccd1 vccd1 _05352_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_133_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09809__B1 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10419__B2 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_3200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09341_ _04207_ _05282_ vssd1 vssd1 vccd1 vccd1 _05283_ sky130_fd_sc_hd__nor2_1
XANTENNA__11616__B1 net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08088__A2 net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_3211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_186_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_186_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_90_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_103_2491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07296__B1 net1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09272_ _03244_ _05145_ net609 vssd1 vssd1 vccd1 vccd1 _05214_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_62_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08493__C1 net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_115_wb_clk_i clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_115_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_30_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_157_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_134_3119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08223_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[945\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[913\]
+ net962 vssd1 vssd1 vccd1 vccd1 _04165_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_706 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10954__A net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09588__A2 _04382_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08154_ team_03_WB.instance_to_wrap.core.decoder.inst\[19\] _02820_ vssd1 vssd1 vccd1
+ vccd1 _04096_ sky130_fd_sc_hd__and2_4
XTAP_TAPCELL_ROW_151_3466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08424__A net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_151_3477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07105_ net1199 team_03_WB.instance_to_wrap.core.register_file.registers_state\[481\]
+ net883 _03045_ net1134 vssd1 vssd1 vccd1 vccd1 _03047_ sky130_fd_sc_hd__a311o_1
XFILLER_0_113_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08085_ net1141 _04022_ _04024_ _04026_ net721 vssd1 vssd1 vccd1 vccd1 _04027_ sky130_fd_sc_hd__o41a_1
XANTENNA__11488__C net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1136_A net1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09954__S net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07036_ _02975_ _02977_ net809 vssd1 vssd1 vccd1 vccd1 _02978_ sky130_fd_sc_hd__o21a_1
XANTENNA__11147__A2 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout596_A net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08548__B1 net1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1303_A net1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07220__B1 net1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout763_A net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08987_ net1046 team_03_WB.instance_to_wrap.core.register_file.registers_state\[202\]
+ net996 team_03_WB.instance_to_wrap.core.register_file.registers_state\[234\] net918
+ vssd1 vssd1 vccd1 vccd1 _04929_ sky130_fd_sc_hd__a221o_1
XANTENNA__07771__A1 net1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout384_X net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07938_ net1162 _03879_ vssd1 vssd1 vccd1 vccd1 _03880_ sky130_fd_sc_hd__nor2_1
XANTENNA__10658__A1 team_03_WB.instance_to_wrap.CPU_DAT_O\[3\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11855__A0 _06468_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_2981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout930_A net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07869_ net1120 _03809_ _03810_ vssd1 vssd1 vccd1 vccd1 _03811_ sky130_fd_sc_hd__nor3_1
XANTENNA_fanout649_X net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11724__S net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09608_ _05464_ _05470_ net569 vssd1 vssd1 vccd1 vccd1 _05550_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_27_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_158_3609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10880_ net314 net309 _05928_ team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[17\]
+ vssd1 vssd1 vccd1 vccd1 _06476_ sky130_fd_sc_hd__or4b_2
XFILLER_0_78_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11607__A0 _06557_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09539_ net580 _04824_ _05125_ vssd1 vssd1 vccd1 vccd1 _05481_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout816_X net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_159_Left_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11025__A net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07287__B1 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12550_ net1300 vssd1 vssd1 vccd1 vccd1 _00314_ sky130_fd_sc_hd__inv_2
XFILLER_0_93_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11501_ _06469_ net2721 net388 vssd1 vssd1 vccd1 vccd1 _02005_ sky130_fd_sc_hd__mux2_1
X_12481_ net1282 vssd1 vssd1 vccd1 vccd1 _00245_ sky130_fd_sc_hd__inv_2
XFILLER_0_163_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13240__A net1380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14220_ clknet_leaf_18_wb_clk_i _01984_ _00585_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[574\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09123__S1 net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11432_ net506 net263 _06756_ net398 net2185 vssd1 vssd1 vccd1 vccd1 _02052_ sky130_fd_sc_hd__a32o_1
XFILLER_0_80_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12032__B1 net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_238 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07134__S0 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11386__A2 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08787__B1 net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14151_ clknet_leaf_113_wb_clk_i _01915_ _00516_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[505\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11363_ net714 net272 net699 vssd1 vssd1 vccd1 vccd1 _06734_ sky130_fd_sc_hd__and3_1
XFILLER_0_21_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13102_ net1303 vssd1 vssd1 vccd1 vccd1 _00866_ sky130_fd_sc_hd__inv_2
X_10314_ _02766_ net677 _06133_ _06155_ vssd1 vssd1 vccd1 vccd1 _02665_ sky130_fd_sc_hd__a2bb2o_1
X_14082_ clknet_leaf_173_wb_clk_i _01846_ _00447_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[436\]
+ sky130_fd_sc_hd__dfrtp_1
X_11294_ net505 net633 _06714_ net410 net2167 vssd1 vssd1 vccd1 vccd1 _02148_ sky130_fd_sc_hd__a32o_1
XPHY_EDGE_ROW_168_Left_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13033_ net1256 vssd1 vssd1 vccd1 vccd1 _00797_ sky130_fd_sc_hd__inv_2
X_10245_ _05991_ _06086_ vssd1 vssd1 vccd1 vccd1 _06087_ sky130_fd_sc_hd__nor2_1
XANTENNA__09200__A1 _02954_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08634__S0 net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1100 net1101 vssd1 vssd1 vccd1 vccd1 net1100 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_119_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1111 net1113 vssd1 vssd1 vccd1 vccd1 net1111 sky130_fd_sc_hd__buf_2
X_10176_ team_03_WB.instance_to_wrap.core.pc.current_pc\[9\] net675 vssd1 vssd1 vccd1
+ vccd1 _06018_ sky130_fd_sc_hd__nand2_1
Xfanout1122 _02786_ vssd1 vssd1 vccd1 vccd1 net1122 sky130_fd_sc_hd__buf_4
Xfanout1133 net1134 vssd1 vssd1 vccd1 vccd1 net1133 sky130_fd_sc_hd__buf_4
Xfanout1144 team_03_WB.EN_VAL_REG vssd1 vssd1 vccd1 vccd1 net1144 sky130_fd_sc_hd__clkbuf_4
Xfanout1155 net1157 vssd1 vssd1 vccd1 vccd1 net1155 sky130_fd_sc_hd__buf_4
XANTENNA__12099__B1 net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1166 net1168 vssd1 vssd1 vccd1 vccd1 net1166 sky130_fd_sc_hd__clkbuf_4
X_14984_ clknet_leaf_81_wb_clk_i net63 _01349_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_156_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1177 net1178 vssd1 vssd1 vccd1 vccd1 net1177 sky130_fd_sc_hd__buf_2
XANTENNA_clkbuf_leaf_12_wb_clk_i_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout1188 net1189 vssd1 vssd1 vccd1 vccd1 net1188 sky130_fd_sc_hd__buf_2
XFILLER_0_156_1134 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1199 net1206 vssd1 vssd1 vccd1 vccd1 net1199 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11846__A0 net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13935_ clknet_leaf_143_wb_clk_i _01699_ _00300_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[289\]
+ sky130_fd_sc_hd__dfrtp_1
X_15091__1477 vssd1 vssd1 vccd1 vccd1 _15091__1477/HI net1477 sky130_fd_sc_hd__conb_1
XANTENNA__08711__B1 net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07514__B2 net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload5_A clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13866_ clknet_leaf_0_wb_clk_i _01630_ _00231_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[220\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_159_658 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12817_ net1274 vssd1 vssd1 vccd1 vccd1 _00581_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_83_2074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13797_ clknet_leaf_12_wb_clk_i _01561_ _00162_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[151\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_173_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_511 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_807 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12748_ net1312 vssd1 vssd1 vccd1 vccd1 _00512_ sky130_fd_sc_hd__inv_2
XFILLER_0_17_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_987 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_330 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12679_ net1368 vssd1 vssd1 vccd1 vccd1 _00443_ sky130_fd_sc_hd__inv_2
XFILLER_0_154_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14418_ clknet_leaf_163_wb_clk_i _02182_ _00783_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[772\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_71_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09114__S1 net1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08227__C1 net1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12023__B1 net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08244__A net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10924__D net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14349_ clknet_leaf_183_wb_clk_i _02113_ _00714_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[703\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_4_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xwire591 _04861_ vssd1 vssd1 vccd1 vccd1 net591 sky130_fd_sc_hd__buf_4
Xhold605 team_03_WB.instance_to_wrap.core.register_file.registers_state\[248\] vssd1
+ vssd1 vccd1 vccd1 net2098 sky130_fd_sc_hd__dlygate4sd3_1
Xhold616 team_03_WB.instance_to_wrap.core.register_file.registers_state\[237\] vssd1
+ vssd1 vccd1 vccd1 net2109 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10585__B1 net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold627 team_03_WB.instance_to_wrap.core.register_file.registers_state\[231\] vssd1
+ vssd1 vccd1 vccd1 net2120 sky130_fd_sc_hd__dlygate4sd3_1
Xhold638 team_03_WB.instance_to_wrap.core.register_file.registers_state\[753\] vssd1
+ vssd1 vccd1 vccd1 net2131 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_150_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold649 team_03_WB.instance_to_wrap.core.register_file.registers_state\[251\] vssd1
+ vssd1 vccd1 vccd1 net2142 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_51_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_08910_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[556\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[524\]
+ net979 vssd1 vssd1 vccd1 vccd1 _04852_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10713__S net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09890_ net320 _05437_ _05770_ net352 _05831_ vssd1 vssd1 vccd1 vccd1 _05832_ sky130_fd_sc_hd__a221o_2
XFILLER_0_111_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10888__A1 _06480_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08841_ _04781_ _04782_ net858 vssd1 vssd1 vccd1 vccd1 _04783_ sky130_fd_sc_hd__o21a_1
XFILLER_0_100_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08772_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[34\] net978
+ vssd1 vssd1 vccd1 vccd1 _04714_ sky130_fd_sc_hd__or2_1
XANTENNA__10014__A net94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07723_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[525\] net778
+ net747 _03664_ vssd1 vssd1 vccd1 vccd1 _03665_ sky130_fd_sc_hd__a211o_1
XANTENNA__11837__B1 net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06939__S0 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_2531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07654_ net1119 _03594_ _03595_ vssd1 vssd1 vccd1 vccd1 _03596_ sky130_fd_sc_hd__or3_1
XFILLER_0_67_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_0_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08419__A net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_0_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_146 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_228 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07585_ team_03_WB.instance_to_wrap.core.decoder.inst\[24\] net1020 vssd1 vssd1 vccd1
+ vccd1 _03527_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout344_A _06805_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1086_A net1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09324_ _04679_ _05252_ vssd1 vssd1 vccd1 vccd1 _05266_ sky130_fd_sc_hd__and2_1
XFILLER_0_47_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_146_831 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_153_3517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09255_ _05069_ _05195_ vssd1 vssd1 vccd1 vccd1 _05197_ sky130_fd_sc_hd__nor2_1
XFILLER_0_118_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10684__A _05429_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout511_A net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1253_A net1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout609_A _02938_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13060__A net1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_90_wb_clk_i_A clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_08206_ _04134_ _04147_ net850 vssd1 vssd1 vccd1 vccd1 _04148_ sky130_fd_sc_hd__mux2_8
XFILLER_0_69_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12014__B1 net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_170_3864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09186_ net434 net429 _04620_ net544 vssd1 vssd1 vccd1 vccd1 _05128_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_170_3875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08154__A team_03_WB.instance_to_wrap.core.decoder.inst\[19\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11368__A2 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_895 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08137_ _03567_ _04076_ _04077_ _04078_ vssd1 vssd1 vccd1 vccd1 _04079_ sky130_fd_sc_hd__nand4b_4
XFILLER_0_114_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10576__B1 net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1041_X net1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1139_X net1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_1998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_83_wb_clk_i clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_83_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__10040__A2 net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07441__B1 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08068_ net1186 team_03_WB.instance_to_wrap.core.register_file.registers_state\[726\]
+ net771 team_03_WB.instance_to_wrap.core.register_file.registers_state\[758\] net745
+ vssd1 vssd1 vccd1 vccd1 _04010_ sky130_fd_sc_hd__o221a_1
XANTENNA__11011__C net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout880_A net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout599_X net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout978_A net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11719__S net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07992__A1 net1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07019_ _02959_ _02960_ net1118 vssd1 vssd1 vccd1 vccd1 _02961_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_12_wb_clk_i clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_12_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__10623__S net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12404__A net1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10030_ team_03_WB.instance_to_wrap.BUSY_O team_03_WB.instance_to_wrap.wb.prev_BUSY_O
+ net1037 vssd1 vssd1 vccd1 vccd1 _05906_ sky130_fd_sc_hd__and3b_1
XFILLER_0_101_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10879__A1 net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout766_X net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11540__A2 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1098 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_1128 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11828__B1 net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout933_X net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11981_ net277 net2626 net444 vssd1 vssd1 vccd1 vccd1 _01563_ sky130_fd_sc_hd__mux2_1
X_13720_ clknet_leaf_186_wb_clk_i _01484_ _00085_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[74\]
+ sky130_fd_sc_hd__dfrtp_1
X_10932_ net838 _06517_ vssd1 vssd1 vccd1 vccd1 _06519_ sky130_fd_sc_hd__nor2_4
XANTENNA__10500__B1 net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_169_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_168_455 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13651_ clknet_leaf_96_wb_clk_i _01415_ _00016_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_10863_ net1252 net1018 net1251 vssd1 vssd1 vccd1 vccd1 _06462_ sky130_fd_sc_hd__and3b_1
XFILLER_0_38_111 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12602_ net1377 vssd1 vssd1 vccd1 vccd1 _00366_ sky130_fd_sc_hd__inv_2
XFILLER_0_112_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13582_ net1343 vssd1 vssd1 vccd1 vccd1 _01346_ sky130_fd_sc_hd__inv_2
XFILLER_0_137_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11056__B2 net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08457__C1 net1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10794_ _05799_ _05867_ vssd1 vssd1 vccd1 vccd1 _06404_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_155_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12533_ net1275 vssd1 vssd1 vccd1 vccd1 _00297_ sky130_fd_sc_hd__inv_2
XFILLER_0_136_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12005__A0 net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07680__B1 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12464_ net1410 vssd1 vssd1 vccd1 vccd1 _00228_ sky130_fd_sc_hd__inv_2
XFILLER_0_34_350 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14203_ clknet_leaf_122_wb_clk_i _01967_ _00568_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[557\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_34_372 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11415_ net272 net2735 net399 vssd1 vssd1 vccd1 vccd1 _02066_ sky130_fd_sc_hd__mux2_1
XANTENNA__09421__A1 net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10567__B1 net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12395_ net1281 vssd1 vssd1 vccd1 vccd1 _00159_ sky130_fd_sc_hd__inv_2
XANTENNA__12020__A3 net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14134_ clknet_leaf_178_wb_clk_i _01898_ _00499_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[488\]
+ sky130_fd_sc_hd__dfrtp_1
X_11346_ net515 net644 _06725_ net403 net2169 vssd1 vssd1 vccd1 vccd1 _02107_ sky130_fd_sc_hd__a32o_1
XFILLER_0_120_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07983__A1 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14065_ clknet_leaf_143_wb_clk_i _01829_ _00430_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[419\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08607__S0 net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12314__A net1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11277_ net1247 net837 net270 net670 vssd1 vssd1 vccd1 vccd1 _06706_ sky130_fd_sc_hd__and4_1
XANTENNA__07408__A net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13016_ net1375 vssd1 vssd1 vccd1 vccd1 _00780_ sky130_fd_sc_hd__inv_2
X_10228_ _06004_ _06069_ vssd1 vssd1 vccd1 vccd1 _06070_ sky130_fd_sc_hd__nor2_1
XANTENNA__07735__A1 team_03_WB.instance_to_wrap.core.decoder.inst\[23\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_135_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11531__A2 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2 team_03_WB.instance_to_wrap.SEL_I\[0\] vssd1 vssd1 vccd1 vccd1 net1495 sky130_fd_sc_hd__dlygate4sd3_1
X_10159_ _05041_ net660 vssd1 vssd1 vccd1 vccd1 _06001_ sky130_fd_sc_hd__and2_1
XFILLER_0_55_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_85_2114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11819__B1 net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14967_ clknet_leaf_91_wb_clk_i _02719_ _01332_ vssd1 vssd1 vccd1 vccd1 net219 sky130_fd_sc_hd__dfrtp_1
XANTENNA__12087__A3 net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1050 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13918_ clknet_leaf_119_wb_clk_i _01682_ _00283_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[272\]
+ sky130_fd_sc_hd__dfrtp_1
X_14898_ clknet_leaf_63_wb_clk_i _02661_ _01263_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.pc.current_pc\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_162_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08160__A1 net1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09910__X _05852_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_18_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13849_ clknet_leaf_162_wb_clk_i _01613_ _00214_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[203\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_119_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12984__A net1380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07370_ net721 _03311_ _03303_ _03296_ vssd1 vssd1 vccd1 vccd1 _03312_ sky130_fd_sc_hd__o2bb2a_4
XANTENNA__08448__C1 net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_174_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_831 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_935 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_155_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07120__C1 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09040_ net874 _04973_ _04976_ vssd1 vssd1 vccd1 vccd1 _04982_ sky130_fd_sc_hd__or3_1
XFILLER_0_154_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07671__B1 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12011__A3 net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold402 team_03_WB.instance_to_wrap.core.register_file.registers_state\[810\] vssd1
+ vssd1 vccd1 vccd1 net1895 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold413 team_03_WB.instance_to_wrap.core.register_file.registers_state\[437\] vssd1
+ vssd1 vccd1 vccd1 net1906 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_174_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_41_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold424 team_03_WB.instance_to_wrap.core.register_file.registers_state\[362\] vssd1
+ vssd1 vccd1 vccd1 net1917 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold435 team_03_WB.instance_to_wrap.core.register_file.registers_state\[49\] vssd1
+ vssd1 vccd1 vccd1 net1928 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold446 team_03_WB.instance_to_wrap.core.register_file.registers_state\[292\] vssd1
+ vssd1 vccd1 vccd1 net1939 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07974__A1 net1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold457 team_03_WB.instance_to_wrap.core.register_file.registers_state\[423\] vssd1
+ vssd1 vccd1 vccd1 net1950 sky130_fd_sc_hd__dlygate4sd3_1
Xhold468 team_03_WB.instance_to_wrap.CPU_DAT_O\[23\] vssd1 vssd1 vccd1 vccd1 net1961
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09942_ _05875_ net1866 net293 vssd1 vssd1 vccd1 vccd1 _02756_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_129_3018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold479 team_03_WB.instance_to_wrap.core.register_file.registers_state\[818\] vssd1
+ vssd1 vccd1 vccd1 net1972 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_3029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout904 _02844_ vssd1 vssd1 vccd1 vccd1 net904 sky130_fd_sc_hd__buf_4
XFILLER_0_0_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout915 net257 vssd1 vssd1 vccd1 vccd1 net915 sky130_fd_sc_hd__buf_2
XANTENNA__09715__A2 _05650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout926 net932 vssd1 vssd1 vccd1 vccd1 net926 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_74_1895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09873_ net352 _05422_ _05814_ net584 vssd1 vssd1 vccd1 vccd1 _05815_ sky130_fd_sc_hd__o22a_1
Xfanout937 net939 vssd1 vssd1 vccd1 vccd1 net937 sky130_fd_sc_hd__buf_4
Xfanout948 net949 vssd1 vssd1 vccd1 vccd1 net948 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout294_A _05859_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_146_3365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout959 net974 vssd1 vssd1 vccd1 vccd1 net959 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08923__B1 net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_146_3376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08824_ net1053 team_03_WB.instance_to_wrap.core.register_file.registers_state\[705\]
+ net1006 team_03_WB.instance_to_wrap.core.register_file.registers_state\[737\] net1077
+ vssd1 vssd1 vccd1 vccd1 _04766_ sky130_fd_sc_hd__a221o_1
Xhold1102 team_03_WB.instance_to_wrap.core.register_file.registers_state\[862\] vssd1
+ vssd1 vccd1 vccd1 net2595 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1113 team_03_WB.instance_to_wrap.core.register_file.registers_state\[149\] vssd1
+ vssd1 vccd1 vccd1 net2606 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1124 team_03_WB.instance_to_wrap.core.register_file.registers_state\[581\] vssd1
+ vssd1 vccd1 vccd1 net2617 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1001_A net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1135 team_03_WB.instance_to_wrap.core.register_file.registers_state\[850\] vssd1
+ vssd1 vccd1 vccd1 net2628 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1146 team_03_WB.instance_to_wrap.core.register_file.registers_state\[605\] vssd1
+ vssd1 vccd1 vccd1 net2639 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1157 team_03_WB.instance_to_wrap.wb.curr_state\[2\] vssd1 vssd1 vccd1 vccd1 net2650
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08755_ net942 _04694_ _04695_ _04696_ vssd1 vssd1 vccd1 vccd1 _04697_ sky130_fd_sc_hd__a22o_1
XFILLER_0_174_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10679__A net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout461_A net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1168 team_03_WB.instance_to_wrap.core.register_file.registers_state\[365\] vssd1
+ vssd1 vccd1 vccd1 net2661 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1179 team_03_WB.instance_to_wrap.core.register_file.registers_state\[894\] vssd1
+ vssd1 vccd1 vccd1 net2672 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout559_A net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07706_ net1104 team_03_WB.instance_to_wrap.core.register_file.registers_state\[237\]
+ net900 vssd1 vssd1 vccd1 vccd1 _03648_ sky130_fd_sc_hd__or3_1
XANTENNA__11286__A1 net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08686_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[1000\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[968\]
+ net975 vssd1 vssd1 vccd1 vccd1 _04628_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_130_wb_clk_i clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_130_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08151__A1 net1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07637_ net1094 team_03_WB.instance_to_wrap.core.register_file.registers_state\[334\]
+ net1157 vssd1 vssd1 vccd1 vccd1 _03579_ sky130_fd_sc_hd__a21o_1
XFILLER_0_95_537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_2837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_120_2848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout726_A net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1370_A net1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout347_X net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1089_X net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08439__C1 net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_172_3904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07568_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[536\] net804
+ net734 _03509_ vssd1 vssd1 vccd1 vccd1 _03510_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_172_3915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09307_ _04565_ _05248_ vssd1 vssd1 vccd1 vccd1 _05249_ sky130_fd_sc_hd__nor2_1
XANTENNA__10618__S net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08155__Y _04097_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout514_X net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07499_ _03433_ _03434_ _03439_ _03440_ net1120 net1140 vssd1 vssd1 vccd1 vccd1 _03441_
+ sky130_fd_sc_hd__mux4_1
X_09238_ _04323_ _05179_ vssd1 vssd1 vccd1 vccd1 _05180_ sky130_fd_sc_hd__nor2_1
XFILLER_0_1_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_160_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11022__B net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09169_ net435 net428 _04647_ net551 vssd1 vssd1 vccd1 vccd1 _05111_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_118_2799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15090__1476 vssd1 vssd1 vccd1 vccd1 _15090__1476/HI net1476 sky130_fd_sc_hd__conb_1
X_11200_ _06409_ net2342 net487 vssd1 vssd1 vccd1 vccd1 _02208_ sky130_fd_sc_hd__mux2_1
XFILLER_0_142_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07414__B1 net1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12180_ net1524 vssd1 vssd1 vccd1 vccd1 _02373_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_fanout883_X net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07965__A1 net1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11131_ net714 net694 net302 vssd1 vssd1 vccd1 vccd1 _06641_ sky130_fd_sc_hd__or3b_1
XFILLER_0_8_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold980 team_03_WB.instance_to_wrap.core.register_file.registers_state\[660\] vssd1
+ vssd1 vccd1 vccd1 net2473 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09167__B1 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold991 team_03_WB.instance_to_wrap.core.register_file.registers_state\[840\] vssd1
+ vssd1 vccd1 vccd1 net2484 sky130_fd_sc_hd__dlygate4sd3_1
X_11062_ net2569 net423 _06608_ net516 vssd1 vssd1 vccd1 vccd1 _02274_ sky130_fd_sc_hd__a22o_1
XFILLER_0_101_296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10013_ _03103_ net1740 net287 vssd1 vssd1 vccd1 vccd1 _02701_ sky130_fd_sc_hd__mux2_1
XANTENNA__08390__A1 net1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14821_ clknet_leaf_95_wb_clk_i net1774 _01186_ vssd1 vssd1 vccd1 vccd1 net141 sky130_fd_sc_hd__dfrtp_1
XANTENNA_input22_A DAT_I[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14752_ clknet_leaf_48_wb_clk_i _02516_ _01117_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_11964_ net640 _06741_ net476 net366 net1951 vssd1 vssd1 vccd1 vccd1 _01579_ sky130_fd_sc_hd__a32o_1
XANTENNA__08059__A net1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13703_ clknet_leaf_109_wb_clk_i _01467_ _00068_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[57\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10915_ net838 _06503_ vssd1 vssd1 vccd1 vccd1 _06505_ sky130_fd_sc_hd__nor2_2
XFILLER_0_169_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14683_ clknet_leaf_67_wb_clk_i _02447_ _01048_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.ADR_I\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_80_2011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09890__A1 net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11895_ net635 _06704_ net468 net373 net1963 vssd1 vssd1 vccd1 vccd1 _01646_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_80_2022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07350__C1 net1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09890__B2 net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11912__S net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13634_ net1434 vssd1 vssd1 vccd1 vccd1 _01398_ sky130_fd_sc_hd__inv_2
X_10846_ _06443_ _06444_ _06445_ net585 vssd1 vssd1 vccd1 vccd1 _06446_ sky130_fd_sc_hd__o211a_2
XFILLER_0_39_464 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13565_ net1421 vssd1 vssd1 vccd1 vccd1 _01329_ sky130_fd_sc_hd__inv_2
XFILLER_0_66_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10777_ net1252 net1018 vssd1 vssd1 vccd1 vccd1 _06387_ sky130_fd_sc_hd__nand2_8
XFILLER_0_171_428 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11213__A _06456_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12516_ net1366 vssd1 vssd1 vccd1 vccd1 _00280_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07653__B1 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13496_ net1341 vssd1 vssd1 vccd1 vccd1 _01260_ sky130_fd_sc_hd__inv_2
XFILLER_0_14_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_1076 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12447_ net1285 vssd1 vssd1 vccd1 vccd1 _00211_ sky130_fd_sc_hd__inv_2
XFILLER_0_152_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07405__B1 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08602__C1 net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12378_ net1372 vssd1 vssd1 vccd1 vccd1 _00142_ sky130_fd_sc_hd__inv_2
XANTENNA__07956__A1 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14117_ clknet_leaf_11_wb_clk_i _01881_ _00482_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[471\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11752__A2 net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11329_ net263 net2563 net406 vssd1 vssd1 vccd1 vccd1 _02116_ sky130_fd_sc_hd__mux2_1
X_15097_ net914 vssd1 vssd1 vccd1 vccd1 net255 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10960__A0 _06541_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07138__A net1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14048_ clknet_leaf_2_wb_clk_i _01812_ _00413_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[402\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07708__A1 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_52_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09173__A3 net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06870_ team_03_WB.instance_to_wrap.core.control_logic.instruction\[3\] team_03_WB.instance_to_wrap.core.control_logic.instruction\[2\]
+ team_03_WB.instance_to_wrap.core.control_logic.instruction\[1\] team_03_WB.instance_to_wrap.core.control_logic.instruction\[0\]
+ vssd1 vssd1 vccd1 vccd1 _02812_ sky130_fd_sc_hd__and4_1
XANTENNA__10712__B1 net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07184__A2 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08381__A1 net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11094__S net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_35 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_141_3262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08540_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[958\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[926\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[830\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[798\]
+ net965 net1072 vssd1 vssd1 vccd1 vccd1 _04482_ sky130_fd_sc_hd__mux4_1
XANTENNA__11268__A1 net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_141_3273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire315_X net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09640__X _05582_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08471_ net1218 _04411_ _04412_ vssd1 vssd1 vccd1 vccd1 _04413_ sky130_fd_sc_hd__o21ai_1
XANTENNA__11107__B _06523_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10786__X _06396_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07304__C net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_159_263 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07422_ net1084 team_03_WB.instance_to_wrap.core.register_file.registers_state\[884\]
+ net889 _03363_ net1125 vssd1 vssd1 vccd1 vccd1 _03364_ sky130_fd_sc_hd__o311a_1
XANTENNA__10491__A2 net1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07892__B1 net1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_163_907 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_1042 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07353_ net1114 _03291_ _03292_ vssd1 vssd1 vccd1 vccd1 _03295_ sky130_fd_sc_hd__or3_1
XFILLER_0_70_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09633__A1 net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_114_Left_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07644__B1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07284_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[9\] net788
+ net753 _03225_ vssd1 vssd1 vccd1 vccd1 _03226_ sky130_fd_sc_hd__a211o_1
XFILLER_0_66_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06998__A2 team_03_WB.instance_to_wrap.core.decoder.inst\[12\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_142_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09023_ net1244 team_03_WB.instance_to_wrap.core.register_file.registers_state\[336\]
+ net989 team_03_WB.instance_to_wrap.core.register_file.registers_state\[368\] net1078
+ vssd1 vssd1 vccd1 vccd1 _04965_ sky130_fd_sc_hd__o221a_1
XFILLER_0_170_450 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_832 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout307_A _06396_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1049_A net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold210 team_03_WB.instance_to_wrap.core.register_file.registers_state\[2\] vssd1
+ vssd1 vccd1 vccd1 net1703 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_76_1935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold221 _02575_ vssd1 vssd1 vccd1 vccd1 net1714 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_76_1946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold232 team_03_WB.instance_to_wrap.CPU_DAT_I\[8\] vssd1 vssd1 vccd1 vccd1 net1725
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_148_3405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold243 _02593_ vssd1 vssd1 vccd1 vccd1 net1736 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10173__S net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_148_3416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold254 _02586_ vssd1 vssd1 vccd1 vccd1 net1747 sky130_fd_sc_hd__dlygate4sd3_1
Xhold265 team_03_WB.instance_to_wrap.CPU_DAT_I\[31\] vssd1 vssd1 vccd1 vccd1 net1758
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold276 net226 vssd1 vssd1 vccd1 vccd1 net1769 sky130_fd_sc_hd__dlygate4sd3_1
Xhold287 _02589_ vssd1 vssd1 vccd1 vccd1 net1780 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_113_2696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1216_A team_03_WB.instance_to_wrap.core.decoder.inst\[17\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09962__S net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout701 _06559_ vssd1 vssd1 vccd1 vccd1 net701 sky130_fd_sc_hd__clkbuf_8
Xhold298 net223 vssd1 vssd1 vccd1 vccd1 net1791 sky130_fd_sc_hd__dlygate4sd3_1
X_09925_ _05646_ _05676_ _05856_ vssd1 vssd1 vccd1 vccd1 _05867_ sky130_fd_sc_hd__and3_1
XANTENNA__09815__X _05757_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout712 net713 vssd1 vssd1 vccd1 vccd1 net712 sky130_fd_sc_hd__clkbuf_4
Xfanout723 _02863_ vssd1 vssd1 vccd1 vccd1 net723 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_165_3763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout734 net737 vssd1 vssd1 vccd1 vccd1 net734 sky130_fd_sc_hd__buf_4
XANTENNA_fanout676_A _05948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_123_Left_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout297_X net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout745 net755 vssd1 vssd1 vccd1 vccd1 net745 sky130_fd_sc_hd__buf_4
Xfanout756 net758 vssd1 vssd1 vccd1 vccd1 net756 sky130_fd_sc_hd__clkbuf_4
X_09856_ _05080_ _05609_ _05791_ _05797_ vssd1 vssd1 vccd1 vccd1 _05798_ sky130_fd_sc_hd__o211a_4
Xfanout767 net770 vssd1 vssd1 vccd1 vccd1 net767 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout1004_X net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout778 net780 vssd1 vssd1 vccd1 vccd1 net778 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10703__B1 net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07335__X _03277_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout789 net790 vssd1 vssd1 vccd1 vccd1 net789 sky130_fd_sc_hd__buf_2
XANTENNA__08372__A1 net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08807_ net1055 team_03_WB.instance_to_wrap.core.register_file.registers_state\[321\]
+ net1004 team_03_WB.instance_to_wrap.core.register_file.registers_state\[353\] net1215
+ vssd1 vssd1 vccd1 vccd1 _04749_ sky130_fd_sc_hd__a221o_1
X_09787_ _02954_ _05508_ _05724_ _05728_ vssd1 vssd1 vccd1 vccd1 _05729_ sky130_fd_sc_hd__a211o_1
Xclkbuf_4_8__f_wb_clk_i clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_8__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_fanout843_A _06304_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06999_ team_03_WB.instance_to_wrap.core.decoder.inst\[13\] _02832_ vssd1 vssd1 vccd1
+ vccd1 _02941_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout464_X net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08738_ net434 net429 _04679_ net544 vssd1 vssd1 vccd1 vccd1 _04680_ sky130_fd_sc_hd__o31a_1
XFILLER_0_96_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_166_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout631_X net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08669_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[935\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[903\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[807\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[775\]
+ net989 net1078 vssd1 vssd1 vccd1 vccd1 _04611_ sky130_fd_sc_hd__mux4_1
XANTENNA__09872__A1 _05736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11732__S net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout729_X net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10700_ _02769_ _06315_ _02768_ vssd1 vssd1 vccd1 vccd1 _06338_ sky130_fd_sc_hd__o21a_1
XFILLER_0_95_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10482__A2 net1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11680_ _06722_ net379 net338 net2033 vssd1 vssd1 vccd1 vccd1 _01854_ sky130_fd_sc_hd__a22o_1
XFILLER_0_165_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_272 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10631_ team_03_WB.instance_to_wrap.core.decoder.inst\[30\] team_03_WB.instance_to_wrap.CPU_DAT_O\[30\]
+ net845 vssd1 vssd1 vccd1 vccd1 _02497_ sky130_fd_sc_hd__mux2_1
XFILLER_0_165_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_870 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11033__A net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13350_ net1342 vssd1 vssd1 vccd1 vccd1 _01114_ sky130_fd_sc_hd__inv_2
XFILLER_0_64_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10562_ net1837 net533 net600 _05872_ vssd1 vssd1 vccd1 vccd1 _02561_ sky130_fd_sc_hd__a22o_1
XANTENNA__08832__C1 net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12301_ net1331 vssd1 vssd1 vccd1 vccd1 _00065_ sky130_fd_sc_hd__inv_2
XFILLER_0_106_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13281_ net1404 vssd1 vssd1 vccd1 vccd1 _01045_ sky130_fd_sc_hd__inv_2
X_10493_ net107 net1029 net906 net1852 vssd1 vssd1 vccd1 vccd1 _02616_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_20_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15020_ clknet_leaf_94_wb_clk_i _02740_ _01385_ vssd1 vssd1 vccd1 vccd1 net176 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_20_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12232_ net1630 vssd1 vssd1 vccd1 vccd1 _01425_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__07884__C net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07399__C1 net1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08286__S1 net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11734__A2 _06519_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12163_ net1539 vssd1 vssd1 vccd1 vccd1 _02390_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_9_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11114_ _06631_ net2695 net418 vssd1 vssd1 vccd1 vccd1 _02245_ sky130_fd_sc_hd__mux2_1
X_12094_ _06792_ net456 net439 net2321 vssd1 vssd1 vccd1 vccd1 _01453_ sky130_fd_sc_hd__a22o_1
XFILLER_0_120_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09155__A3 _04267_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11045_ net2334 net422 _06599_ net503 vssd1 vssd1 vccd1 vccd1 _02282_ sky130_fd_sc_hd__a22o_1
XFILLER_0_127_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08363__A1 net1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07797__S0 net1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_48 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06913__A2 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14804_ clknet_leaf_83_wb_clk_i _02568_ _01169_ vssd1 vssd1 vccd1 vccd1 net135 sky130_fd_sc_hd__dfrtp_1
X_12996_ net1384 vssd1 vssd1 vccd1 vccd1 _00760_ sky130_fd_sc_hd__inv_2
XANTENNA__08115__B2 net1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14735_ clknet_leaf_31_wb_clk_i _02499_ _01100_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_8_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11947_ net620 _06724_ net452 net363 net2049 vssd1 vssd1 vccd1 vccd1 _01596_ sky130_fd_sc_hd__a32o_1
XFILLER_0_157_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1015 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_583 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14666_ clknet_leaf_7_wb_clk_i _02430_ _01031_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1020\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_74_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11878_ net627 _06687_ net458 net371 net2298 vssd1 vssd1 vccd1 vccd1 _01663_ sky130_fd_sc_hd__a32o_1
XANTENNA__07421__A net1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13617_ net1429 vssd1 vssd1 vccd1 vccd1 _01381_ sky130_fd_sc_hd__inv_2
X_10829_ net311 net310 net317 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[24\]
+ vssd1 vssd1 vccd1 vccd1 _06432_ sky130_fd_sc_hd__a31o_1
XANTENNA__09615__A1 _04778_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09076__C1 net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14597_ clknet_leaf_40_wb_clk_i _02361_ _00962_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[951\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_156_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_45_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13548_ net1324 vssd1 vssd1 vccd1 vccd1 _01312_ sky130_fd_sc_hd__inv_2
XFILLER_0_27_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08823__C1 net1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_2360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_2371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13479_ net1425 vssd1 vssd1 vccd1 vccd1 _01243_ sky130_fd_sc_hd__inv_2
XFILLER_0_113_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11089__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07929__A1 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_2279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11725__A2 _06479_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_68 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10933__B1 net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_1832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07971_ net750 _03911_ _03912_ net808 vssd1 vssd1 vccd1 vccd1 _03913_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_71_1843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09710_ _03682_ _05041_ _05651_ net666 vssd1 vssd1 vccd1 vccd1 _05652_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_143_3302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06922_ team_03_WB.instance_to_wrap.core.decoder.inst\[24\] net876 vssd1 vssd1 vccd1
+ vccd1 _02864_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_143_3313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09000__C1 net1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08398__S net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09083__A net1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09641_ net581 _05338_ _05564_ _05582_ vssd1 vssd1 vccd1 vccd1 _05583_ sky130_fd_sc_hd__a31o_4
X_06853_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[12\] vssd1
+ vssd1 vccd1 vccd1 _02796_ sky130_fd_sc_hd__inv_2
XFILLER_0_93_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_160_3660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11118__A net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09572_ _05513_ vssd1 vssd1 vccd1 vccd1 _05514_ sky130_fd_sc_hd__inv_2
XANTENNA__10022__A net84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09811__A net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08523_ net1227 team_03_WB.instance_to_wrap.core.register_file.registers_state\[95\]
+ net952 team_03_WB.instance_to_wrap.core.register_file.registers_state\[127\] net916
+ vssd1 vssd1 vccd1 vccd1 _04465_ sky130_fd_sc_hd__o221a_1
XFILLER_0_132_1007 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_183 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07034__C net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11661__A1 _06624_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08454_ net1062 _04394_ _04395_ net1074 vssd1 vssd1 vccd1 vccd1 _04396_ sky130_fd_sc_hd__a211o_1
XFILLER_0_37_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07969__C net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07405_ net1171 team_03_WB.instance_to_wrap.core.register_file.registers_state\[607\]
+ net758 team_03_WB.instance_to_wrap.core.register_file.registers_state\[639\] net1124
+ vssd1 vssd1 vccd1 vccd1 _03347_ sky130_fd_sc_hd__o221a_1
XFILLER_0_46_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08385_ _04150_ _04210_ _04269_ _04326_ net554 net567 vssd1 vssd1 vccd1 vccd1 _04327_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__09606__A1 _05547_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout424_A net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1166_A net1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07336_ team_03_WB.instance_to_wrap.core.decoder.inst\[31\] net826 vssd1 vssd1 vccd1
+ vccd1 _03278_ sky130_fd_sc_hd__and2_1
XANTENNA__07617__B1 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_951 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07267_ net1108 team_03_WB.instance_to_wrap.core.register_file.registers_state\[873\]
+ net902 vssd1 vssd1 vccd1 vccd1 _03209_ sky130_fd_sc_hd__or3_1
XFILLER_0_116_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_2736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11003__D net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07632__A3 net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1333_A net1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_314 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_115_2747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09006_ net1046 team_03_WB.instance_to_wrap.core.register_file.registers_state\[682\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[650\] net996 net933
+ vssd1 vssd1 vccd1 vccd1 _04948_ sky130_fd_sc_hd__o221a_1
XFILLER_0_61_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_170_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07198_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[50\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[18\]
+ net756 vssd1 vssd1 vccd1 vccd1 _03140_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_167_3803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout793_A net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1121_X net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_131_Left_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1219_X net1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09790__B1 net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout581_X net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout960_A net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout520 _06395_ vssd1 vssd1 vccd1 vccd1 net520 sky130_fd_sc_hd__clkbuf_8
Xfanout531 net532 vssd1 vssd1 vccd1 vccd1 net531 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout679_X net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11727__S net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout542 net543 vssd1 vssd1 vccd1 vccd1 net542 sky130_fd_sc_hd__clkbuf_2
X_09908_ _05518_ _05583_ _05849_ vssd1 vssd1 vccd1 vccd1 _05850_ sky130_fd_sc_hd__nand3_1
XANTENNA__10631__S net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout553 net554 vssd1 vssd1 vccd1 vccd1 net553 sky130_fd_sc_hd__clkbuf_4
Xfanout564 _03025_ vssd1 vssd1 vccd1 vccd1 net564 sky130_fd_sc_hd__clkbuf_4
Xfanout575 net576 vssd1 vssd1 vccd1 vccd1 net575 sky130_fd_sc_hd__buf_2
XANTENNA__08345__A1 net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout586 _06400_ vssd1 vssd1 vccd1 vccd1 net586 sky130_fd_sc_hd__clkbuf_4
X_09839_ net578 _05778_ _05779_ _05780_ _05078_ vssd1 vssd1 vccd1 vccd1 _05781_ sky130_fd_sc_hd__a311o_1
Xfanout597 _06464_ vssd1 vssd1 vccd1 vccd1 net597 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout846_X net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12850_ net1395 vssd1 vssd1 vccd1 vccd1 _00614_ sky130_fd_sc_hd__inv_2
XFILLER_0_69_824 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11801_ net2757 _06629_ net330 vssd1 vssd1 vccd1 vccd1 _01737_ sky130_fd_sc_hd__mux2_1
XANTENNA__11101__A0 _06505_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_3_1_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_1_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_12781_ net1275 vssd1 vssd1 vccd1 vccd1 _00545_ sky130_fd_sc_hd__inv_2
XANTENNA__07305__C1 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_140_Left_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14520_ clknet_leaf_187_wb_clk_i _02284_ _00885_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[874\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13243__A net1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11732_ net1938 _06509_ net335 vssd1 vssd1 vccd1 vccd1 _01804_ sky130_fd_sc_hd__mux2_1
XFILLER_0_139_745 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_827 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07320__A2 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07241__A net1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14451_ clknet_leaf_98_wb_clk_i _02215_ _00816_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[805\]
+ sky130_fd_sc_hd__dfrtp_1
X_11663_ net2047 _06626_ net344 vssd1 vssd1 vccd1 vccd1 _01870_ sky130_fd_sc_hd__mux2_1
XANTENNA__09058__C1 net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_153_Right_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_25_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13402_ net1406 vssd1 vssd1 vccd1 vccd1 _01166_ sky130_fd_sc_hd__inv_2
X_10614_ net2645 net1849 net840 vssd1 vssd1 vccd1 vccd1 _02514_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07608__B1 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14382_ clknet_leaf_128_wb_clk_i _02146_ _00747_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[736\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11594_ net298 net2482 net449 vssd1 vssd1 vccd1 vccd1 _01935_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13333_ net1325 vssd1 vssd1 vccd1 vccd1 _01097_ sky130_fd_sc_hd__inv_2
X_10545_ team_03_WB.instance_to_wrap.wb.curr_state\[0\] _06288_ vssd1 vssd1 vccd1
+ vccd1 _06289_ sky130_fd_sc_hd__nand2_1
XFILLER_0_122_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13264_ net1413 vssd1 vssd1 vccd1 vccd1 _01028_ sky130_fd_sc_hd__inv_2
XFILLER_0_122_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10476_ net1823 net1027 net905 team_03_WB.instance_to_wrap.ADR_I\[30\] vssd1 vssd1
+ vccd1 vccd1 _02633_ sky130_fd_sc_hd__a22o_1
XFILLER_0_33_982 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08072__A net1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15003_ clknet_leaf_59_wb_clk_i net51 _01368_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_150_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11707__A2 net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12215_ net1569 vssd1 vssd1 vccd1 vccd1 _02338_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_122_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13195_ net1287 vssd1 vssd1 vccd1 vccd1 _00959_ sky130_fd_sc_hd__inv_2
XFILLER_0_20_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07387__A2 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12146_ net1582 vssd1 vssd1 vccd1 vccd1 _02407_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__10391__A1 net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_159_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09128__A3 net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12077_ net619 _06640_ net452 net439 net1793 vssd1 vssd1 vccd1 vccd1 _01470_ sky130_fd_sc_hd__a32o_1
XFILLER_0_47_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11028_ net504 net653 _06588_ net422 net2044 vssd1 vssd1 vccd1 vccd1 _02288_ sky130_fd_sc_hd__a32o_1
XANTENNA__07416__A net1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_1018 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10143__A1 _04148_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11340__B1 net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10694__A2 _06316_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11891__A1 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12979_ net1265 vssd1 vssd1 vccd1 vccd1 _00743_ sky130_fd_sc_hd__inv_2
XFILLER_0_63_79 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14718_ clknet_leaf_50_wb_clk_i _02482_ _01083_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.decoder.inst\[15\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_86_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_99_2400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_2411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09049__C1 net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14649_ clknet_leaf_175_wb_clk_i _02413_ _01014_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1003\]
+ sky130_fd_sc_hd__dfstp_1
XPHY_EDGE_ROW_120_Right_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_64_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08170_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[820\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[788\]
+ net958 vssd1 vssd1 vccd1 vccd1 _04112_ sky130_fd_sc_hd__mux2_1
XANTENNA__08534__X _04476_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_136_3161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_3172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08498__S1 net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_95_2319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07121_ net614 _03059_ _03061_ vssd1 vssd1 vccd1 vccd1 _03063_ sky130_fd_sc_hd__a21o_1
XFILLER_0_6_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08272__B1 net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07052_ net1153 _02818_ _02809_ net1042 vssd1 vssd1 vccd1 vccd1 _02994_ sky130_fd_sc_hd__o2bb2a_4
XANTENNA__09078__A net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_54 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_876 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput112 net112 vssd1 vssd1 vccd1 vccd1 ADR_O[18] sky130_fd_sc_hd__buf_2
Xoutput123 net123 vssd1 vssd1 vccd1 vccd1 ADR_O[28] sky130_fd_sc_hd__clkbuf_4
XANTENNA__11120__B net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08024__B1 net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput134 net134 vssd1 vssd1 vccd1 vccd1 ADR_O[9] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_63_5 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput145 net145 vssd1 vssd1 vccd1 vccd1 DAT_O[18] sky130_fd_sc_hd__clkbuf_4
XANTENNA__10017__A net71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput156 net156 vssd1 vssd1 vccd1 vccd1 DAT_O[28] sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_110_2633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08575__A1 net1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput167 net167 vssd1 vssd1 vccd1 vccd1 DAT_O[9] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_110_2644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput178 net178 vssd1 vssd1 vccd1 vccd1 gpio_oeb[13] sky130_fd_sc_hd__buf_2
XFILLER_0_10_164 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput189 net189 vssd1 vssd1 vccd1 vccd1 gpio_oeb[24] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_162_3700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_162_3711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07954_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[823\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[791\]
+ net766 vssd1 vssd1 vccd1 vccd1 _03896_ sky130_fd_sc_hd__mux2_1
XANTENNA__07326__A net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06905_ net1148 net881 vssd1 vssd1 vccd1 vccd1 _02847_ sky130_fd_sc_hd__nand2_1
X_07885_ net1187 team_03_WB.instance_to_wrap.core.register_file.registers_state\[143\]
+ net877 net1152 vssd1 vssd1 vccd1 vccd1 _03827_ sky130_fd_sc_hd__o211a_1
XANTENNA__07535__C1 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout374_A _06813_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09624_ net575 _05565_ vssd1 vssd1 vccd1 vccd1 _05566_ sky130_fd_sc_hd__nand2_1
X_06836_ team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[17\] vssd1 vssd1 vccd1
+ vccd1 _02779_ sky130_fd_sc_hd__inv_2
XANTENNA__08856__S net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11882__A1 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_2584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09555_ _04778_ _05106_ _05489_ _05492_ _05496_ vssd1 vssd1 vccd1 vccd1 _05497_ sky130_fd_sc_hd__o2111ai_1
XFILLER_0_77_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_37_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_37_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__06884__B team_03_WB.instance_to_wrap.core.decoder.inst\[28\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1283_A net1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout639_A net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08506_ net548 _04417_ _04447_ vssd1 vssd1 vccd1 vccd1 _04448_ sky130_fd_sc_hd__o21ai_1
XANTENNA__10880__D_N team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[17\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13063__A net1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09486_ _05371_ _05404_ _05412_ _05427_ vssd1 vssd1 vccd1 vccd1 _05428_ sky130_fd_sc_hd__a211o_1
XFILLER_0_148_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08437_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[890\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[858\]
+ net964 vssd1 vssd1 vccd1 vccd1 _04379_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout1071_X net1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout806_A net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1169_X net1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08368_ net1236 team_03_WB.instance_to_wrap.core.register_file.registers_state\[598\]
+ net970 team_03_WB.instance_to_wrap.core.register_file.registers_state\[630\] net921
+ vssd1 vssd1 vccd1 vccd1 _04310_ sky130_fd_sc_hd__o221a_1
XFILLER_0_33_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07319_ net1185 team_03_WB.instance_to_wrap.core.register_file.registers_state\[61\]
+ net876 vssd1 vssd1 vccd1 vccd1 _03261_ sky130_fd_sc_hd__and3_1
XANTENNA__10626__S net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08299_ _04239_ _04240_ net864 vssd1 vssd1 vccd1 vccd1 _04241_ sky130_fd_sc_hd__a21o_1
XANTENNA__10070__B1 net1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10330_ team_03_WB.instance_to_wrap.core.pc.current_pc\[28\] _06168_ net678 vssd1
+ vssd1 vccd1 vccd1 _02662_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout796_X net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10261_ _06093_ _06102_ vssd1 vssd1 vccd1 vccd1 _06103_ sky130_fd_sc_hd__nand2_1
XFILLER_0_14_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08566__A1 net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12000_ net265 _06756_ net469 net444 net2516 vssd1 vssd1 vccd1 vccd1 _01544_ sky130_fd_sc_hd__a32o_1
XFILLER_0_100_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10192_ _04565_ net676 vssd1 vssd1 vccd1 vccd1 _06034_ sky130_fd_sc_hd__or2_1
XANTENNA__08620__A net1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout963_X net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1304 net1305 vssd1 vssd1 vccd1 vccd1 net1304 sky130_fd_sc_hd__clkbuf_4
Xfanout1315 net1330 vssd1 vssd1 vccd1 vccd1 net1315 sky130_fd_sc_hd__clkbuf_4
Xfanout1326 net1329 vssd1 vssd1 vccd1 vccd1 net1326 sky130_fd_sc_hd__buf_4
Xfanout1337 net1338 vssd1 vssd1 vccd1 vccd1 net1337 sky130_fd_sc_hd__buf_4
XANTENNA__08318__A1 net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1348 net1349 vssd1 vssd1 vccd1 vccd1 net1348 sky130_fd_sc_hd__buf_4
Xfanout361 _06817_ vssd1 vssd1 vccd1 vccd1 net361 sky130_fd_sc_hd__buf_6
Xfanout1359 net1364 vssd1 vssd1 vccd1 vccd1 net1359 sky130_fd_sc_hd__buf_4
Xfanout372 _06813_ vssd1 vssd1 vccd1 vccd1 net372 sky130_fd_sc_hd__clkbuf_4
Xfanout383 net387 vssd1 vssd1 vccd1 vccd1 net383 sky130_fd_sc_hd__buf_4
X_13951_ clknet_leaf_166_wb_clk_i _01715_ _00316_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[305\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11322__A0 _06628_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout394 net395 vssd1 vssd1 vccd1 vccd1 net394 sky130_fd_sc_hd__buf_4
XANTENNA__07526__C1 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12902_ net1300 vssd1 vssd1 vccd1 vccd1 _00666_ sky130_fd_sc_hd__inv_2
X_13882_ clknet_leaf_142_wb_clk_i _01646_ _00247_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[236\]
+ sky130_fd_sc_hd__dfrtp_1
X_12833_ net1262 vssd1 vssd1 vccd1 vccd1 _00597_ sky130_fd_sc_hd__inv_2
XFILLER_0_154_1062 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12764_ net1419 vssd1 vssd1 vccd1 vccd1 _00528_ sky130_fd_sc_hd__inv_2
XFILLER_0_57_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08067__A net1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14503_ clknet_leaf_110_wb_clk_i _02267_ _00868_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[857\]
+ sky130_fd_sc_hd__dfrtp_1
X_11715_ net1857 net302 net336 vssd1 vssd1 vccd1 vccd1 _01821_ sky130_fd_sc_hd__mux2_1
X_12695_ net1390 vssd1 vssd1 vccd1 vccd1 _00459_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_540 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11920__S net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14434_ clknet_leaf_174_wb_clk_i _02198_ _00799_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[788\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_42_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11646_ net2646 _06612_ net342 vssd1 vssd1 vccd1 vccd1 _01887_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_962 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput14 DAT_I[20] vssd1 vssd1 vccd1 vccd1 net14 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_142_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput25 DAT_I[30] vssd1 vssd1 vccd1 vccd1 net25 sky130_fd_sc_hd__buf_1
XANTENNA__08254__B1 net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14365_ clknet_leaf_24_wb_clk_i _02129_ _00730_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[719\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput36 gpio_in[11] vssd1 vssd1 vccd1 vccd1 net36 sky130_fd_sc_hd__clkbuf_1
X_11577_ net280 net2458 net447 vssd1 vssd1 vccd1 vccd1 _01952_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput47 gpio_in[22] vssd1 vssd1 vccd1 vccd1 net47 sky130_fd_sc_hd__clkbuf_1
Xinput58 gpio_in[33] vssd1 vssd1 vccd1 vccd1 net58 sky130_fd_sc_hd__clkbuf_1
X_13316_ net1326 vssd1 vssd1 vccd1 vccd1 _01080_ sky130_fd_sc_hd__inv_2
XFILLER_0_80_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10528_ net138 net1032 net1024 net1754 vssd1 vssd1 vccd1 vccd1 _02582_ sky130_fd_sc_hd__a22o_1
Xinput69 wbs_adr_i[11] vssd1 vssd1 vccd1 vccd1 net69 sky130_fd_sc_hd__buf_1
Xhold809 team_03_WB.instance_to_wrap.core.register_file.registers_state\[652\] vssd1
+ vssd1 vccd1 vccd1 net2302 sky130_fd_sc_hd__dlygate4sd3_1
X_14296_ clknet_leaf_19_wb_clk_i _02060_ _00661_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[650\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_90_2216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13247_ net1347 vssd1 vssd1 vccd1 vccd1 _01011_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_90_2227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_41_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_10459_ team_03_WB.instance_to_wrap.core.pc.current_pc\[4\] _06273_ net683 vssd1
+ vssd1 vccd1 vccd1 _02638_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08557__A1 net1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13178_ net1377 vssd1 vssd1 vccd1 vccd1 _00942_ sky130_fd_sc_hd__inv_2
XANTENNA__08530__A net1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10271__S net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12129_ net1502 vssd1 vssd1 vccd1 vccd1 _02424_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__08309__A1 net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12105__A2 net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_88_2178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07670_ net1177 team_03_WB.instance_to_wrap.core.register_file.registers_state\[222\]
+ vssd1 vssd1 vccd1 vccd1 _03612_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_88_2189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06985__A net1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09340_ _03170_ _05151_ vssd1 vssd1 vccd1 vccd1 _05282_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_90_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_3201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_3212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11040__C_N net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_902 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09271_ _05211_ _05212_ vssd1 vssd1 vccd1 vccd1 _05213_ sky130_fd_sc_hd__nand2_1
XANTENNA__07296__A1 net1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_2492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08493__B1 net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13611__A net1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08222_ net1241 team_03_WB.instance_to_wrap.core.register_file.registers_state\[977\]
+ net961 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1009\] net1225
+ vssd1 vssd1 vccd1 vccd1 _04164_ sky130_fd_sc_hd__o221a_1
XFILLER_0_62_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_236 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_80_wb_clk_i_A clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__08705__A _04646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10954__B _06536_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_578 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07048__A1 team_03_WB.instance_to_wrap.core.decoder.inst\[10\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07048__B2 net1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08153_ net860 _04091_ _04094_ vssd1 vssd1 vccd1 vccd1 _04095_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_71_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_155_wb_clk_i clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_155_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_151_3467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10052__B1 net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11131__A net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07104_ net1100 team_03_WB.instance_to_wrap.core.register_file.registers_state\[321\]
+ net801 team_03_WB.instance_to_wrap.core.register_file.registers_state\[353\] net1155
+ vssd1 vssd1 vccd1 vccd1 _03046_ sky130_fd_sc_hd__a221oi_1
XTAP_TAPCELL_ROW_151_3478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08084_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[790\] net793
+ net1041 _04025_ vssd1 vssd1 vccd1 vccd1 _04026_ sky130_fd_sc_hd__o211a_1
XANTENNA__11488__D _06463_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_941 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07035_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[3\] net801
+ net731 _02976_ vssd1 vssd1 vccd1 vccd1 _02977_ sky130_fd_sc_hd__o211a_1
XFILLER_0_3_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1031_A net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1129_A net1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09536__A _05477_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_294 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout491_A net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07756__C1 net1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10181__S net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08986_ net1045 team_03_WB.instance_to_wrap.core.register_file.registers_state\[74\]
+ net996 team_03_WB.instance_to_wrap.core.register_file.registers_state\[106\] net933
+ vssd1 vssd1 vccd1 vccd1 _04928_ sky130_fd_sc_hd__a221o_1
XANTENNA__09970__S net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07937_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[439\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[407\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[311\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[279\]
+ net766 net1128 vssd1 vssd1 vccd1 vccd1 _03879_ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout377_X net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout756_A net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07868_ net1201 team_03_WB.instance_to_wrap.core.register_file.registers_state\[475\]
+ net783 team_03_WB.instance_to_wrap.core.register_file.registers_state\[507\] net1158
+ vssd1 vssd1 vccd1 vccd1 _03810_ sky130_fd_sc_hd__o221a_1
XFILLER_0_39_1132 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_2982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08181__C1 net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08720__A1 net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09607_ _05548_ _05371_ vssd1 vssd1 vccd1 vccd1 _05549_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_27_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07799_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[11\] net797
+ net730 _03740_ vssd1 vssd1 vccd1 vccd1 _03741_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout923_A _04088_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09538_ _05306_ _05307_ _05311_ _05329_ vssd1 vssd1 vccd1 vccd1 _05480_ sky130_fd_sc_hd__nor4_1
XANTENNA__10210__A _02889_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08079__A3 net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09469_ _05410_ vssd1 vssd1 vccd1 vccd1 _05411_ sky130_fd_sc_hd__inv_2
XFILLER_0_148_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout711_X net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout809_X net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11500_ _06454_ net2246 net388 vssd1 vssd1 vccd1 vccd1 _02006_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12480_ net1400 vssd1 vssd1 vccd1 vccd1 _00244_ sky130_fd_sc_hd__inv_2
XFILLER_0_47_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11431_ net268 net2586 net398 vssd1 vssd1 vccd1 vccd1 _02053_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10043__B1 net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08787__A1 net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07134__S1 net1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11041__A net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14150_ clknet_leaf_28_wb_clk_i _01914_ _00515_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[504\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_34_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11362_ net495 net624 _06733_ net400 net1957 vssd1 vssd1 vccd1 vccd1 _02099_ sky130_fd_sc_hd__a32o_1
XFILLER_0_46_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13101_ net1292 vssd1 vssd1 vccd1 vccd1 _00865_ sky130_fd_sc_hd__inv_2
X_10313_ net282 _06154_ net677 vssd1 vssd1 vccd1 vccd1 _06155_ sky130_fd_sc_hd__o21a_1
XFILLER_0_0_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14081_ clknet_leaf_183_wb_clk_i _01845_ _00446_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[435\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_104_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09717__Y _05659_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10880__A net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11293_ net1249 net839 _06545_ net671 vssd1 vssd1 vccd1 vccd1 _06714_ sky130_fd_sc_hd__and4_1
XANTENNA__07518__X _03460_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13032_ net1297 vssd1 vssd1 vccd1 vccd1 _00796_ sky130_fd_sc_hd__inv_2
XANTENNA_input52_A gpio_in[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10244_ _05996_ _05999_ _06084_ _05994_ _05992_ vssd1 vssd1 vccd1 vccd1 _06086_ sky130_fd_sc_hd__o311a_2
XFILLER_0_30_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11543__B1 net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08634__S1 net1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1101 net1105 vssd1 vssd1 vccd1 vccd1 net1101 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07211__A1 net1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_125_wb_clk_i_A clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_100_670 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1112 net1113 vssd1 vssd1 vccd1 vccd1 net1112 sky130_fd_sc_hd__clkbuf_4
X_10175_ _03789_ _06015_ vssd1 vssd1 vccd1 vccd1 _06017_ sky130_fd_sc_hd__xnor2_1
Xfanout1123 net1124 vssd1 vssd1 vccd1 vccd1 net1123 sky130_fd_sc_hd__buf_4
Xfanout1134 net1137 vssd1 vssd1 vccd1 vccd1 net1134 sky130_fd_sc_hd__buf_4
Xfanout1145 team_03_WB.instance_to_wrap.core.ru.state\[0\] vssd1 vssd1 vccd1 vccd1
+ net1145 sky130_fd_sc_hd__buf_2
Xfanout1156 net1157 vssd1 vssd1 vccd1 vccd1 net1156 sky130_fd_sc_hd__buf_2
Xfanout1167 net1168 vssd1 vssd1 vccd1 vccd1 net1167 sky130_fd_sc_hd__buf_4
X_14983_ clknet_leaf_66_wb_clk_i net62 _01348_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1178 net1179 vssd1 vssd1 vccd1 vccd1 net1178 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_89_705 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1189 net1190 vssd1 vssd1 vccd1 vccd1 net1189 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11915__S net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13934_ clknet_leaf_126_wb_clk_i _01698_ _00299_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[288\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_44_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08172__C1 net1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08711__A1 net1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13865_ clknet_leaf_117_wb_clk_i _01629_ _00230_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[219\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_8_wb_clk_i_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_57_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12816_ net1411 vssd1 vssd1 vccd1 vccd1 _00580_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_83_2075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13796_ clknet_leaf_30_wb_clk_i _01560_ _00161_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[150\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_167_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12747_ net1288 vssd1 vssd1 vccd1 vccd1 _00511_ sky130_fd_sc_hd__inv_2
XFILLER_0_127_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11650__S net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_13_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12678_ net1300 vssd1 vssd1 vccd1 vccd1 _00442_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_13_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08525__A net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09120__S net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_404 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14417_ clknet_leaf_141_wb_clk_i _02181_ _00782_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[771\]
+ sky130_fd_sc_hd__dfrtp_1
X_11629_ _06703_ net384 net348 net2544 vssd1 vssd1 vccd1 vccd1 _01903_ sky130_fd_sc_hd__a22o_1
XANTENNA__12023__A1 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_163_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09975__A0 _02921_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10034__B1 net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08778__A1 net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14348_ clknet_leaf_16_wb_clk_i _02112_ _00713_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[702\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_164_wb_clk_i_A clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold606 team_03_WB.instance_to_wrap.core.register_file.registers_state\[38\] vssd1
+ vssd1 vccd1 vccd1 net2099 sky130_fd_sc_hd__dlygate4sd3_1
Xhold617 team_03_WB.instance_to_wrap.core.register_file.registers_state\[174\] vssd1
+ vssd1 vccd1 vccd1 net2110 sky130_fd_sc_hd__dlygate4sd3_1
Xwire592 _04739_ vssd1 vssd1 vccd1 vccd1 net592 sky130_fd_sc_hd__buf_4
XANTENNA__10585__B2 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold628 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[5\] vssd1 vssd1 vccd1
+ vccd1 net2121 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07450__A1 net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold639 team_03_WB.instance_to_wrap.core.register_file.registers_state\[483\] vssd1
+ vssd1 vccd1 vccd1 net2132 sky130_fd_sc_hd__dlygate4sd3_1
X_14279_ clknet_leaf_106_wb_clk_i _02043_ _00644_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[633\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_59_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09356__A net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07202__A1 net1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08840_ net1240 team_03_WB.instance_to_wrap.core.register_file.registers_state\[128\]
+ net990 team_03_WB.instance_to_wrap.core.register_file.registers_state\[160\] net946
+ vssd1 vssd1 vccd1 vccd1 _04782_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_55_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08771_ net551 _04712_ _04680_ vssd1 vssd1 vccd1 vccd1 _04713_ sky130_fd_sc_hd__a21o_1
XFILLER_0_109_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15059__1445 vssd1 vssd1 vccd1 vccd1 _15059__1445/HI net1445 sky130_fd_sc_hd__conb_1
XFILLER_0_97_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07722_ net1197 team_03_WB.instance_to_wrap.core.register_file.registers_state\[557\]
+ net884 vssd1 vssd1 vccd1 vccd1 _03664_ sky130_fd_sc_hd__and3_1
XANTENNA__11837__A1 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07163__X _03105_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08702__A1 net1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06939__S1 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_2532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07653_ net1094 team_03_WB.instance_to_wrap.core.register_file.registers_state\[974\]
+ net796 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1006\] net1131
+ vssd1 vssd1 vccd1 vccd1 _03595_ sky130_fd_sc_hd__a221oi_1
XTAP_TAPCELL_ROW_0_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11126__A net1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07584_ net722 _03500_ _03506_ _03525_ vssd1 vssd1 vccd1 vccd1 _03526_ sky130_fd_sc_hd__o31a_4
XFILLER_0_149_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09323_ _05263_ _05264_ _05256_ vssd1 vssd1 vccd1 vccd1 _05265_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_122_2890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_146_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10965__A net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_153_3507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_153_3518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09254_ _05069_ _05195_ vssd1 vssd1 vccd1 vccd1 _05196_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout1079_A net1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_145_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08205_ net867 _04145_ _04146_ vssd1 vssd1 vccd1 vccd1 _04147_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_106_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09185_ _04824_ _04831_ _05126_ _05123_ vssd1 vssd1 vccd1 vccd1 _05127_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout504_A net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_170_3865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1246_A team_03_WB.instance_to_wrap.core.decoder.inst\[15\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08136_ _03352_ _03391_ _03428_ _03903_ vssd1 vssd1 vccd1 vccd1 _04078_ sky130_fd_sc_hd__and4_1
XANTENNA__10576__B2 _05886_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11773__B1 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07441__A1 net1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_1999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08067_ net1186 team_03_WB.instance_to_wrap.core.register_file.registers_state\[598\]
+ vssd1 vssd1 vccd1 vccd1 _04009_ sky130_fd_sc_hd__or2_1
XANTENNA__10904__S net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1034_X net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1413_A net1436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07338__X _03280_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09266__A _05041_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07018_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[931\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[899\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[803\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[771\]
+ net780 net1133 vssd1 vssd1 vccd1 vccd1 _02960_ sky130_fd_sc_hd__mux4_1
XANTENNA_clkbuf_4_15__f_wb_clk_i_X clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout494_X net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout873_A net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07729__C1 net1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09194__A1 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10879__A2 net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1201_X net1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08941__A1 net1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_52_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_52_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout661_X net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08969_ _04909_ _04910_ net1223 vssd1 vssd1 vccd1 vccd1 _04911_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout759_X net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11735__S net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11980_ _06426_ net2614 net443 vssd1 vssd1 vccd1 vccd1 _01564_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_546 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10931_ _06517_ vssd1 vssd1 vccd1 vccd1 _06518_ sky130_fd_sc_hd__inv_2
XFILLER_0_168_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout926_X net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11036__A net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10862_ net1248 _06388_ _06459_ vssd1 vssd1 vccd1 vccd1 _06461_ sky130_fd_sc_hd__o21ai_1
X_13650_ clknet_leaf_117_wb_clk_i _01414_ _00015_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_156_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12601_ net1357 vssd1 vssd1 vccd1 vccd1 _00365_ sky130_fd_sc_hd__inv_2
XFILLER_0_38_123 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13581_ net1433 vssd1 vssd1 vccd1 vccd1 _01345_ sky130_fd_sc_hd__inv_2
XANTENNA__11056__A2 net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10793_ _05799_ _05867_ vssd1 vssd1 vccd1 vccd1 _06403_ sky130_fd_sc_hd__and2b_1
XFILLER_0_137_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_1124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13251__A net1358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12532_ net1310 vssd1 vssd1 vccd1 vccd1 _00296_ sky130_fd_sc_hd__inv_2
XFILLER_0_81_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_163_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07680__A1 net1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12463_ net1336 vssd1 vssd1 vccd1 vccd1 _00227_ sky130_fd_sc_hd__inv_2
XFILLER_0_152_835 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14202_ clknet_leaf_148_wb_clk_i _01966_ _00567_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[556\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_34_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11414_ net2521 net396 _06753_ net501 vssd1 vssd1 vccd1 vccd1 _02067_ sky130_fd_sc_hd__a22o_1
X_12394_ net1279 vssd1 vssd1 vccd1 vccd1 _00158_ sky130_fd_sc_hd__inv_2
XANTENNA__09421__A2 net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10881__Y _06477_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11764__B1 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07968__C1 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14133_ clknet_leaf_129_wb_clk_i _01897_ _00498_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[487\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_104_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11345_ net277 net715 net699 vssd1 vssd1 vccd1 vccd1 _06725_ sky130_fd_sc_hd__and3_1
XFILLER_0_1_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15119__1488 vssd1 vssd1 vccd1 vccd1 _15119__1488/HI net1488 sky130_fd_sc_hd__conb_1
XFILLER_0_132_592 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07395__S net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09709__B1 net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14064_ clknet_leaf_121_wb_clk_i _01828_ _00429_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[418\]
+ sky130_fd_sc_hd__dfrtp_1
X_11276_ net505 net633 _06705_ net410 net2079 vssd1 vssd1 vccd1 vccd1 _02157_ sky130_fd_sc_hd__a32o_1
XANTENNA__11516__A0 net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08607__S1 net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_18_Left_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13015_ net1385 vssd1 vssd1 vccd1 vccd1 _00779_ sky130_fd_sc_hd__inv_2
X_10227_ _06009_ _06012_ _06065_ _06006_ _06002_ vssd1 vssd1 vccd1 vccd1 _06069_ sky130_fd_sc_hd__a311oi_4
XANTENNA__08393__C1 net1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10158_ team_03_WB.instance_to_wrap.core.pc.current_pc\[13\] net660 vssd1 vssd1 vccd1
+ vccd1 _06000_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_33_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3 team_03_WB.instance_to_wrap.core.register_file.registers_state\[944\] vssd1
+ vssd1 vccd1 vccd1 net1496 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11645__S net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10089_ net594 _05519_ _05540_ _05932_ vssd1 vssd1 vccd1 vccd1 _05933_ sky130_fd_sc_hd__o211a_1
X_14966_ clknet_leaf_101_wb_clk_i _02718_ _01331_ vssd1 vssd1 vccd1 vccd1 net218 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_85_2126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08145__C1 net1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07043__S0 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13917_ clknet_leaf_26_wb_clk_i _01681_ _00282_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[271\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14897_ clknet_leaf_63_wb_clk_i _02660_ _01262_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.pc.current_pc\[26\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_18_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08954__S net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13848_ clknet_leaf_173_wb_clk_i _01612_ _00213_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[202\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08448__B1 net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13779_ clknet_leaf_109_wb_clk_i _01543_ _00144_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[133\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_100_2440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07671__A1 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10007__A0 _03488_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_142_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10791__Y _06401_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1011 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10558__B2 _05868_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11755__B1 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_3_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold403 team_03_WB.instance_to_wrap.core.register_file.registers_state\[696\] vssd1
+ vssd1 vccd1 vccd1 net1896 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold414 team_03_WB.instance_to_wrap.core.register_file.registers_state\[699\] vssd1
+ vssd1 vccd1 vccd1 net1907 sky130_fd_sc_hd__dlygate4sd3_1
Xhold425 team_03_WB.instance_to_wrap.core.register_file.registers_state\[804\] vssd1
+ vssd1 vccd1 vccd1 net1918 sky130_fd_sc_hd__dlygate4sd3_1
Xhold436 team_03_WB.instance_to_wrap.core.register_file.registers_state\[318\] vssd1
+ vssd1 vccd1 vccd1 net1929 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_57_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold447 team_03_WB.instance_to_wrap.core.register_file.registers_state\[311\] vssd1
+ vssd1 vccd1 vccd1 net1940 sky130_fd_sc_hd__dlygate4sd3_1
Xhold458 team_03_WB.instance_to_wrap.core.register_file.registers_state\[169\] vssd1
+ vssd1 vccd1 vccd1 net1951 sky130_fd_sc_hd__dlygate4sd3_1
X_09941_ _03900_ net663 vssd1 vssd1 vccd1 vccd1 _05875_ sky130_fd_sc_hd__nor2_1
Xhold469 net208 vssd1 vssd1 vccd1 vccd1 net1962 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_3019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout905 net906 vssd1 vssd1 vccd1 vccd1 net905 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_0_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout916 net923 vssd1 vssd1 vccd1 vccd1 net916 sky130_fd_sc_hd__clkbuf_4
Xfanout927 net932 vssd1 vssd1 vccd1 vccd1 net927 sky130_fd_sc_hd__clkbuf_4
X_09872_ _05734_ _05736_ net573 vssd1 vssd1 vccd1 vccd1 _05814_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_286 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_1896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout938 net939 vssd1 vssd1 vccd1 vccd1 net938 sky130_fd_sc_hd__buf_2
Xfanout949 _04087_ vssd1 vssd1 vccd1 vccd1 net949 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_146_3366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08823_ net1053 team_03_WB.instance_to_wrap.core.register_file.registers_state\[577\]
+ net1006 team_03_WB.instance_to_wrap.core.register_file.registers_state\[609\] net1215
+ vssd1 vssd1 vccd1 vccd1 _04765_ sky130_fd_sc_hd__a221o_1
Xhold1103 team_03_WB.instance_to_wrap.core.register_file.registers_state\[583\] vssd1
+ vssd1 vccd1 vccd1 net2596 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_146_3377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1114 team_03_WB.instance_to_wrap.core.register_file.registers_state\[879\] vssd1
+ vssd1 vccd1 vccd1 net2607 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06934__B1 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_7__f_wb_clk_i clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_7__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_fanout287_A net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1125 team_03_WB.instance_to_wrap.core.register_file.registers_state\[927\] vssd1
+ vssd1 vccd1 vccd1 net2618 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_31_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1136 team_03_WB.instance_to_wrap.core.register_file.registers_state\[133\] vssd1
+ vssd1 vccd1 vccd1 net2629 sky130_fd_sc_hd__dlygate4sd3_1
X_08754_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[515\] net1004
+ net926 vssd1 vssd1 vccd1 vccd1 _04696_ sky130_fd_sc_hd__o21a_1
Xhold1147 team_03_WB.instance_to_wrap.core.register_file.registers_state\[836\] vssd1
+ vssd1 vccd1 vccd1 net2640 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1158 team_03_WB.instance_to_wrap.core.register_file.registers_state\[732\] vssd1
+ vssd1 vccd1 vccd1 net2651 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1169 team_03_WB.instance_to_wrap.core.register_file.registers_state\[641\] vssd1
+ vssd1 vccd1 vccd1 net2662 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_124_2930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07705_ net1197 team_03_WB.instance_to_wrap.core.register_file.registers_state\[77\]
+ net778 team_03_WB.instance_to_wrap.core.register_file.registers_state\[109\] net731
+ vssd1 vssd1 vccd1 vccd1 _03647_ sky130_fd_sc_hd__o221a_1
X_08685_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[936\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[904\]
+ net975 vssd1 vssd1 vccd1 vccd1 _04627_ sky130_fd_sc_hd__mux2_1
XANTENNA__11286__A2 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout454_A net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1196_A net1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10494__B1 net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07053__B _02994_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07636_ net1192 team_03_WB.instance_to_wrap.core.register_file.registers_state\[366\]
+ net881 vssd1 vssd1 vccd1 vccd1 _03578_ sky130_fd_sc_hd__and3_1
XFILLER_0_49_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_120_2838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_120_2849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_165_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07621__X _03563_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07567_ net1106 team_03_WB.instance_to_wrap.core.register_file.registers_state\[568\]
+ net903 vssd1 vssd1 vccd1 vccd1 _03509_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_172_3905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10695__A _05583_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_170_wb_clk_i clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_170_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout621_A net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1363_A net1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_172_3916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09306_ net526 _05247_ vssd1 vssd1 vccd1 vccd1 _05248_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_119_843 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout719_A net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13071__A net1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07498_ _03435_ _03436_ net752 vssd1 vssd1 vccd1 vccd1 _03440_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11994__A0 net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09237_ _04032_ _05154_ vssd1 vssd1 vccd1 vccd1 _05179_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_17_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07662__A1 net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1151_X net1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07500__C net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10982__X _06560_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout507_X net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1249_X net1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09168_ _05108_ _05109_ vssd1 vssd1 vccd1 vccd1 _05110_ sky130_fd_sc_hd__nor2_1
XFILLER_0_16_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11022__C net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_2789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_160_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout990_A net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_687 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11746__B1 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07414__A1 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08119_ net1087 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1018\]
+ net892 _04060_ net1151 vssd1 vssd1 vccd1 vccd1 _04061_ sky130_fd_sc_hd__o311a_1
XFILLER_0_82_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10634__S net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08611__B1 net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09099_ net852 _05027_ _05040_ vssd1 vssd1 vccd1 vccd1 _05041_ sky130_fd_sc_hd__o21ba_4
XFILLER_0_160_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11130_ net491 net647 _06640_ net412 net1816 vssd1 vssd1 vccd1 vccd1 _02238_ sky130_fd_sc_hd__a32o_1
XANTENNA__07965__A2 net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11761__A3 net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold970 team_03_WB.instance_to_wrap.core.register_file.registers_state\[486\] vssd1
+ vssd1 vccd1 vccd1 net2463 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout876_X net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold981 team_03_WB.instance_to_wrap.core.register_file.registers_state\[269\] vssd1
+ vssd1 vccd1 vccd1 net2474 sky130_fd_sc_hd__dlygate4sd3_1
Xhold992 team_03_WB.instance_to_wrap.core.register_file.registers_state\[129\] vssd1
+ vssd1 vccd1 vccd1 net2485 sky130_fd_sc_hd__dlygate4sd3_1
X_11061_ net657 net707 net266 net830 vssd1 vssd1 vccd1 vccd1 _06608_ sky130_fd_sc_hd__and4_1
X_10012_ _03059_ net1704 net287 vssd1 vssd1 vccd1 vccd1 _02702_ sky130_fd_sc_hd__mux2_1
XANTENNA__10721__A1 _05623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14820_ clknet_leaf_104_wb_clk_i net1719 _01185_ vssd1 vssd1 vccd1 vccd1 net140 sky130_fd_sc_hd__dfrtp_1
XANTENNA__13246__A net1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input15_A DAT_I[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14751_ clknet_leaf_50_wb_clk_i _02515_ _01116_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11963_ net624 _06740_ net455 net363 net2092 vssd1 vssd1 vccd1 vccd1 _01580_ sky130_fd_sc_hd__a32o_1
XFILLER_0_98_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_169_743 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10485__B1 net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13702_ clknet_leaf_74_wb_clk_i _01466_ _00067_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[56\]
+ sky130_fd_sc_hd__dfrtp_1
X_10914_ _06503_ vssd1 vssd1 vccd1 vccd1 _06504_ sky130_fd_sc_hd__inv_2
XFILLER_0_98_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14682_ clknet_leaf_81_wb_clk_i _02446_ _01047_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.ADR_I\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_168_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11894_ net637 _06703_ net469 net373 net2109 vssd1 vssd1 vccd1 vccd1 _01647_ sky130_fd_sc_hd__a32o_1
XFILLER_0_58_229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_2012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_538 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10876__Y _06473_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_2023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10845_ net685 _05596_ vssd1 vssd1 vccd1 vccd1 _06445_ sky130_fd_sc_hd__nand2_1
X_13633_ net1417 vssd1 vssd1 vccd1 vccd1 _01397_ sky130_fd_sc_hd__inv_2
XFILLER_0_41_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_651 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10776_ net1252 net1018 vssd1 vssd1 vccd1 vccd1 _06386_ sky130_fd_sc_hd__and2_1
X_13564_ net1416 vssd1 vssd1 vccd1 vccd1 _01328_ sky130_fd_sc_hd__inv_2
XANTENNA__10788__A1 team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[31\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11985__A0 _06446_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07653__A1 net1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12515_ net1356 vssd1 vssd1 vccd1 vccd1 _00279_ sky130_fd_sc_hd__inv_2
XANTENNA__11213__B _06478_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13495_ net1340 vssd1 vssd1 vccd1 vccd1 _01259_ sky130_fd_sc_hd__inv_2
XFILLER_0_54_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15058__1444 vssd1 vssd1 vccd1 vccd1 _15058__1444/HI net1444 sky130_fd_sc_hd__conb_1
XFILLER_0_152_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12446_ net1390 vssd1 vssd1 vccd1 vccd1 _00210_ sky130_fd_sc_hd__inv_2
XFILLER_0_152_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07405__A1 net1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_738 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12377_ net1365 vssd1 vssd1 vccd1 vccd1 _00141_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_26_Left_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11328_ _06631_ net2422 net406 vssd1 vssd1 vccd1 vccd1 _02117_ sky130_fd_sc_hd__mux2_1
X_14116_ clknet_leaf_29_wb_clk_i _01880_ _00481_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[470\]
+ sky130_fd_sc_hd__dfrtp_1
X_15096_ net912 vssd1 vssd1 vccd1 vccd1 net248 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11259_ net709 _06468_ net827 vssd1 vssd1 vccd1 vccd1 _06697_ sky130_fd_sc_hd__and3_1
X_14047_ clknet_leaf_170_wb_clk_i _01811_ _00412_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[401\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07853__S net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06916__B1 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_167_Right_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_173_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_141_3263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14949_ clknet_leaf_101_wb_clk_i _02701_ _01314_ vssd1 vssd1 vccd1 vccd1 net206 sky130_fd_sc_hd__dfrtp_1
XANTENNA__11268__A2 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_141_3274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_35_Left_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10476__B1 net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_516 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08470_ net1062 _04409_ _04410_ vssd1 vssd1 vccd1 vccd1 _04412_ sky130_fd_sc_hd__or3_1
XFILLER_0_89_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14983__Q team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[2\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07421_ net1176 team_03_WB.instance_to_wrap.core.register_file.registers_state\[852\]
+ vssd1 vssd1 vccd1 vccd1 _03363_ sky130_fd_sc_hd__or2_1
XFILLER_0_159_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07352_ net1160 _03293_ vssd1 vssd1 vccd1 vccd1 _03294_ sky130_fd_sc_hd__or2_1
XFILLER_0_163_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11976__A0 net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_174_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07644__A1 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_312 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07283_ net1205 team_03_WB.instance_to_wrap.core.register_file.registers_state\[41\]
+ net886 vssd1 vssd1 vccd1 vccd1 _03225_ sky130_fd_sc_hd__and3_1
XFILLER_0_31_1098 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08841__B1 net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_142_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09022_ net856 _04962_ _04963_ _04961_ vssd1 vssd1 vccd1 vccd1 _04964_ sky130_fd_sc_hd__o31a_1
XFILLER_0_170_462 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold200 net179 vssd1 vssd1 vccd1 vccd1 net1693 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold211 net233 vssd1 vssd1 vccd1 vccd1 net1704 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_354 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_1936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold222 team_03_WB.instance_to_wrap.CPU_DAT_O\[13\] vssd1 vssd1 vccd1 vccd1 net1715
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_76_1947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold233 _02579_ vssd1 vssd1 vccd1 vccd1 net1726 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_148_3406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold244 team_03_WB.instance_to_wrap.core.register_file.registers_state\[52\] vssd1
+ vssd1 vccd1 vccd1 net1737 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07329__A net1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold255 net211 vssd1 vssd1 vccd1 vccd1 net1748 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_148_3417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold266 _02602_ vssd1 vssd1 vccd1 vccd1 net1759 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10951__A1 team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[4\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09149__A1 net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_2697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold277 team_03_WB.instance_to_wrap.core.register_file.registers_state\[302\] vssd1
+ vssd1 vccd1 vccd1 net1770 sky130_fd_sc_hd__dlygate4sd3_1
Xhold288 net219 vssd1 vssd1 vccd1 vccd1 net1781 sky130_fd_sc_hd__dlygate4sd3_1
X_09924_ net313 _05863_ _05864_ _05429_ vssd1 vssd1 vccd1 vccd1 _05866_ sky130_fd_sc_hd__or4b_1
Xhold299 team_03_WB.instance_to_wrap.core.register_file.registers_state\[167\] vssd1
+ vssd1 vccd1 vccd1 net1792 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout702 _06559_ vssd1 vssd1 vccd1 vccd1 net702 sky130_fd_sc_hd__buf_2
Xfanout713 net716 vssd1 vssd1 vccd1 vccd1 net713 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_165_3753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout724 _02863_ vssd1 vssd1 vccd1 vccd1 net724 sky130_fd_sc_hd__buf_4
XFILLER_0_0_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1111_A net1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout735 net737 vssd1 vssd1 vccd1 vccd1 net735 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_165_3764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout746 net749 vssd1 vssd1 vccd1 vccd1 net746 sky130_fd_sc_hd__buf_4
X_09855_ _05795_ _05796_ _05081_ _05794_ vssd1 vssd1 vccd1 vccd1 _05797_ sky130_fd_sc_hd__a211o_1
Xfanout757 net758 vssd1 vssd1 vccd1 vccd1 net757 sky130_fd_sc_hd__buf_2
XANTENNA_input7_A DAT_I[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10703__A1 net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout571_A net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout768 net769 vssd1 vssd1 vccd1 vccd1 net768 sky130_fd_sc_hd__clkbuf_4
Xfanout779 net780 vssd1 vssd1 vccd1 vccd1 net779 sky130_fd_sc_hd__clkbuf_2
XANTENNA__11900__B1 net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout669_A _06564_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08806_ _04744_ _04747_ net868 vssd1 vssd1 vccd1 vccd1 _04748_ sky130_fd_sc_hd__o21ai_1
X_09786_ net322 _05384_ _05727_ vssd1 vssd1 vccd1 vccd1 _05728_ sky130_fd_sc_hd__a21o_1
X_06998_ _02792_ team_03_WB.instance_to_wrap.core.decoder.inst\[12\] _02939_ vssd1
+ vssd1 vccd1 vccd1 _02940_ sky130_fd_sc_hd__o21ba_1
XPHY_EDGE_ROW_134_Right_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08737_ net852 _04663_ _04678_ vssd1 vssd1 vccd1 vccd1 _04679_ sky130_fd_sc_hd__o21ai_4
XANTENNA_fanout457_X net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout836_A net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1199_X net1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08124__A2 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08668_ _04608_ _04609_ vssd1 vssd1 vccd1 vccd1 _04610_ sky130_fd_sc_hd__and2_1
XANTENNA__11017__C net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07332__B1 net1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07883__A1 net1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07619_ net808 _03549_ _03550_ vssd1 vssd1 vccd1 vccd1 _03561_ sky130_fd_sc_hd__or3_1
X_08599_ _04539_ _04540_ net856 vssd1 vssd1 vccd1 vccd1 _04541_ sky130_fd_sc_hd__a21o_1
XANTENNA__10629__S net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout624_X net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_165_245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10630_ team_03_WB.instance_to_wrap.core.decoder.inst\[31\] net2228 net845 vssd1
+ vssd1 vccd1 vccd1 _02498_ sky130_fd_sc_hd__mux2_1
XFILLER_0_113_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_284 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11967__B1 net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07096__C1 net1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10561_ net1925 net531 net598 _05871_ vssd1 vssd1 vccd1 vccd1 _02562_ sky130_fd_sc_hd__a22o_1
XANTENNA__07635__A1 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07230__C net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12300_ net1333 vssd1 vssd1 vccd1 vccd1 _00064_ sky130_fd_sc_hd__inv_2
XFILLER_0_91_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13280_ net1407 vssd1 vssd1 vccd1 vccd1 _01044_ sky130_fd_sc_hd__inv_2
X_10492_ net108 net1029 net907 net1658 vssd1 vssd1 vccd1 vccd1 _02617_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout993_X net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12231_ net1652 vssd1 vssd1 vccd1 vccd1 _01426_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_161_484 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11195__B2 net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12162_ net1547 vssd1 vssd1 vccd1 vccd1 _02391_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__11734__A3 net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10942__A1 _06524_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11113_ net835 _06541_ vssd1 vssd1 vccd1 vccd1 _06631_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_9_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12093_ _06791_ net468 net441 net2149 vssd1 vssd1 vccd1 vccd1 _01454_ sky130_fd_sc_hd__a22o_1
X_11044_ net632 _06598_ vssd1 vssd1 vccd1 vccd1 _06599_ sky130_fd_sc_hd__nor2_1
XANTENNA__07797__S1 net1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07571__B1 net1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14803_ clknet_leaf_55_wb_clk_i _02567_ _01168_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.BUSY_O
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA_input18_X net18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_101_Right_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_157_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12995_ net1371 vssd1 vssd1 vccd1 vccd1 _00759_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11923__S net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14734_ clknet_leaf_44_wb_clk_i _02498_ _01099_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.decoder.inst\[31\]
+ sky130_fd_sc_hd__dfrtp_4
X_11946_ net640 _06723_ net463 net364 net1935 vssd1 vssd1 vccd1 vccd1 _01597_ sky130_fd_sc_hd__a32o_1
XFILLER_0_143_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07323__B1 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09863__A2 net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_169_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14665_ clknet_leaf_78_wb_clk_i _02429_ _01030_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1019\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_129_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11877_ net625 _06686_ net455 net371 net2058 vssd1 vssd1 vccd1 vccd1 _01664_ sky130_fd_sc_hd__a32o_1
XFILLER_0_28_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11224__A _06456_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13616_ net1417 vssd1 vssd1 vccd1 vccd1 _01380_ sky130_fd_sc_hd__inv_2
X_10828_ net692 _05499_ vssd1 vssd1 vccd1 vccd1 _06431_ sky130_fd_sc_hd__or2_1
XANTENNA__09076__B1 net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09615__A2 _05551_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14596_ clknet_leaf_22_wb_clk_i _02360_ _00961_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[950\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_54_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11958__B1 net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_171_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_45_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13547_ net1324 vssd1 vssd1 vccd1 vccd1 _01311_ sky130_fd_sc_hd__inv_2
XANTENNA__08823__B1 net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07140__C net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10759_ _02774_ _06294_ vssd1 vssd1 vccd1 vccd1 _06373_ sky130_fd_sc_hd__nand2_1
XFILLER_0_54_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07848__S net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10630__A0 team_03_WB.instance_to_wrap.core.decoder.inst\[31\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09629__A _03314_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_2361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11973__A3 net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_2372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13478_ net1424 vssd1 vssd1 vccd1 vccd1 _01242_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12429_ net1311 vssd1 vssd1 vccd1 vccd1 _00193_ sky130_fd_sc_hd__inv_2
XFILLER_0_168_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10933__A1 net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07970_ net1193 team_03_WB.instance_to_wrap.core.register_file.registers_state\[208\]
+ vssd1 vssd1 vccd1 vccd1 _03912_ sky130_fd_sc_hd__or2_1
X_15079_ net1465 vssd1 vssd1 vccd1 vccd1 la_data_out[15] sky130_fd_sc_hd__buf_2
XANTENNA__06988__A team_03_WB.instance_to_wrap.core.decoder.inst\[14\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_1833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06921_ team_03_WB.instance_to_wrap.core.decoder.inst\[24\] net876 vssd1 vssd1 vccd1
+ vccd1 _02863_ sky130_fd_sc_hd__and2_4
XTAP_TAPCELL_ROW_143_3303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09000__B1 net995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_143_3314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07157__A3 net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09640_ _05371_ _05569_ _05581_ vssd1 vssd1 vccd1 vccd1 _05582_ sky130_fd_sc_hd__a21bo_1
X_06852_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[44\] vssd1
+ vssd1 vccd1 vccd1 _02795_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_109_wb_clk_i clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_109_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_160_3650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_160_3661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09571_ net576 _05371_ vssd1 vssd1 vccd1 vccd1 _05513_ sky130_fd_sc_hd__and2_2
XANTENNA__11118__B net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08522_ net934 _04462_ _04463_ vssd1 vssd1 vccd1 vccd1 _04464_ sky130_fd_sc_hd__o21a_1
XFILLER_0_77_302 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_171_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_1019 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07314__B1 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_195 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08511__C1 net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08453_ net1228 team_03_WB.instance_to_wrap.core.register_file.registers_state\[988\]
+ net954 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1020\] net1218
+ vssd1 vssd1 vccd1 vccd1 _04395_ sky130_fd_sc_hd__o221a_1
XFILLER_0_147_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_519 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07404_ net1124 _03342_ _03343_ _03345_ net1138 vssd1 vssd1 vccd1 vccd1 _03346_ sky130_fd_sc_hd__a311o_1
XANTENNA__11134__A net1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_163_705 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08384_ net548 _04296_ _04325_ vssd1 vssd1 vccd1 vccd1 _04326_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_147_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_163_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11949__B1 net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07617__A1 net1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07335_ net722 _03260_ _03269_ _03276_ vssd1 vssd1 vccd1 vccd1 _03277_ sky130_fd_sc_hd__o2bb2a_4
XFILLER_0_46_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10973__A team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[0\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1061_A net1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout417_A _06610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09539__A net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07266_ net612 _03205_ _03207_ vssd1 vssd1 vccd1 vccd1 _03208_ sky130_fd_sc_hd__o21ai_2
XANTENNA__11964__A3 net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_115_2737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09005_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[554\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[522\]
+ net955 vssd1 vssd1 vccd1 vccd1 _04947_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_624 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07197_ _03138_ vssd1 vssd1 vccd1 vccd1 _03139_ sky130_fd_sc_hd__inv_2
XANTENNA__08162__B net995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_167_3804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1326_A net1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11177__B2 net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08578__C1 net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_460 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09973__S net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09826__X _05768_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08042__A1 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout786_A net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1114_X net1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout510 net517 vssd1 vssd1 vccd1 vccd1 net510 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07493__S net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09274__A _04953_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout521 _06395_ vssd1 vssd1 vccd1 vccd1 net521 sky130_fd_sc_hd__buf_4
Xfanout532 net533 vssd1 vssd1 vccd1 vccd1 net532 sky130_fd_sc_hd__clkbuf_4
X_09907_ _05541_ _05842_ vssd1 vssd1 vccd1 vccd1 _05849_ sky130_fd_sc_hd__nor2_1
Xfanout543 _03106_ vssd1 vssd1 vccd1 vccd1 net543 sky130_fd_sc_hd__buf_2
Xfanout554 _03064_ vssd1 vssd1 vccd1 vccd1 net554 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout953_A net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout565 _03025_ vssd1 vssd1 vccd1 vccd1 net565 sky130_fd_sc_hd__buf_2
XANTENNA__10688__B1 net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout576 net577 vssd1 vssd1 vccd1 vccd1 net576 sky130_fd_sc_hd__clkbuf_2
X_09838_ net578 _05670_ vssd1 vssd1 vccd1 vccd1 _05780_ sky130_fd_sc_hd__nor2_1
Xfanout598 net599 vssd1 vssd1 vccd1 vccd1 net598 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07553__B1 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15057__1443 vssd1 vssd1 vccd1 vccd1 _15057__1443/HI net1443 sky130_fd_sc_hd__conb_1
X_09769_ _04775_ _05106_ vssd1 vssd1 vccd1 vccd1 _05711_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout741_X net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout839_X net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11800_ net2127 _06519_ net328 vssd1 vssd1 vccd1 vccd1 _01738_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12780_ net1333 vssd1 vssd1 vccd1 vccd1 _00544_ sky130_fd_sc_hd__inv_2
XANTENNA__08177__X _04119_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07305__B1 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10867__B net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07081__X _03023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11731_ net596 _06505_ net456 _06808_ net1745 vssd1 vssd1 vccd1 vccd1 _01805_ sky130_fd_sc_hd__a32o_1
XFILLER_0_68_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_139_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_711 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_96_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11044__A net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14450_ clknet_leaf_163_wb_clk_i _02214_ _00815_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[804\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11662_ net2696 _06625_ net344 vssd1 vssd1 vccd1 vccd1 _01871_ sky130_fd_sc_hd__mux2_1
XANTENNA__09058__B1 net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13401_ net1424 vssd1 vssd1 vccd1 vccd1 _01165_ sky130_fd_sc_hd__inv_2
XFILLER_0_154_738 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_850 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10613_ net1606 team_03_WB.instance_to_wrap.CPU_DAT_O\[16\] net841 vssd1 vssd1 vccd1
+ vccd1 _02515_ sky130_fd_sc_hd__mux2_1
XANTENNA__07608__A1 net1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11593_ net271 net2309 net449 vssd1 vssd1 vccd1 vccd1 _01936_ sky130_fd_sc_hd__mux2_1
X_14381_ clknet_leaf_188_wb_clk_i _02145_ _00746_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[735\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10883__A net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_148_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_1123 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10544_ team_03_WB.instance_to_wrap.WRITE_I team_03_WB.instance_to_wrap.READ_I vssd1
+ vssd1 vccd1 vccd1 _06288_ sky130_fd_sc_hd__xnor2_1
X_13332_ net1319 vssd1 vssd1 vccd1 vccd1 _01096_ sky130_fd_sc_hd__inv_2
XANTENNA_input82_A wbs_adr_i[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11955__A3 net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08353__A _04294_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10475_ net127 net1027 net905 net1587 vssd1 vssd1 vccd1 vccd1 _02634_ sky130_fd_sc_hd__a22o_1
XFILLER_0_161_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13263_ net1339 vssd1 vssd1 vccd1 vccd1 _01027_ sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_31_wb_clk_i_A clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15002_ clknet_leaf_51_wb_clk_i net50 _01367_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_33_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12214_ net1498 vssd1 vssd1 vccd1 vccd1 _02339_ sky130_fd_sc_hd__clkbuf_1
X_13194_ net1284 vssd1 vssd1 vccd1 vccd1 _00958_ sky130_fd_sc_hd__inv_2
XANTENNA__10107__B net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_7_wb_clk_i clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_7_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_12145_ net1727 vssd1 vssd1 vccd1 vccd1 _02408_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__11918__S net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1070 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10822__S net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10391__A2 _06144_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12076_ _06782_ net458 net439 net1932 vssd1 vssd1 vccd1 vccd1 _01471_ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_1020 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11027_ net706 net271 net831 vssd1 vssd1 vccd1 vccd1 _06588_ sky130_fd_sc_hd__and3_1
XFILLER_0_21_1075 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11340__A1 net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08741__C1 net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09912__A _05706_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11653__S net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08087__X _04029_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12978_ net1395 vssd1 vssd1 vccd1 vccd1 _00742_ sky130_fd_sc_hd__inv_2
XANTENNA__07432__A net1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14717_ clknet_leaf_68_wb_clk_i _02481_ _01082_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.decoder.inst\[14\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_47_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11929_ _06505_ net2633 net369 vssd1 vssd1 vccd1 vccd1 _01613_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_47_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_908 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_2401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14648_ clknet_leaf_3_wb_clk_i _02412_ _01013_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1002\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__09049__B1 net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_2412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_716 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_70_wb_clk_i_A clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_27_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_738 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14579_ clknet_leaf_98_wb_clk_i _02343_ _00944_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[933\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_136_3162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_136_3173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07120_ net723 _03058_ _03043_ net617 vssd1 vssd1 vccd1 vccd1 _03062_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_103_75 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11946__A3 net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire587_A _05883_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08263__A net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07051_ net614 net593 _02991_ vssd1 vssd1 vccd1 vccd1 _02993_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_3_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_140_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_112 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_408 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_600 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_66 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput113 net113 vssd1 vssd1 vccd1 vccd1 ADR_O[19] sky130_fd_sc_hd__clkbuf_4
Xoutput124 net124 vssd1 vssd1 vccd1 vccd1 ADR_O[29] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_3_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08024__A1 net1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput135 net135 vssd1 vssd1 vccd1 vccd1 CYC_O sky130_fd_sc_hd__clkbuf_4
XANTENNA__10906__A1 net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10017__B net70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput146 net146 vssd1 vssd1 vccd1 vccd1 DAT_O[19] sky130_fd_sc_hd__buf_2
Xoutput157 net157 vssd1 vssd1 vccd1 vccd1 DAT_O[29] sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_110_2634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput168 net168 vssd1 vssd1 vccd1 vccd1 SEL_O[0] sky130_fd_sc_hd__clkbuf_4
Xoutput179 net179 vssd1 vssd1 vccd1 vccd1 gpio_oeb[14] sky130_fd_sc_hd__clkbuf_4
XANTENNA__10732__S net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_2645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_176 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_162_3701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08202__S net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07953_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[919\] net793
+ _03892_ net1152 vssd1 vssd1 vccd1 vccd1 _03895_ sky130_fd_sc_hd__o211a_1
XANTENNA__11129__A net1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06904_ net1139 net901 vssd1 vssd1 vccd1 vccd1 _02846_ sky130_fd_sc_hd__nor2_1
X_07884_ net1090 team_03_WB.instance_to_wrap.core.register_file.registers_state\[175\]
+ net894 vssd1 vssd1 vccd1 vccd1 _03826_ sky130_fd_sc_hd__or3_1
XFILLER_0_173_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07535__B1 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08732__C1 net1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09623_ _05482_ _05494_ net570 vssd1 vssd1 vccd1 vccd1 _05565_ sky130_fd_sc_hd__mux2_1
X_06835_ team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[29\] vssd1 vssd1 vccd1
+ vccd1 _02778_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_108_2585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout367_A _06814_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13344__A net1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_2596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09554_ net320 _05495_ vssd1 vssd1 vccd1 vccd1 _05496_ sky130_fd_sc_hd__nand2_1
XANTENNA__06884__C team_03_WB.instance_to_wrap.core.decoder.inst\[27\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08505_ net541 net431 net425 _04444_ vssd1 vssd1 vccd1 vccd1 _04447_ sky130_fd_sc_hd__or4_1
X_09485_ net320 _05419_ _05422_ net583 _05426_ vssd1 vssd1 vccd1 vccd1 _05427_ sky130_fd_sc_hd__a221o_1
XANTENNA__11634__A2 net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout534_A _06298_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10842__A0 net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09968__S net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08436_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[1018\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[986\]
+ net964 vssd1 vssd1 vccd1 vccd1 _04378_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_77_wb_clk_i clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_77_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_148_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_22_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08367_ _04303_ _04308_ net872 vssd1 vssd1 vccd1 vccd1 _04309_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1064_X net1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07318_ net817 _03258_ _03259_ _03251_ _03254_ vssd1 vssd1 vccd1 vccd1 _03260_ sky130_fd_sc_hd__a32o_1
XANTENNA__09269__A net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07066__A2 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08298_ net1242 team_03_WB.instance_to_wrap.core.register_file.registers_state\[184\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[152\] net987 net928
+ vssd1 vssd1 vccd1 vccd1 _04240_ sky130_fd_sc_hd__a221o_1
XFILLER_0_2_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07249_ net1191 team_03_WB.instance_to_wrap.core.register_file.registers_state\[168\]
+ vssd1 vssd1 vccd1 vccd1 _03191_ sky130_fd_sc_hd__and2_1
XFILLER_0_171_590 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_983 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_588 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_966 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1329_X net1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10260_ _06098_ _06101_ vssd1 vssd1 vccd1 vccd1 _06102_ sky130_fd_sc_hd__nor2_1
XFILLER_0_131_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09212__B1 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout691_X net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout789_X net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09763__A1 net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10191_ team_03_WB.instance_to_wrap.core.pc.current_pc\[5\] net675 vssd1 vssd1 vccd1
+ vccd1 _06033_ sky130_fd_sc_hd__nand2_1
XANTENNA__10642__S net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_115_wb_clk_i_A clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_79_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1305 net1309 vssd1 vssd1 vccd1 vccd1 net1305 sky130_fd_sc_hd__clkbuf_4
Xfanout1316 net1317 vssd1 vssd1 vccd1 vccd1 net1316 sky130_fd_sc_hd__buf_4
Xfanout1327 net1328 vssd1 vssd1 vccd1 vccd1 net1327 sky130_fd_sc_hd__buf_4
XANTENNA_fanout956_X net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout340 _06806_ vssd1 vssd1 vccd1 vccd1 net340 sky130_fd_sc_hd__clkbuf_8
Xfanout1338 net1339 vssd1 vssd1 vccd1 vccd1 net1338 sky130_fd_sc_hd__buf_4
Xfanout351 _04831_ vssd1 vssd1 vccd1 vccd1 net351 sky130_fd_sc_hd__clkbuf_4
Xfanout1349 net1358 vssd1 vssd1 vccd1 vccd1 net1349 sky130_fd_sc_hd__clkbuf_4
Xfanout362 _06817_ vssd1 vssd1 vccd1 vccd1 net362 sky130_fd_sc_hd__clkbuf_4
Xfanout373 _06813_ vssd1 vssd1 vccd1 vccd1 net373 sky130_fd_sc_hd__clkbuf_8
X_13950_ clknet_leaf_118_wb_clk_i _01714_ _00315_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[304\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout384 net387 vssd1 vssd1 vccd1 vccd1 net384 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07526__B1 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout395 _06757_ vssd1 vssd1 vccd1 vccd1 net395 sky130_fd_sc_hd__clkbuf_8
X_12901_ net1351 vssd1 vssd1 vccd1 vccd1 _00665_ sky130_fd_sc_hd__inv_2
XFILLER_0_88_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13881_ clknet_leaf_162_wb_clk_i _01645_ _00246_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[235\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07541__A3 net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13254__A net1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12832_ net1399 vssd1 vssd1 vccd1 vccd1 _00596_ sky130_fd_sc_hd__inv_2
XANTENNA__09818__A2 _04679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_1074 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11086__A0 _06454_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_1047 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11625__A2 net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12763_ net1360 vssd1 vssd1 vccd1 vccd1 _00527_ sky130_fd_sc_hd__inv_2
XFILLER_0_84_603 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_863 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14502_ clknet_leaf_72_wb_clk_i _02266_ _00867_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[856\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10833__B1 _06401_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11714_ net1891 net279 net335 vssd1 vssd1 vccd1 vccd1 _01822_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12694_ net1281 vssd1 vssd1 vccd1 vccd1 _00458_ sky130_fd_sc_hd__inv_2
XFILLER_0_127_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14433_ clknet_leaf_181_wb_clk_i _02197_ _00798_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[787\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10817__S net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11645_ net2372 _06611_ net343 vssd1 vssd1 vccd1 vccd1 _01888_ sky130_fd_sc_hd__mux2_1
XFILLER_0_140_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_42_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14364_ clknet_leaf_153_wb_clk_i _02128_ _00729_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[718\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput15 DAT_I[21] vssd1 vssd1 vccd1 vccd1 net15 sky130_fd_sc_hd__buf_1
Xinput26 DAT_I[31] vssd1 vssd1 vccd1 vccd1 net26 sky130_fd_sc_hd__clkbuf_1
XANTENNA_clkbuf_leaf_154_wb_clk_i_A clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_11576_ net281 net2119 net447 vssd1 vssd1 vccd1 vccd1 _01953_ sky130_fd_sc_hd__mux2_1
XANTENNA__08083__A net1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput37 gpio_in[12] vssd1 vssd1 vccd1 vccd1 net37 sky130_fd_sc_hd__clkbuf_1
Xinput48 gpio_in[23] vssd1 vssd1 vccd1 vccd1 net48 sky130_fd_sc_hd__clkbuf_1
X_13315_ net1335 vssd1 vssd1 vccd1 vccd1 _01079_ sky130_fd_sc_hd__inv_2
Xinput59 gpio_in[34] vssd1 vssd1 vccd1 vccd1 net59 sky130_fd_sc_hd__clkbuf_1
X_10527_ net139 net1032 net1024 net1821 vssd1 vssd1 vccd1 vccd1 _02583_ sky130_fd_sc_hd__a22o_1
XFILLER_0_150_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14295_ clknet_leaf_78_wb_clk_i _02059_ _00660_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[649\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_131_3070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09907__A _05541_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10458_ _06272_ _06271_ net286 vssd1 vssd1 vccd1 vccd1 _06273_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_90_2217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13246_ net1413 vssd1 vssd1 vccd1 vccd1 _01010_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_2228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11648__S net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09754__A1 net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10389_ _05994_ _05995_ _06085_ vssd1 vssd1 vccd1 vccd1 _06217_ sky130_fd_sc_hd__and3_1
XFILLER_0_0_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13177_ net1365 vssd1 vssd1 vccd1 vccd1 _00941_ sky130_fd_sc_hd__inv_2
XANTENNA__11875__C net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07765__B1 net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08962__C1 net1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12128_ net1637 vssd1 vssd1 vccd1 vccd1 _02425_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__09506__A1 _04778_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12059_ _06625_ net2641 net357 vssd1 vssd1 vccd1 vccd1 _01487_ sky130_fd_sc_hd__mux2_1
XANTENNA__07517__A0 _03430_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08714__C1 net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_2179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_318 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09809__A2 _04565_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11077__A0 _06616_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_66_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11616__A2 net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_3202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_138_3213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_157_340 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09270_ net591 _05210_ vssd1 vssd1 vccd1 vccd1 _05212_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_103_2482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08493__A1 net1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_2493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09690__B1 _05631_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14991__Q team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[10\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08221_ _04157_ _04162_ net871 vssd1 vssd1 vccd1 vccd1 _04163_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_155_3560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08152_ net854 _04092_ _04093_ vssd1 vssd1 vccd1 vccd1 _04094_ sky130_fd_sc_hd__or3_1
XANTENNA__08245__A1 net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_99_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07103_ net1100 team_03_WB.instance_to_wrap.core.register_file.registers_state\[449\]
+ vssd1 vssd1 vccd1 vccd1 _03045_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_151_3468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11131__B net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1004 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_706 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_151_3479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10052__B2 team_03_WB.instance_to_wrap.CPU_DAT_O\[11\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07453__C1 net1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08083_ net1088 team_03_WB.instance_to_wrap.core.register_file.registers_state\[822\]
+ net894 vssd1 vssd1 vccd1 vccd1 _04025_ sky130_fd_sc_hd__or3_1
X_15056__1442 vssd1 vssd1 vccd1 vccd1 _15056__1442/HI net1442 sky130_fd_sc_hd__conb_1
XFILLER_0_141_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07034_ net1099 team_03_WB.instance_to_wrap.core.register_file.registers_state\[35\]
+ net898 vssd1 vssd1 vccd1 vccd1 _02976_ sky130_fd_sc_hd__or3_1
XFILLER_0_113_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07205__C1 net1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_124_wb_clk_i clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_124_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout1024_A net1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09028__S net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08985_ _04925_ _04926_ net855 vssd1 vssd1 vccd1 vccd1 _04927_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout484_A _06779_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07771__A3 net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07936_ net1181 team_03_WB.instance_to_wrap.core.register_file.registers_state\[471\]
+ net766 team_03_WB.instance_to_wrap.core.register_file.registers_state\[503\] net1152
+ vssd1 vssd1 vccd1 vccd1 _03878_ sky130_fd_sc_hd__o221a_1
XFILLER_0_39_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07508__B1 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout651_A net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout272_X net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07867_ net1201 team_03_WB.instance_to_wrap.core.register_file.registers_state\[347\]
+ net784 team_03_WB.instance_to_wrap.core.register_file.registers_state\[379\] net1136
+ vssd1 vssd1 vccd1 vccd1 _03809_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_127_2983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1144 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1393_A net1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout749_A net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09606_ _05546_ _05547_ net574 vssd1 vssd1 vccd1 vccd1 _05548_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07798_ net1097 team_03_WB.instance_to_wrap.core.register_file.registers_state\[43\]
+ net900 vssd1 vssd1 vccd1 vccd1 _03740_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_27_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07072__A net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1079 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09537_ net594 _05456_ _05457_ _05478_ vssd1 vssd1 vccd1 vccd1 _05479_ sky130_fd_sc_hd__o31a_1
XANTENNA_fanout537_X net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout916_A net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1181_X net1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10815__B1 _06401_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09468_ net559 _05101_ _05103_ _05409_ net569 vssd1 vssd1 vccd1 vccd1 _05410_ sky130_fd_sc_hd__o311a_1
XANTENNA__09681__B1 _05622_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07800__A net1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_308 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08419_ net854 _04359_ _04360_ vssd1 vssd1 vccd1 vccd1 _04361_ sky130_fd_sc_hd__or3_1
XFILLER_0_81_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10637__S _06303_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout704_X net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09399_ _03352_ _04475_ vssd1 vssd1 vccd1 vccd1 _05341_ sky130_fd_sc_hd__nor2_1
XFILLER_0_93_488 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09659__S1 net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_708 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08236__A1 net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11430_ net511 _06537_ _06756_ net398 net2027 vssd1 vssd1 vccd1 vccd1 _02054_ sky130_fd_sc_hd__a32o_1
XFILLER_0_34_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12032__A2 net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10043__A1 net14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11361_ net1249 net838 _06477_ net669 vssd1 vssd1 vccd1 vccd1 _06733_ sky130_fd_sc_hd__and4_1
XANTENNA__11240__B1 net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10312_ team_03_WB.instance_to_wrap.core.pc.current_pc\[31\] _06153_ vssd1 vssd1
+ vccd1 vccd1 _06154_ sky130_fd_sc_hd__xnor2_1
X_13100_ net1313 vssd1 vssd1 vccd1 vccd1 _00864_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11791__A1 _06479_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14080_ clknet_leaf_187_wb_clk_i _01844_ _00445_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[434\]
+ sky130_fd_sc_hd__dfrtp_1
X_11292_ net507 net635 _06713_ net410 net2020 vssd1 vssd1 vccd1 vccd1 _02149_ sky130_fd_sc_hd__a32o_1
XFILLER_0_132_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10880__B net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09197__C1 net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10243_ _05999_ _06084_ vssd1 vssd1 vccd1 vccd1 _06085_ sky130_fd_sc_hd__or2_1
XFILLER_0_120_958 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13031_ net1369 vssd1 vssd1 vccd1 vccd1 _00795_ sky130_fd_sc_hd__inv_2
XANTENNA__11543__A1 net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07247__A net1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08944__C1 net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input45_A gpio_in[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10174_ team_03_WB.instance_to_wrap.core.decoder.inst\[30\] net826 _06015_ vssd1
+ vssd1 vccd1 vccd1 _06016_ sky130_fd_sc_hd__and3_1
Xfanout1102 net1104 vssd1 vssd1 vccd1 vccd1 net1102 sky130_fd_sc_hd__buf_2
Xfanout1113 _02787_ vssd1 vssd1 vccd1 vccd1 net1113 sky130_fd_sc_hd__buf_2
Xfanout1124 net1127 vssd1 vssd1 vccd1 vccd1 net1124 sky130_fd_sc_hd__buf_4
XFILLER_0_100_682 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1135 net1136 vssd1 vssd1 vccd1 vccd1 net1135 sky130_fd_sc_hd__buf_4
Xfanout1146 net1147 vssd1 vssd1 vccd1 vccd1 net1146 sky130_fd_sc_hd__clkbuf_8
X_14982_ clknet_leaf_66_wb_clk_i net61 _01347_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12099__A2 net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1157 net1159 vssd1 vssd1 vccd1 vccd1 net1157 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06970__A1 _02871_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1168 net1169 vssd1 vssd1 vccd1 vccd1 net1168 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_35_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1179 net1180 vssd1 vssd1 vccd1 vccd1 net1179 sky130_fd_sc_hd__buf_2
XANTENNA__06970__B2 _02869_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13933_ clknet_leaf_187_wb_clk_i _01697_ _00298_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[287\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10401__A net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13864_ clknet_leaf_7_wb_clk_i _01628_ _00229_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[218\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08078__A net1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12815_ net1394 vssd1 vssd1 vccd1 vccd1 _00579_ sky130_fd_sc_hd__inv_2
XFILLER_0_158_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_83_2076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13795_ clknet_leaf_35_wb_clk_i _01559_ _00160_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[149\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_2087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11931__S net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_159 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12746_ net1286 vssd1 vssd1 vccd1 vccd1 _00510_ sky130_fd_sc_hd__inv_2
XFILLER_0_155_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_173_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_170 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_168 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12677_ net1355 vssd1 vssd1 vccd1 vccd1 _00441_ sky130_fd_sc_hd__inv_2
XFILLER_0_25_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_13_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_3110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14416_ clknet_leaf_161_wb_clk_i _02180_ _00781_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[770\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08227__A1 net1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11628_ _06702_ net383 net348 net2316 vssd1 vssd1 vccd1 vccd1 _01904_ sky130_fd_sc_hd__a22o_1
XFILLER_0_4_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10034__A1 net23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11231__A0 _06545_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14347_ clknet_leaf_34_wb_clk_i _02111_ _00712_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[701\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_672 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11559_ net653 _06669_ vssd1 vssd1 vccd1 vccd1 _06794_ sky130_fd_sc_hd__nor2_1
Xhold607 team_03_WB.instance_to_wrap.core.register_file.registers_state\[866\] vssd1
+ vssd1 vccd1 vccd1 net2100 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10585__A2 net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwire593 _02989_ vssd1 vssd1 vccd1 vccd1 net593 sky130_fd_sc_hd__buf_4
Xhold618 team_03_WB.instance_to_wrap.core.register_file.registers_state\[42\] vssd1
+ vssd1 vccd1 vccd1 net2111 sky130_fd_sc_hd__dlygate4sd3_1
Xhold629 team_03_WB.instance_to_wrap.core.register_file.registers_state\[447\] vssd1
+ vssd1 vccd1 vccd1 net2122 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07450__A2 net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14278_ clknet_leaf_117_wb_clk_i _02042_ _00643_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[632\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_110_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_750 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13229_ net1292 vssd1 vssd1 vccd1 vccd1 _00993_ sky130_fd_sc_hd__inv_2
XANTENNA__08134__B_N _03489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_4_6__f_wb_clk_i clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_6__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
X_08770_ net434 net429 _04711_ vssd1 vssd1 vccd1 vccd1 _04712_ sky130_fd_sc_hd__or3_2
XFILLER_0_58_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09372__A _04382_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14986__Q team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[5\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07721_ net1122 _03661_ _03662_ vssd1 vssd1 vccd1 vccd1 _03663_ sky130_fd_sc_hd__nor3_1
XANTENNA__11298__B1 net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11837__A2 _06675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08163__B1 net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_2533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07652_ net1094 team_03_WB.instance_to_wrap.core.register_file.registers_state\[846\]
+ net798 team_03_WB.instance_to_wrap.core.register_file.registers_state\[878\] net1154
+ vssd1 vssd1 vccd1 vccd1 _03594_ sky130_fd_sc_hd__a221oi_1
XTAP_TAPCELL_ROW_0_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_157_3600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11126__B net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07583_ net1148 _03514_ _03524_ net722 vssd1 vssd1 vccd1 vccd1 _03525_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_76_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09322_ _04711_ _05255_ vssd1 vssd1 vccd1 vccd1 _05264_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_122_2880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_122_2891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08466__A1 net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06935__S net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07958__A1_N net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10965__B _06545_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_153_3508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_861 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_153_3519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09253_ _03604_ _05194_ vssd1 vssd1 vccd1 vccd1 _05195_ sky130_fd_sc_hd__xnor2_1
XANTENNA__11470__B1 net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07674__C1 net1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08204_ net872 _04137_ _04140_ vssd1 vssd1 vccd1 vccd1 _04146_ sky130_fd_sc_hd__or3_1
X_09184_ net579 net572 _05124_ vssd1 vssd1 vccd1 vccd1 _05126_ sky130_fd_sc_hd__and3_2
XFILLER_0_8_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12014__A2 net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_170_3855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_544 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_170_3866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08135_ _03641_ _03823_ _04031_ _04071_ vssd1 vssd1 vccd1 vccd1 _04077_ sky130_fd_sc_hd__and4_1
XANTENNA__10576__A2 net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11773__A1 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07977__B1 net1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1239_A net1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08066_ net1090 team_03_WB.instance_to_wrap.core.register_file.registers_state\[630\]
+ net894 vssd1 vssd1 vccd1 vccd1 _04008_ sky130_fd_sc_hd__or3_1
XFILLER_0_70_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07017_ net1133 _02956_ _02957_ _02958_ vssd1 vssd1 vccd1 vccd1 _02959_ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout699_A net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_794 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07729__B1 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08926__C1 net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11525__B2 net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07067__A net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10879__A3 net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout487_X net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08968_ net1242 team_03_WB.instance_to_wrap.core.register_file.registers_state\[713\]
+ net984 team_03_WB.instance_to_wrap.core.register_file.registers_state\[745\] net944
+ vssd1 vssd1 vccd1 vccd1 _04910_ sky130_fd_sc_hd__o221a_1
X_07919_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[783\] net781
+ _03860_ vssd1 vssd1 vccd1 vccd1 _03861_ sky130_fd_sc_hd__a21o_1
XFILLER_0_98_503 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11828__A2 net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08899_ net857 _04839_ _04840_ _04838_ vssd1 vssd1 vccd1 vccd1 _04841_ sky130_fd_sc_hd__o31a_1
XANTENNA_fanout1396_X net1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10930_ net692 _06515_ _06516_ _06514_ vssd1 vssd1 vccd1 vccd1 _06517_ sky130_fd_sc_hd__a31o_4
Xclkbuf_leaf_92_wb_clk_i clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_92_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_98_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10500__A2 net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07901__B1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10861_ net1248 _06388_ _06459_ vssd1 vssd1 vccd1 vccd1 _06460_ sky130_fd_sc_hd__o21a_1
Xclkbuf_leaf_21_wb_clk_i clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_21_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout821_X net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09103__C1 net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout919_X net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12600_ net1379 vssd1 vssd1 vccd1 vccd1 _00364_ sky130_fd_sc_hd__inv_2
XANTENNA__08457__A1 net1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13580_ net1426 vssd1 vssd1 vccd1 vccd1 _01344_ sky130_fd_sc_hd__inv_2
XFILLER_0_151_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09654__B1 _05595_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10792_ net685 net313 vssd1 vssd1 vccd1 vccd1 _06402_ sky130_fd_sc_hd__nand2_1
XFILLER_0_38_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_1136 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12531_ net1260 vssd1 vssd1 vccd1 vccd1 _00295_ sky130_fd_sc_hd__inv_2
XANTENNA__10803__A3 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_164_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12462_ net1269 vssd1 vssd1 vccd1 vccd1 _00226_ sky130_fd_sc_hd__inv_2
XFILLER_0_151_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_152_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_538 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14201_ clknet_leaf_169_wb_clk_i _01965_ _00566_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[555\]
+ sky130_fd_sc_hd__dfrtp_1
X_11413_ _06478_ _06751_ vssd1 vssd1 vccd1 vccd1 _06753_ sky130_fd_sc_hd__nor2_1
XFILLER_0_152_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12393_ net1254 vssd1 vssd1 vccd1 vccd1 _00157_ sky130_fd_sc_hd__inv_2
XFILLER_0_35_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10567__A2 net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07968__B1 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14132_ clknet_leaf_133_wb_clk_i _01896_ _00497_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[486\]
+ sky130_fd_sc_hd__dfrtp_1
X_11344_ net498 net626 _06724_ net401 net2108 vssd1 vssd1 vccd1 vccd1 _02108_ sky130_fd_sc_hd__a32o_1
XFILLER_0_162_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_284 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14063_ clknet_leaf_135_wb_clk_i _01827_ _00428_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[417\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_120_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11275_ net713 _06504_ net828 vssd1 vssd1 vccd1 vccd1 _06705_ sky130_fd_sc_hd__and3_1
XFILLER_0_120_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_37_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_148_Right_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09744__X _05686_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13014_ net1259 vssd1 vssd1 vccd1 vccd1 _00778_ sky130_fd_sc_hd__inv_2
X_10226_ _06006_ _06067_ vssd1 vssd1 vccd1 vccd1 _06068_ sky130_fd_sc_hd__or2_1
XANTENNA__07196__A1 net1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08393__B1 net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11926__S net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10157_ _03943_ _05998_ vssd1 vssd1 vccd1 vccd1 _05999_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_33_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4 team_03_WB.instance_to_wrap.core.register_file.registers_state\[945\] vssd1
+ vssd1 vccd1 vccd1 net1497 sky130_fd_sc_hd__dlygate4sd3_1
X_10088_ net594 _05456_ _05457_ _05478_ _05499_ vssd1 vssd1 vccd1 vccd1 _05932_ sky130_fd_sc_hd__o311a_1
X_14965_ clknet_leaf_101_wb_clk_i _02717_ _01330_ vssd1 vssd1 vccd1 vccd1 net217 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_85_2116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11819__A2 net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13916_ clknet_leaf_157_wb_clk_i _01680_ _00281_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[270\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_50_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10131__A _03313_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07043__S1 net1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14896_ clknet_leaf_64_wb_clk_i _02659_ _01261_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.pc.current_pc\[25\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__09893__B1 net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15055__1441 vssd1 vssd1 vccd1 vccd1 _15055__1441/HI net1441 sky130_fd_sc_hd__conb_1
XFILLER_0_89_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_159_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_18_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13847_ clknet_leaf_114_wb_clk_i _01611_ _00212_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[201\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_18_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11661__S net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08448__A1 net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13778_ clknet_leaf_118_wb_clk_i _01542_ _00143_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[132\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_100_2430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_174_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_3_0_0_wb_clk_i_X clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12729_ net1357 vssd1 vssd1 vccd1 vccd1 _00493_ sky130_fd_sc_hd__inv_2
XANTENNA__07120__A1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_143_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11204__A0 _06426_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_142_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10558__A2 net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07959__B1 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11755__A1 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold404 team_03_WB.instance_to_wrap.core.register_file.registers_state\[410\] vssd1
+ vssd1 vccd1 vccd1 net1897 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1023 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold415 team_03_WB.instance_to_wrap.core.register_file.registers_state\[185\] vssd1
+ vssd1 vccd1 vccd1 net1908 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold426 team_03_WB.instance_to_wrap.core.register_file.registers_state\[885\] vssd1
+ vssd1 vccd1 vccd1 net1919 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold437 team_03_WB.instance_to_wrap.core.register_file.registers_state\[820\] vssd1
+ vssd1 vccd1 vccd1 net1930 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold448 team_03_WB.instance_to_wrap.core.register_file.registers_state\[34\] vssd1
+ vssd1 vccd1 vccd1 net1941 sky130_fd_sc_hd__dlygate4sd3_1
X_09940_ _05874_ net2252 net292 vssd1 vssd1 vccd1 vccd1 _02757_ sky130_fd_sc_hd__mux2_1
Xhold459 team_03_WB.instance_to_wrap.core.register_file.registers_state\[402\] vssd1
+ vssd1 vccd1 vccd1 net1952 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07974__A3 net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09654__X _05596_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout906 _06285_ vssd1 vssd1 vccd1 vccd1 net906 sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_115_Right_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09871_ _05198_ _05634_ net595 vssd1 vssd1 vccd1 vccd1 _05813_ sky130_fd_sc_hd__a21o_1
XFILLER_0_111_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout917 net923 vssd1 vssd1 vccd1 vccd1 net917 sky130_fd_sc_hd__buf_4
XANTENNA__07187__A1 net1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout928 net932 vssd1 vssd1 vccd1 vccd1 net928 sky130_fd_sc_hd__buf_4
XFILLER_0_110_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_74_1897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout939 net949 vssd1 vssd1 vccd1 vccd1 net939 sky130_fd_sc_hd__buf_4
XFILLER_0_29_71 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08822_ net1053 team_03_WB.instance_to_wrap.core.register_file.registers_state\[673\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[641\] net1006 net1214
+ vssd1 vssd1 vccd1 vccd1 _04764_ sky130_fd_sc_hd__o221a_1
XANTENNA__08923__A2 net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10740__S net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_146_3367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_146_3378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1104 team_03_WB.instance_to_wrap.core.register_file.registers_state\[85\] vssd1
+ vssd1 vccd1 vccd1 net2597 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06934__A1 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1115 team_03_WB.instance_to_wrap.core.register_file.registers_state\[601\] vssd1
+ vssd1 vccd1 vccd1 net2608 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1126 team_03_WB.instance_to_wrap.core.register_file.registers_state\[719\] vssd1
+ vssd1 vccd1 vccd1 net2619 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07615__A net1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1137 team_03_WB.instance_to_wrap.core.register_file.registers_state\[468\] vssd1
+ vssd1 vccd1 vccd1 net2630 sky130_fd_sc_hd__dlygate4sd3_1
X_08753_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[547\] net980
+ vssd1 vssd1 vccd1 vccd1 _04695_ sky130_fd_sc_hd__or2_1
Xhold1148 team_03_WB.instance_to_wrap.core.register_file.registers_state\[77\] vssd1
+ vssd1 vccd1 vccd1 net2641 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1159 team_03_WB.instance_to_wrap.core.register_file.registers_state\[5\] vssd1
+ vssd1 vccd1 vccd1 net2652 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_124_2920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_124_2931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07704_ net747 _03642_ _03643_ _03644_ _03645_ vssd1 vssd1 vccd1 vccd1 _03646_ sky130_fd_sc_hd__o32a_1
X_08684_ _04622_ _04623_ _04624_ _04625_ net862 net924 vssd1 vssd1 vccd1 vccd1 _04626_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__09884__B1 net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07635_ net809 _03572_ _03575_ _03576_ vssd1 vssd1 vccd1 vccd1 _03577_ sky130_fd_sc_hd__a22o_1
XANTENNA__11691__B1 net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07895__C1 net1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1091_A net1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_2839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout447_A _06801_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1189_A net1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08439__A1 net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07566_ net1188 team_03_WB.instance_to_wrap.core.register_file.registers_state\[728\]
+ net781 team_03_WB.instance_to_wrap.core.register_file.registers_state\[760\] net745
+ vssd1 vssd1 vccd1 vccd1 _03508_ sky130_fd_sc_hd__o221a_1
XFILLER_0_165_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_172_3906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09305_ net609 _05144_ vssd1 vssd1 vccd1 vccd1 _05247_ sky130_fd_sc_hd__nor2_1
XFILLER_0_76_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07647__C1 net1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10187__S net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_628 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout614_A net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07497_ _03437_ _03438_ vssd1 vssd1 vccd1 vccd1 _03439_ sky130_fd_sc_hd__and2_1
XANTENNA__09976__S net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09236_ _05176_ _05177_ vssd1 vssd1 vccd1 vccd1 _05178_ sky130_fd_sc_hd__and2b_1
XFILLER_0_63_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07662__A2 _03600_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_17_Right_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09167_ net436 net428 _04953_ net552 vssd1 vssd1 vccd1 vccd1 _05109_ sky130_fd_sc_hd__o31a_1
XFILLER_0_134_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout402_X net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1144_X net1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08118_ net1181 team_03_WB.instance_to_wrap.core.register_file.registers_state\[986\]
+ vssd1 vssd1 vccd1 vccd1 _04060_ sky130_fd_sc_hd__or2_1
XFILLER_0_161_699 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_571 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09098_ net868 _05039_ _05034_ net852 vssd1 vssd1 vccd1 vccd1 _05040_ sky130_fd_sc_hd__o211a_1
XFILLER_0_82_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout983_A net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08049_ net1186 team_03_WB.instance_to_wrap.core.register_file.registers_state\[54\]
+ net879 vssd1 vssd1 vccd1 vccd1 _03991_ sky130_fd_sc_hd__and3_1
Xhold960 team_03_WB.instance_to_wrap.core.register_file.registers_state\[326\] vssd1
+ vssd1 vccd1 vccd1 net2453 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold971 team_03_WB.instance_to_wrap.core.register_file.registers_state\[920\] vssd1
+ vssd1 vccd1 vccd1 net2464 sky130_fd_sc_hd__dlygate4sd3_1
X_11060_ net2530 net422 _06607_ net510 vssd1 vssd1 vccd1 vccd1 _02275_ sky130_fd_sc_hd__a22o_1
Xhold982 team_03_WB.instance_to_wrap.core.register_file.registers_state\[745\] vssd1
+ vssd1 vccd1 vccd1 net2475 sky130_fd_sc_hd__dlygate4sd3_1
Xhold993 team_03_WB.instance_to_wrap.core.register_file.registers_state\[469\] vssd1
+ vssd1 vccd1 vccd1 net2486 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout771_X net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout869_X net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10011_ _03023_ net1672 net287 vssd1 vssd1 vccd1 vccd1 _02703_ sky130_fd_sc_hd__mux2_1
XANTENNA__13527__A net1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10650__S net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_26_Right_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_4_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1106 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11047__A net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14750_ clknet_leaf_50_wb_clk_i _02514_ _01115_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_169_711 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11962_ net633 _06739_ net466 net365 net2143 vssd1 vssd1 vccd1 vccd1 _01581_ sky130_fd_sc_hd__a32o_1
XFILLER_0_153_1128 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09875__B1 _03601_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13701_ clknet_leaf_14_wb_clk_i _01465_ _00066_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[55\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_168_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10913_ net693 _06501_ _06502_ _06500_ vssd1 vssd1 vccd1 vccd1 _06503_ sky130_fd_sc_hd__a31o_4
X_14681_ clknet_leaf_81_wb_clk_i _02445_ _01046_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.ADR_I\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11682__B1 net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11893_ net634 _06702_ net465 net373 net2031 vssd1 vssd1 vccd1 vccd1 _01648_ sky130_fd_sc_hd__a32o_1
XANTENNA__07350__A1 net1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_2013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13632_ net1433 vssd1 vssd1 vccd1 vccd1 _01396_ sky130_fd_sc_hd__inv_2
XFILLER_0_156_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10844_ team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[21\] net307 net685 vssd1
+ vssd1 vccd1 vccd1 _06444_ sky130_fd_sc_hd__a21o_1
XFILLER_0_67_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11434__A0 _06557_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13563_ net1427 vssd1 vssd1 vccd1 vccd1 _01327_ sky130_fd_sc_hd__inv_2
X_10775_ _02930_ _06384_ _06383_ _02942_ _02934_ vssd1 vssd1 vccd1 vccd1 _06385_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_87_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_35_Right_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12514_ net1296 vssd1 vssd1 vccd1 vccd1 _00278_ sky130_fd_sc_hd__inv_2
XANTENNA__08790__S net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13494_ net1328 vssd1 vssd1 vccd1 vccd1 _01258_ sky130_fd_sc_hd__inv_2
XFILLER_0_81_244 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12445_ net1388 vssd1 vssd1 vccd1 vccd1 _00209_ sky130_fd_sc_hd__inv_2
XFILLER_0_81_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11737__A1 net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08602__A1 net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08063__C1 net1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12376_ net1374 vssd1 vssd1 vccd1 vccd1 _00140_ sky130_fd_sc_hd__inv_2
XANTENNA__08091__A net1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14115_ clknet_leaf_35_wb_clk_i _01879_ _00480_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[469\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11327_ net264 net2690 net404 vssd1 vssd1 vccd1 vccd1 _02118_ sky130_fd_sc_hd__mux2_1
X_15095_ net1481 vssd1 vssd1 vccd1 vccd1 la_data_out[31] sky130_fd_sc_hd__buf_2
XANTENNA__10126__A _03279_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_574 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09915__A _05646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14046_ clknet_leaf_119_wb_clk_i _01810_ _00411_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[400\]
+ sky130_fd_sc_hd__dfrtp_1
X_11258_ net493 net622 _06696_ net408 net2250 vssd1 vssd1 vccd1 vccd1 _02166_ sky130_fd_sc_hd__a32o_1
XFILLER_0_5_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_44_Right_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11656__S net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10209_ _06043_ _06050_ _06042_ vssd1 vssd1 vccd1 vccd1 _06051_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_52_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10173__A0 _04954_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11189_ net505 net654 _06675_ net414 net1918 vssd1 vssd1 vccd1 vccd1 _02214_ sky130_fd_sc_hd__a32o_1
XANTENNA__10712__A2 net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14948_ clknet_leaf_55_wb_clk_i _02700_ _01313_ vssd1 vssd1 vccd1 vccd1 team_03_WB.EN_VAL_REG
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_141_3264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_141_3275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07877__C1 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14879_ clknet_leaf_84_wb_clk_i _02642_ _01244_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.pc.current_pc\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_77_528 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07341__A1 net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07420_ _03355_ _03356_ _03361_ net1161 vssd1 vssd1 vccd1 vccd1 _03362_ sky130_fd_sc_hd__o22a_1
XFILLER_0_58_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_53_Right_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07629__C1 net1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07351_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[444\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[412\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[316\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[284\]
+ net757 net1123 vssd1 vssd1 vccd1 vccd1 _03293_ sky130_fd_sc_hd__mux4_1
XFILLER_0_70_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_414 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09633__A3 _05570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_211 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07282_ net823 _03222_ _03223_ vssd1 vssd1 vccd1 vccd1 _03224_ sky130_fd_sc_hd__or3_1
XFILLER_0_143_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10087__A_N _05686_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_324 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09021_ net1244 team_03_WB.instance_to_wrap.core.register_file.registers_state\[208\]
+ net989 team_03_WB.instance_to_wrap.core.register_file.registers_state\[240\] net944
+ vssd1 vssd1 vccd1 vccd1 _04963_ sky130_fd_sc_hd__o221a_1
XFILLER_0_116_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11728__A1 _06491_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11420__A _06503_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08054__C1 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold201 team_03_WB.instance_to_wrap.core.register_file.registers_state\[14\] vssd1
+ vssd1 vccd1 vccd1 net1694 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold212 team_03_WB.instance_to_wrap.core.register_file.registers_state\[565\] vssd1
+ vssd1 vccd1 vccd1 net1705 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_76_1937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold223 team_03_WB.instance_to_wrap.CPU_DAT_I\[24\] vssd1 vssd1 vccd1 vccd1 net1716
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_76_1948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold234 team_03_WB.instance_to_wrap.core.register_file.registers_state\[998\] vssd1
+ vssd1 vccd1 vccd1 net1727 sky130_fd_sc_hd__dlygate4sd3_1
Xhold245 net224 vssd1 vssd1 vccd1 vccd1 net1738 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_148_3407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_148_3418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold256 team_03_WB.instance_to_wrap.core.register_file.registers_state\[913\] vssd1
+ vssd1 vccd1 vccd1 net1749 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_62_Right_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold267 net202 vssd1 vssd1 vccd1 vccd1 net1760 sky130_fd_sc_hd__dlygate4sd3_1
Xhold278 net178 vssd1 vssd1 vccd1 vccd1 net1771 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_113_2687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09923_ _05863_ _05864_ net311 _05429_ vssd1 vssd1 vccd1 vccd1 _05865_ sky130_fd_sc_hd__and4bb_1
XTAP_TAPCELL_ROW_113_2698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold289 team_03_WB.instance_to_wrap.CPU_DAT_I\[10\] vssd1 vssd1 vccd1 vccd1 net1782
+ sky130_fd_sc_hd__dlygate4sd3_1
Xfanout703 net704 vssd1 vssd1 vccd1 vccd1 net703 sky130_fd_sc_hd__buf_4
Xfanout714 net716 vssd1 vssd1 vccd1 vccd1 net714 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_165_3754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout725 net727 vssd1 vssd1 vccd1 vccd1 net725 sky130_fd_sc_hd__buf_4
XANTENNA_fanout397_A _06752_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_165_3765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13347__A net1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout736 net737 vssd1 vssd1 vccd1 vccd1 net736 sky130_fd_sc_hd__buf_2
X_09854_ net565 _05792_ _05793_ net579 vssd1 vssd1 vccd1 vccd1 _05796_ sky130_fd_sc_hd__o31a_1
Xfanout747 net748 vssd1 vssd1 vccd1 vccd1 net747 sky130_fd_sc_hd__buf_4
Xfanout758 net761 vssd1 vssd1 vccd1 vccd1 net758 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout1104_A net1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout769 net770 vssd1 vssd1 vccd1 vccd1 net769 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11900__A1 net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09036__S net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07345__A net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08805_ net863 _04745_ _04746_ vssd1 vssd1 vccd1 vccd1 _04747_ sky130_fd_sc_hd__and3_1
X_09785_ _03459_ _04619_ _04820_ _05726_ vssd1 vssd1 vccd1 vccd1 _05727_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout564_A _03025_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06997_ _02927_ _02929_ vssd1 vssd1 vccd1 vccd1 _02939_ sky130_fd_sc_hd__or2_1
XANTENNA__08109__B1 net1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_0_Left_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_1_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08736_ net1081 _04670_ _04677_ net848 vssd1 vssd1 vccd1 vccd1 _04678_ sky130_fd_sc_hd__a211o_1
XANTENNA__07868__C1 net1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout731_A net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08667_ net1058 team_03_WB.instance_to_wrap.core.register_file.registers_state\[967\]
+ net1011 team_03_WB.instance_to_wrap.core.register_file.registers_state\[999\] net1080
+ vssd1 vssd1 vccd1 vccd1 _04609_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout352_X net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07332__A1 net1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1094_X net1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout829_A net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_71_Right_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07618_ _03558_ _03559_ net814 vssd1 vssd1 vccd1 vccd1 _03560_ sky130_fd_sc_hd__a21o_1
X_08598_ net1058 team_03_WB.instance_to_wrap.core.register_file.registers_state\[709\]
+ net1011 team_03_WB.instance_to_wrap.core.register_file.registers_state\[741\] net931
+ vssd1 vssd1 vccd1 vccd1 _04540_ sky130_fd_sc_hd__a221o_1
XANTENNA__07883__A2 net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11416__A0 net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07549_ _03459_ _03489_ vssd1 vssd1 vccd1 vccd1 _03491_ sky130_fd_sc_hd__nor2_1
XFILLER_0_49_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout617_X net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11967__A1 net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_211 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10560_ net1876 net531 net598 _05870_ vssd1 vssd1 vccd1 vccd1 _02563_ sky130_fd_sc_hd__a22o_1
X_09219_ net607 _05160_ vssd1 vssd1 vccd1 vccd1 _05161_ sky130_fd_sc_hd__nor2_1
XFILLER_0_161_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_132 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10645__S net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10491_ net109 net1029 net906 net1803 vssd1 vssd1 vccd1 vccd1 _02618_ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_21_wb_clk_i_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11719__A1 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12230_ net1540 vssd1 vssd1 vccd1 vccd1 _01427_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_20_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08045__C1 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_20_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_130 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout986_X net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07399__A1 net1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15054__1440 vssd1 vssd1 vccd1 vccd1 _15054__1440/HI net1440 sky130_fd_sc_hd__conb_1
XANTENNA__11195__A2 net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_80_Right_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12161_ net1506 vssd1 vssd1 vccd1 vccd1 _02392_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07954__S net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11112_ net264 net2640 net418 vssd1 vssd1 vccd1 vccd1 _02246_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12092_ _06790_ net469 net441 net1920 vssd1 vssd1 vccd1 vccd1 _01455_ sky130_fd_sc_hd__a22o_1
Xhold790 team_03_WB.instance_to_wrap.core.register_file.registers_state\[655\] vssd1
+ vssd1 vccd1 vccd1 net2283 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_120_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11043_ net710 _06517_ net701 vssd1 vssd1 vccd1 vccd1 _06598_ sky130_fd_sc_hd__or3_1
XANTENNA__08899__A1 net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07571__A1 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14802_ clknet_leaf_92_wb_clk_i _02566_ _01167_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_I\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_157_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12994_ net1352 vssd1 vssd1 vccd1 vccd1 _00758_ sky130_fd_sc_hd__inv_2
XFILLER_0_98_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14733_ clknet_leaf_48_wb_clk_i _02497_ _01098_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.decoder.inst\[30\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_59_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11945_ net619 _06722_ net452 net363 net2432 vssd1 vssd1 vccd1 vccd1 _01598_ sky130_fd_sc_hd__a32o_1
XANTENNA_output114_A net114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11064__X _06610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14664_ clknet_leaf_10_wb_clk_i _02428_ _01029_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1018\]
+ sky130_fd_sc_hd__dfstp_1
X_11876_ net621 _06685_ net453 net371 net2050 vssd1 vssd1 vccd1 vccd1 _01665_ sky130_fd_sc_hd__a32o_1
XANTENNA_clkbuf_leaf_60_wb_clk_i_A clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_55_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11407__A0 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13615_ net1422 vssd1 vssd1 vccd1 vccd1 _01379_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10827_ net277 net2400 net521 vssd1 vssd1 vccd1 vccd1 _02331_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11224__B _06517_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09076__A1 net1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14595_ clknet_leaf_47_wb_clk_i _02359_ _00960_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[949\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_27_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11958__A1 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13546_ net1324 vssd1 vssd1 vccd1 vccd1 _01310_ sky130_fd_sc_hd__inv_2
XANTENNA__12080__B1 net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10758_ net1638 net529 net524 _06372_ vssd1 vssd1 vccd1 vccd1 _02438_ sky130_fd_sc_hd__a22o_1
XFILLER_0_137_471 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08823__A1 net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13477_ net1431 vssd1 vssd1 vccd1 vccd1 _01241_ sky130_fd_sc_hd__inv_2
XANTENNA__09629__B _04415_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_97_2362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10689_ _05563_ _06312_ vssd1 vssd1 vccd1 vccd1 _06329_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_97_2373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12428_ net1331 vssd1 vssd1 vccd1 vccd1 _00192_ sky130_fd_sc_hd__inv_2
XFILLER_0_50_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_168_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12359_ net1368 vssd1 vssd1 vccd1 vccd1 _00123_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10933__A2 net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15078_ net1464 vssd1 vssd1 vccd1 vccd1 la_data_out[14] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_71_1834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13167__A net1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14029_ clknet_leaf_187_wb_clk_i _01793_ _00394_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[383\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_71_1845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06920_ _02858_ _02861_ net819 vssd1 vssd1 vccd1 vccd1 _02862_ sky130_fd_sc_hd__o21a_1
XANTENNA__09000__A1 net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_143_3304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_3315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10697__B2 net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06851_ team_03_WB.instance_to_wrap.core.control_logic.instruction\[4\] vssd1 vssd1
+ vccd1 vccd1 _02794_ sky130_fd_sc_hd__inv_2
XANTENNA__11894__B1 net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_160_3651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09570_ net320 _05378_ _05510_ _05511_ vssd1 vssd1 vccd1 vccd1 _05512_ sky130_fd_sc_hd__a211o_1
XFILLER_0_171_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_160_3662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1134 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08521_ net1230 team_03_WB.instance_to_wrap.core.register_file.registers_state\[191\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[159\] net959 net916
+ vssd1 vssd1 vccd1 vccd1 _04463_ sky130_fd_sc_hd__a221o_1
XANTENNA__14994__Q team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[13\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_69_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08511__B1 net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_149_wb_clk_i clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_149_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_69_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08452_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[956\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[924\]
+ net953 vssd1 vssd1 vccd1 vccd1 _04394_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07403_ net1082 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1023\]
+ net888 _03344_ net1149 vssd1 vssd1 vccd1 vccd1 _03345_ sky130_fd_sc_hd__o311a_1
XFILLER_0_58_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11134__B net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08383_ net432 net424 _04323_ net542 vssd1 vssd1 vccd1 vccd1 _04325_ sky130_fd_sc_hd__o31a_1
XFILLER_0_133_73 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11949__A1 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07078__B1 net1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07334_ net817 _03275_ net717 vssd1 vssd1 vccd1 vccd1 _03276_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_73_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10973__B net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_789 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10621__A1 team_03_WB.instance_to_wrap.CPU_DAT_O\[8\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_07265_ net615 _03206_ vssd1 vssd1 vccd1 vccd1 _03207_ sky130_fd_sc_hd__or2_1
XFILLER_0_33_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout312_A _05388_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1054_A net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11150__A net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09004_ net1045 team_03_WB.instance_to_wrap.core.register_file.registers_state\[714\]
+ net995 team_03_WB.instance_to_wrap.core.register_file.registers_state\[746\] net916
+ vssd1 vssd1 vccd1 vccd1 _04946_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_115_2738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07196_ net1207 net1015 _03107_ vssd1 vssd1 vccd1 vccd1 _03138_ sky130_fd_sc_hd__a21o_2
XFILLER_0_131_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11177__A2 net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08578__B1 net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_167_3805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1221_A net1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_105_wb_clk_i_A clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__07250__B1 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_894 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout681_A _05915_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout500 net517 vssd1 vssd1 vccd1 vccd1 net500 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_6_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout779_A net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout511 net513 vssd1 vssd1 vccd1 vccd1 net511 sky130_fd_sc_hd__clkbuf_4
Xfanout522 _06322_ vssd1 vssd1 vccd1 vccd1 net522 sky130_fd_sc_hd__clkbuf_4
X_09906_ _05596_ _05833_ _05847_ _05500_ vssd1 vssd1 vccd1 vccd1 _05848_ sky130_fd_sc_hd__or4b_1
Xfanout533 _06298_ vssd1 vssd1 vccd1 vccd1 net533 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_158_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout544 net545 vssd1 vssd1 vccd1 vccd1 net544 sky130_fd_sc_hd__buf_2
XANTENNA_fanout1107_X net1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout555 net558 vssd1 vssd1 vccd1 vccd1 net555 sky130_fd_sc_hd__buf_4
XANTENNA__10688__A1 net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout566 _03025_ vssd1 vssd1 vccd1 vccd1 net566 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09842__X _05784_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09837_ net566 _05721_ vssd1 vssd1 vccd1 vccd1 _05779_ sky130_fd_sc_hd__nand2_1
Xfanout577 _02993_ vssd1 vssd1 vccd1 vccd1 net577 sky130_fd_sc_hd__buf_2
XANTENNA__11885__B1 net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout599 net600 vssd1 vssd1 vccd1 vccd1 net599 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout946_A net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09768_ _05092_ _05120_ net578 vssd1 vssd1 vccd1 vccd1 _05710_ sky130_fd_sc_hd__mux2_1
X_08719_ net1223 _04658_ _04659_ vssd1 vssd1 vccd1 vccd1 _04661_ sky130_fd_sc_hd__and3_1
XANTENNA__11637__B1 net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09699_ _04816_ _05639_ net664 vssd1 vssd1 vccd1 vccd1 _05641_ sky130_fd_sc_hd__o21a_1
XANTENNA__07305__A1 net1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout734_X net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11730_ net1910 net297 net336 vssd1 vssd1 vccd1 vccd1 _01806_ sky130_fd_sc_hd__mux2_1
XANTENNA__07856__A2 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11661_ net2064 _06624_ net344 vssd1 vssd1 vccd1 vccd1 _01872_ sky130_fd_sc_hd__mux2_1
XANTENNA__07241__C net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09058__A1 net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout901_X net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13400_ net1424 vssd1 vssd1 vccd1 vccd1 _01164_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_25_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10612_ net2218 team_03_WB.instance_to_wrap.CPU_DAT_O\[17\] net841 vssd1 vssd1 vccd1
+ vccd1 _02516_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_25_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07069__B1 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_54_Left_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14380_ clknet_leaf_16_wb_clk_i _02144_ _00745_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[734\]
+ sky130_fd_sc_hd__dfrtp_1
X_11592_ net299 net2419 net448 vssd1 vssd1 vccd1 vccd1 _01937_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_929 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10883__B _06478_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_144_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_13331_ net1326 vssd1 vssd1 vccd1 vccd1 _01095_ sky130_fd_sc_hd__inv_2
XFILLER_0_146_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10612__A1 team_03_WB.instance_to_wrap.CPU_DAT_O\[17\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10543_ net2427 net1030 net908 vssd1 vssd1 vccd1 vccd1 _02568_ sky130_fd_sc_hd__a21o_1
XFILLER_0_52_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_1135 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_150_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08018__C1 net1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input75_A wbs_adr_i[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13262_ net1303 vssd1 vssd1 vccd1 vccd1 _01026_ sky130_fd_sc_hd__inv_2
X_10474_ net1 net1027 vssd1 vssd1 vccd1 vccd1 _06285_ sky130_fd_sc_hd__nor2_4
XTAP_TAPCELL_ROW_40_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08072__C net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15001_ clknet_leaf_40_wb_clk_i net49 _01366_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_12213_ net1566 vssd1 vssd1 vccd1 vccd1 _02340_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_122_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13193_ net1256 vssd1 vssd1 vccd1 vccd1 _00957_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_92_2270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12144_ net1570 vssd1 vssd1 vccd1 vccd1 _02409_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_138_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09184__B net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_63_Left_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10128__B1 _03279_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12075_ _06781_ net452 net439 net1944 vssd1 vssd1 vccd1 vccd1 _01472_ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_1032 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input30_X net30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09533__A2 _04354_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11026_ net2607 net421 _06587_ net502 vssd1 vssd1 vccd1 vccd1 _02289_ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11876__B1 net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10898__X _06491_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07416__C net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1087 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08741__B1 net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11340__A2 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07544__B2 net1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11934__S net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09912__B _05730_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11891__A3 net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07713__A net1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11628__B1 net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12977_ net1268 vssd1 vssd1 vccd1 vccd1 _00741_ sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_183_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11235__A _06405_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14716_ clknet_leaf_62_wb_clk_i _02480_ _01081_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.decoder.inst\[13\]
+ sky130_fd_sc_hd__dfrtp_4
X_11928_ _06626_ net2724 net369 vssd1 vssd1 vccd1 vccd1 _01614_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_47_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_47_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_72_Left_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_170_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14647_ clknet_leaf_110_wb_clk_i _02411_ _01012_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1001\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__09049__A1 net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_2402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11859_ _06487_ net2211 net376 vssd1 vssd1 vccd1 vccd1 _01681_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_99_2413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_64_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08257__C1 net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14578_ clknet_leaf_160_wb_clk_i _02342_ _00943_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[932\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__10793__B _05867_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08544__A net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_3163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_3174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13529_ net1316 vssd1 vssd1 vccd1 vccd1 _01293_ sky130_fd_sc_hd__inv_2
XFILLER_0_103_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_153_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07050_ net614 net593 _02991_ vssd1 vssd1 vccd1 vccd1 _02992_ sky130_fd_sc_hd__a21o_2
XFILLER_0_153_794 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07480__B1 net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput103 net103 vssd1 vssd1 vccd1 vccd1 ADR_O[0] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_11_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput114 net114 vssd1 vssd1 vccd1 vccd1 ADR_O[1] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_23_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput125 net125 vssd1 vssd1 vccd1 vccd1 ADR_O[2] sky130_fd_sc_hd__clkbuf_4
XANTENNA__06999__A team_03_WB.instance_to_wrap.core.decoder.inst\[13\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput136 net136 vssd1 vssd1 vccd1 vccd1 DAT_O[0] sky130_fd_sc_hd__buf_2
XANTENNA__10906__A2 net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput147 net147 vssd1 vssd1 vccd1 vccd1 DAT_O[1] sky130_fd_sc_hd__buf_2
XFILLER_0_2_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07447__X _03389_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14989__Q team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[8\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_81_Left_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_1100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_2635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput158 net158 vssd1 vssd1 vccd1 vccd1 DAT_O[2] sky130_fd_sc_hd__buf_2
Xoutput169 net169 vssd1 vssd1 vccd1 vccd1 SEL_O[1] sky130_fd_sc_hd__clkbuf_4
X_15117__1487 vssd1 vssd1 vccd1 vccd1 _15117__1487/HI net1487 sky130_fd_sc_hd__conb_1
XFILLER_0_103_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_162_3702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12005__S net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07952_ net1147 _03884_ _03885_ _03893_ net1162 vssd1 vssd1 vccd1 vccd1 _03894_ sky130_fd_sc_hd__o311a_1
X_06903_ net1017 net1015 net1018 vssd1 vssd1 vccd1 vccd1 _02845_ sky130_fd_sc_hd__o21ai_1
XANTENNA__11129__B net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07883_ net1187 net877 team_03_WB.instance_to_wrap.core.register_file.registers_state\[15\]
+ vssd1 vssd1 vccd1 vccd1 _03825_ sky130_fd_sc_hd__a21o_1
XANTENNA__11844__S net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09622_ _05331_ _05335_ _05337_ vssd1 vssd1 vccd1 vccd1 _05564_ sky130_fd_sc_hd__or3_1
X_06834_ team_03_WB.instance_to_wrap.READ_I vssd1 vssd1 vccd1 vccd1 _02777_ sky130_fd_sc_hd__inv_2
XANTENNA__06938__S net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08719__A net1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11882__A3 net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09553_ _05493_ _05494_ net567 vssd1 vssd1 vccd1 vccd1 _05495_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_108_2586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11619__B1 net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_2597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08504_ _04080_ _04444_ vssd1 vssd1 vccd1 vccd1 _04446_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_90_Left_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09484_ _05425_ vssd1 vssd1 vccd1 vccd1 _05426_ sky130_fd_sc_hd__inv_2
XANTENNA__08496__C1 net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08435_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[954\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[922\]
+ net964 vssd1 vssd1 vccd1 vccd1 _04377_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout527_A net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1171_A net1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1269_A net1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08366_ net1219 _04306_ _04307_ vssd1 vssd1 vccd1 vccd1 _04308_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_163_547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07317_ net807 _03247_ _03248_ vssd1 vssd1 vccd1 vccd1 _03259_ sky130_fd_sc_hd__or3_1
XFILLER_0_18_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08297_ net944 _04238_ vssd1 vssd1 vccd1 vccd1 _04239_ sky130_fd_sc_hd__or2_1
XANTENNA__09984__S net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1436_A net1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07471__B1 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07248_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[8\] net774
+ net746 _03189_ vssd1 vssd1 vccd1 vccd1 _03190_ sky130_fd_sc_hd__a211o_1
Xclkbuf_leaf_46_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_46_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_103_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout896_A net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_995 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09556__Y _05498_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09212__A1 _03391_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10358__B1 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07179_ net1161 _03119_ _03120_ vssd1 vssd1 vccd1 vccd1 _03121_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout1224_X net1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_291 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10190_ _06030_ _06031_ vssd1 vssd1 vccd1 vccd1 _06032_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout684_X net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07774__A1 net1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1306 net1309 vssd1 vssd1 vccd1 vccd1 net1306 sky130_fd_sc_hd__buf_4
XFILLER_0_100_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1317 net1320 vssd1 vssd1 vccd1 vccd1 net1317 sky130_fd_sc_hd__buf_4
Xfanout1328 net1329 vssd1 vssd1 vccd1 vccd1 net1328 sky130_fd_sc_hd__buf_4
Xfanout330 _06810_ vssd1 vssd1 vccd1 vccd1 net330 sky130_fd_sc_hd__buf_4
Xfanout341 _06806_ vssd1 vssd1 vccd1 vccd1 net341 sky130_fd_sc_hd__buf_2
Xfanout1339 net1346 vssd1 vssd1 vccd1 vccd1 net1339 sky130_fd_sc_hd__clkbuf_4
Xfanout352 _04776_ vssd1 vssd1 vccd1 vccd1 net352 sky130_fd_sc_hd__buf_4
XANTENNA__11858__A0 _06483_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout363 _06815_ vssd1 vssd1 vccd1 vccd1 net363 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout851_X net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07526__A1 net1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout374 _06813_ vssd1 vssd1 vccd1 vccd1 net374 sky130_fd_sc_hd__clkbuf_4
Xfanout385 net387 vssd1 vssd1 vccd1 vccd1 net385 sky130_fd_sc_hd__buf_4
XANTENNA_fanout949_X net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12900_ net1366 vssd1 vssd1 vccd1 vccd1 _00664_ sky130_fd_sc_hd__inv_2
Xfanout396 _06752_ vssd1 vssd1 vccd1 vccd1 net396 sky130_fd_sc_hd__clkbuf_8
X_13880_ clknet_leaf_185_wb_clk_i _01644_ _00245_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[234\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10530__B1 net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12831_ net1347 vssd1 vssd1 vccd1 vccd1 _00595_ sky130_fd_sc_hd__inv_2
XFILLER_0_115_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11055__A net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12762_ net1372 vssd1 vssd1 vccd1 vccd1 _00526_ sky130_fd_sc_hd__inv_2
XFILLER_0_115_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14501_ clknet_leaf_40_wb_clk_i _02265_ _00866_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[855\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_90_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11713_ net1880 _06413_ net335 vssd1 vssd1 vccd1 vccd1 _01823_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12693_ net1275 vssd1 vssd1 vccd1 vccd1 _00457_ sky130_fd_sc_hd__inv_2
XFILLER_0_49_380 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_166_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14432_ clknet_leaf_2_wb_clk_i _02196_ _00797_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[786\]
+ sky130_fd_sc_hd__dfrtp_1
X_11644_ net2459 _06609_ net342 vssd1 vssd1 vccd1 vccd1 _01889_ sky130_fd_sc_hd__mux2_1
XANTENNA__12035__B1 net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_3_5_0_wb_clk_i_X clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14363_ clknet_leaf_124_wb_clk_i _02127_ _00728_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[717\]
+ sky130_fd_sc_hd__dfrtp_1
X_11575_ _06390_ _06394_ vssd1 vssd1 vccd1 vccd1 _06801_ sky130_fd_sc_hd__nand2_4
Xinput16 DAT_I[22] vssd1 vssd1 vccd1 vccd1 net16 sky130_fd_sc_hd__clkbuf_2
Xinput27 DAT_I[3] vssd1 vssd1 vccd1 vccd1 net27 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_2310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput38 gpio_in[13] vssd1 vssd1 vccd1 vccd1 net38 sky130_fd_sc_hd__clkbuf_1
X_13314_ net1325 vssd1 vssd1 vccd1 vccd1 _01078_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10526_ net140 net1034 net1026 net1718 vssd1 vssd1 vccd1 vccd1 _02584_ sky130_fd_sc_hd__a22o_1
Xinput49 gpio_in[24] vssd1 vssd1 vccd1 vccd1 net49 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_109_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14294_ clknet_leaf_154_wb_clk_i _02058_ _00659_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[648\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11929__S net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_3060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13245_ net1388 vssd1 vssd1 vccd1 vccd1 _01009_ sky130_fd_sc_hd__inv_2
X_10457_ team_03_WB.instance_to_wrap.core.pc.current_pc\[4\] _06134_ vssd1 vssd1 vccd1
+ vccd1 _06272_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_131_3071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_932 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_2218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_2229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_1019 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08411__C1 net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13176_ net1380 vssd1 vssd1 vccd1 vccd1 _00940_ sky130_fd_sc_hd__inv_2
XANTENNA__11010__B2 net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10388_ _05994_ _05995_ _06085_ vssd1 vssd1 vccd1 vccd1 _06216_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07765__A1 net1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08962__B1 net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12127_ net1518 vssd1 vssd1 vccd1 vccd1 _02426_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_4_5__f_wb_clk_i clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_5__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__06973__C1 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11849__A0 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12058_ _06624_ net2399 net357 vssd1 vssd1 vccd1 vccd1 _01488_ sky130_fd_sc_hd__mux2_1
XANTENNA__07517__A1 _03458_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11664__S net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08714__B1 net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11009_ net630 _06577_ vssd1 vssd1 vccd1 vccd1 _06578_ sky130_fd_sc_hd__nor2_1
XANTENNA__10521__B1 net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08539__A net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_66_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08478__C1 net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_3203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_3214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10824__A1 net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_2483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09690__A1 net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_2494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08220_ net1217 _04160_ _04161_ vssd1 vssd1 vccd1 vccd1 _04162_ sky130_fd_sc_hd__o21a_1
XFILLER_0_118_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12026__B1 net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_155_3550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_155_3561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_22 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08151_ net1230 team_03_WB.instance_to_wrap.core.register_file.registers_state\[212\]
+ net960 team_03_WB.instance_to_wrap.core.register_file.registers_state\[244\] net936
+ vssd1 vssd1 vccd1 vccd1 _04093_ sky130_fd_sc_hd__o221a_1
XANTENNA__10588__B1 net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_160_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07102_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[417\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[385\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[289\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[257\]
+ net780 net1133 vssd1 vssd1 vccd1 vccd1 _03044_ sky130_fd_sc_hd__mux4_1
XANTENNA__10052__A2 net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07453__B1 net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_151_3469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08561__X _04503_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08082_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[918\] net793
+ net1014 _04023_ vssd1 vssd1 vccd1 vccd1 _04024_ sky130_fd_sc_hd__o211a_1
XFILLER_0_28_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10028__B net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_141_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07033_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[163\] net780
+ net748 _02974_ vssd1 vssd1 vccd1 vccd1 _02975_ sky130_fd_sc_hd__o211a_1
XFILLER_0_2_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08402__C1 net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07756__A1 net1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08984_ net1232 team_03_WB.instance_to_wrap.core.register_file.registers_state\[138\]
+ net960 team_03_WB.instance_to_wrap.core.register_file.registers_state\[170\] net935
+ vssd1 vssd1 vccd1 vccd1 _04926_ sky130_fd_sc_hd__o221a_1
X_07935_ net1181 team_03_WB.instance_to_wrap.core.register_file.registers_state\[343\]
+ net766 team_03_WB.instance_to_wrap.core.register_file.registers_state\[375\] vssd1
+ vssd1 vccd1 vccd1 _03877_ sky130_fd_sc_hd__o22a_1
XANTENNA__09053__S0 net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_164_wb_clk_i clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_164_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout477_A net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13355__A net1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11427__X _06756_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07866_ net1167 _03807_ vssd1 vssd1 vccd1 vccd1 _03808_ sky130_fd_sc_hd__nor2_1
XANTENNA__10512__B1 net1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08181__A1 net1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09605_ _05459_ _05466_ net571 vssd1 vssd1 vccd1 vccd1 _05547_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_127_2984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08181__B2 net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07353__A net1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_1156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07797_ _03731_ _03732_ _03737_ _03738_ net1119 net1139 vssd1 vssd1 vccd1 vccd1 _03739_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_79_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout644_A net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout265_X net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1386_A net1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09536_ _05477_ vssd1 vssd1 vccd1 vccd1 _05478_ sky130_fd_sc_hd__inv_2
XANTENNA__09979__S net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10985__Y _06563_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09467_ net559 _05408_ vssd1 vssd1 vccd1 vccd1 _05409_ sky130_fd_sc_hd__nand2_1
XANTENNA__09681__A1 net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout811_A net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout909_A net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1174_X net1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08418_ net1229 team_03_WB.instance_to_wrap.core.register_file.registers_state\[218\]
+ net954 team_03_WB.instance_to_wrap.core.register_file.registers_state\[250\] net933
+ vssd1 vssd1 vccd1 vccd1 _04360_ sky130_fd_sc_hd__o221a_1
XANTENNA__12017__B1 net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_311 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09398_ _05170_ _05174_ _05338_ _05172_ _05167_ vssd1 vssd1 vccd1 vccd1 _05340_ sky130_fd_sc_hd__a311oi_4
XFILLER_0_46_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_1042 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08349_ net1063 _04288_ _04289_ vssd1 vssd1 vccd1 vccd1 _04291_ sky130_fd_sc_hd__or3_1
XANTENNA_fanout1341_X net1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10579__B1 net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_129_Right_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_128_Left_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_1075 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_539 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11240__A1 net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_794 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11360_ net490 net618 _06732_ net400 net2041 vssd1 vssd1 vccd1 vccd1 _02100_ sky130_fd_sc_hd__a32o_1
XFILLER_0_34_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08912__A net1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout899_X net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10311_ team_03_WB.instance_to_wrap.core.pc.current_pc\[30\] _06152_ vssd1 vssd1
+ vccd1 vccd1 _06153_ sky130_fd_sc_hd__nand2_1
XANTENNA__10653__S net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11291_ net712 net268 net829 vssd1 vssd1 vccd1 vccd1 _06713_ sky130_fd_sc_hd__and3_1
XFILLER_0_46_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08619__S0 net992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12434__A net1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13030_ net1300 vssd1 vssd1 vccd1 vccd1 _00794_ sky130_fd_sc_hd__inv_2
X_10242_ _06080_ _06081_ _06083_ vssd1 vssd1 vccd1 vccd1 _06084_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_104_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11543__A2 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08944__B1 net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10173_ _04954_ team_03_WB.instance_to_wrap.core.pc.current_pc\[10\] net675 vssd1
+ vssd1 vccd1 vccd1 _06015_ sky130_fd_sc_hd__mux2_1
Xfanout1103 net1104 vssd1 vssd1 vccd1 vccd1 net1103 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_28_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10751__B1 net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06955__C1 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1114 net1117 vssd1 vssd1 vccd1 vccd1 net1114 sky130_fd_sc_hd__buf_4
XFILLER_0_121_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1125 net1127 vssd1 vssd1 vccd1 vccd1 net1125 sky130_fd_sc_hd__buf_4
Xfanout1136 net1137 vssd1 vssd1 vccd1 vccd1 net1136 sky130_fd_sc_hd__buf_4
XFILLER_0_100_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input38_A gpio_in[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1147 net1148 vssd1 vssd1 vccd1 vccd1 net1147 sky130_fd_sc_hd__buf_6
X_14981_ clknet_leaf_65_wb_clk_i net34 _01346_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1158 net1159 vssd1 vssd1 vccd1 vccd1 net1158 sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_137_Left_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_156_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1169 team_03_WB.instance_to_wrap.core.decoder.inst\[21\] vssd1 vssd1 vccd1
+ vccd1 net1169 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_35_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13932_ clknet_leaf_16_wb_clk_i _01696_ _00297_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[286\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10503__B1 net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08172__A1 net1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13863_ clknet_leaf_114_wb_clk_i _01627_ _00228_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[217\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12814_ net1310 vssd1 vssd1 vccd1 vccd1 _00578_ sky130_fd_sc_hd__inv_2
X_13794_ clknet_leaf_172_wb_clk_i _01558_ _00159_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[148\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_83_2077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09632__A1_N team_03_WB.instance_to_wrap.core.decoder.inst\[28\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_486 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_2088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12745_ net1254 vssd1 vssd1 vccd1 vccd1 _00509_ sky130_fd_sc_hd__inv_2
XFILLER_0_57_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_151_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12008__B1 net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12676_ net1366 vssd1 vssd1 vccd1 vccd1 _00440_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_61_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_350 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_146_Left_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_13_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_133_3100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14415_ clknet_leaf_135_wb_clk_i _02179_ _00780_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[769\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_133_3111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11627_ _06701_ net382 net347 net2383 vssd1 vssd1 vccd1 vccd1 _01905_ sky130_fd_sc_hd__a22o_1
XFILLER_0_154_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10034__A2 net1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14346_ clknet_leaf_3_wb_clk_i _02110_ _00711_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[700\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07435__B1 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11558_ net2074 net485 _06793_ net513 vssd1 vssd1 vccd1 vccd1 _01963_ sky130_fd_sc_hd__a22o_1
XANTENNA__08632__C1 net1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08381__X _04323_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_684 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11659__S net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold608 team_03_WB.instance_to_wrap.core.register_file.registers_state\[854\] vssd1
+ vssd1 vccd1 vccd1 net2101 sky130_fd_sc_hd__dlygate4sd3_1
X_10509_ net159 net1030 net1025 net1729 vssd1 vssd1 vccd1 vccd1 _02601_ sky130_fd_sc_hd__a22o_1
XFILLER_0_40_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold619 team_03_WB.instance_to_wrap.core.register_file.registers_state\[874\] vssd1
+ vssd1 vccd1 vccd1 net2112 sky130_fd_sc_hd__dlygate4sd3_1
X_14277_ clknet_leaf_11_wb_clk_i _02041_ _00642_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[631\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_150_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11489_ _06609_ net2664 net388 vssd1 vssd1 vccd1 vccd1 _02017_ sky130_fd_sc_hd__mux2_1
XFILLER_0_40_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13228_ net1315 vssd1 vssd1 vccd1 vccd1 _00992_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_59_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08935__B1 net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13159_ net1395 vssd1 vssd1 vccd1 vccd1 _00923_ sky130_fd_sc_hd__inv_2
X_15052__1493 vssd1 vssd1 vccd1 vccd1 net1493 _15052__1493/LO sky130_fd_sc_hd__conb_1
XPHY_EDGE_ROW_155_Left_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07720_ net1197 team_03_WB.instance_to_wrap.core.register_file.registers_state\[589\]
+ net778 team_03_WB.instance_to_wrap.core.register_file.registers_state\[621\] net731
+ vssd1 vssd1 vccd1 vccd1 _03662_ sky130_fd_sc_hd__o221a_1
XANTENNA__11298__A1 net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08699__C1 net1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11837__A3 net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07173__A net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07651_ net746 _03590_ _03592_ net1119 vssd1 vssd1 vccd1 vccd1 _03593_ sky130_fd_sc_hd__o211ai_1
Xclkbuf_0_wb_clk_i wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_0_wb_clk_i sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_105_2523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07910__A1 net1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_116 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07582_ net1163 _03519_ _03521_ _03523_ net1138 vssd1 vssd1 vccd1 vccd1 _03524_ sky130_fd_sc_hd__a2111o_1
XANTENNA__11126__C _06414_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_157_3601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09321_ _05260_ _05261_ _05259_ vssd1 vssd1 vccd1 vccd1 _05263_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_122_2881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10738__S net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_153_3509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09252_ _03728_ _05147_ net608 vssd1 vssd1 vccd1 vccd1 _05194_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_8_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11470__A1 net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07674__B1 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_174_3970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08203_ _04141_ _04142_ _04143_ _04144_ net860 net935 vssd1 vssd1 vccd1 vccd1 _04145_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_173_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09183_ net572 _05124_ vssd1 vssd1 vccd1 vccd1 _05125_ sky130_fd_sc_hd__and2_1
XFILLER_0_90_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_170_3856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11710__X _06808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_170_3867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08134_ _03459_ _03489_ _03280_ _03314_ vssd1 vssd1 vccd1 vccd1 _04076_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_43_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_940 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10981__B net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08065_ net820 _04006_ vssd1 vssd1 vccd1 vccd1 _04007_ sky130_fd_sc_hd__nor2_1
XFILLER_0_102_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1134_A net1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09179__B1 net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07016_ net1099 team_03_WB.instance_to_wrap.core.register_file.registers_state\[835\]
+ net1155 vssd1 vssd1 vccd1 vccd1 _02958_ sky130_fd_sc_hd__a21o_1
XFILLER_0_144_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07729__A1 net1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout594_A net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11525__A2 net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08926__B1 net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1301_A net1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10733__B1 net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08967_ net1243 team_03_WB.instance_to_wrap.core.register_file.registers_state\[585\]
+ net986 team_03_WB.instance_to_wrap.core.register_file.registers_state\[617\] net928
+ vssd1 vssd1 vccd1 vccd1 _04909_ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout761_A net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout382_X net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout859_A net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07918_ net1187 team_03_WB.instance_to_wrap.core.register_file.registers_state\[815\]
+ net878 _02872_ vssd1 vssd1 vccd1 vccd1 _03860_ sky130_fd_sc_hd__a31o_1
X_08898_ net1239 team_03_WB.instance_to_wrap.core.register_file.registers_state\[76\]
+ net979 team_03_WB.instance_to_wrap.core.register_file.registers_state\[108\] net926
+ vssd1 vssd1 vccd1 vccd1 _04840_ sky130_fd_sc_hd__o221a_1
XFILLER_0_75_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07849_ net1189 team_03_WB.instance_to_wrap.core.register_file.registers_state\[699\]
+ net878 vssd1 vssd1 vccd1 vccd1 _03791_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout1291_X net1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout647_X net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07901__A1 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10860_ net1042 net1251 net1252 _02808_ vssd1 vssd1 vccd1 vccd1 _06459_ sky130_fd_sc_hd__or4_2
XFILLER_0_39_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09103__B1 net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07370__X _03312_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09519_ net565 _05460_ vssd1 vssd1 vccd1 vccd1 _05461_ sky130_fd_sc_hd__nand2_1
XFILLER_0_94_721 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10648__S net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09654__A1 net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10791_ _02829_ net688 _06399_ vssd1 vssd1 vccd1 vccd1 _06401_ sky130_fd_sc_hd__o21ai_4
XANTENNA_fanout814_X net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12530_ net1394 vssd1 vssd1 vccd1 vccd1 _00294_ sky130_fd_sc_hd__inv_2
XANTENNA__11333__A net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1148 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_404 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_61_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_61_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_137_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_990 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12461_ net1332 vssd1 vssd1 vccd1 vccd1 _00225_ sky130_fd_sc_hd__inv_2
X_14200_ clknet_leaf_4_wb_clk_i _01964_ _00565_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[554\]
+ sky130_fd_sc_hd__dfrtp_1
X_11412_ net273 net2462 net396 vssd1 vssd1 vccd1 vccd1 _02068_ sky130_fd_sc_hd__mux2_1
XANTENNA__09738__A net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08614__C1 net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12392_ net1293 vssd1 vssd1 vccd1 vccd1 _00156_ sky130_fd_sc_hd__inv_2
XFILLER_0_50_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07968__A1 net1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07512__S0 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11764__A2 net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14131_ clknet_leaf_105_wb_clk_i _01895_ _00496_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[485\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11343_ net1247 net836 net278 net668 vssd1 vssd1 vccd1 vccd1 _06724_ sky130_fd_sc_hd__and4_1
XFILLER_0_120_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09709__A2 _05041_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14062_ clknet_leaf_124_wb_clk_i _01826_ _00427_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[416\]
+ sky130_fd_sc_hd__dfrtp_1
X_11274_ net507 net635 _06704_ net410 net2148 vssd1 vssd1 vccd1 vccd1 _02158_ sky130_fd_sc_hd__a32o_1
XFILLER_0_123_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_37_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13013_ net1291 vssd1 vssd1 vccd1 vccd1 _00777_ sky130_fd_sc_hd__inv_2
X_10225_ _06008_ _06066_ vssd1 vssd1 vccd1 vccd1 _06067_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_37_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09185__A3 _05126_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08393__A1 net1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10156_ net590 net674 _05997_ vssd1 vssd1 vccd1 vccd1 _05998_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07264__Y _03206_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold5 team_03_WB.instance_to_wrap.core.register_file.registers_state\[929\] vssd1
+ vssd1 vccd1 vccd1 net1498 sky130_fd_sc_hd__dlygate4sd3_1
X_10087_ _05686_ _05697_ _05706_ _05930_ vssd1 vssd1 vccd1 vccd1 _05931_ sky130_fd_sc_hd__and4bb_1
X_14964_ clknet_leaf_101_wb_clk_i _02716_ _01329_ vssd1 vssd1 vccd1 vccd1 net216 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_85_2117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_169_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13915_ clknet_leaf_159_wb_clk_i _01679_ _00280_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[269\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_50_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14895_ clknet_leaf_64_wb_clk_i _02658_ _01260_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.pc.current_pc\[24\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA_clkload3_A clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09920__B _05596_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13846_ clknet_leaf_179_wb_clk_i _01610_ _00211_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[200\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_18_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09412__S net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07721__A net1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13777_ clknet_leaf_141_wb_clk_i _01541_ _00142_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[131\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07105__C1 net1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10989_ net280 net651 net704 net828 vssd1 vssd1 vccd1 vccd1 _06566_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_100_2420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08536__B _04476_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_2431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11243__A net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09860__D_N _05697_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07656__B1 net1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12728_ net1380 vssd1 vssd1 vccd1 vccd1 _00492_ sky130_fd_sc_hd__inv_2
XANTENNA__08853__C1 net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_704 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12659_ net1261 vssd1 vssd1 vccd1 vccd1 _00423_ sky130_fd_sc_hd__inv_2
XFILLER_0_115_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_167_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09648__A net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07959__A1 net1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold405 team_03_WB.instance_to_wrap.core.register_file.registers_state\[291\] vssd1
+ vssd1 vccd1 vccd1 net1898 sky130_fd_sc_hd__dlygate4sd3_1
X_14329_ clknet_leaf_168_wb_clk_i _02093_ _00694_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[683\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold416 team_03_WB.instance_to_wrap.core.register_file.registers_state\[252\] vssd1
+ vssd1 vccd1 vccd1 net1909 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold427 team_03_WB.instance_to_wrap.core.register_file.registers_state\[45\] vssd1
+ vssd1 vccd1 vccd1 net1920 sky130_fd_sc_hd__dlygate4sd3_1
Xhold438 team_03_WB.instance_to_wrap.core.register_file.registers_state\[816\] vssd1
+ vssd1 vccd1 vccd1 net1931 sky130_fd_sc_hd__dlygate4sd3_1
Xhold449 team_03_WB.instance_to_wrap.core.register_file.registers_state\[415\] vssd1
+ vssd1 vccd1 vccd1 net1942 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08908__B1 net1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout907 _06285_ vssd1 vssd1 vccd1 vccd1 net907 sky130_fd_sc_hd__clkbuf_4
X_09870_ _05811_ vssd1 vssd1 vccd1 vccd1 _05812_ sky130_fd_sc_hd__inv_2
XANTENNA__09176__A3 _05041_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout918 net923 vssd1 vssd1 vccd1 vccd1 net918 sky130_fd_sc_hd__buf_4
XANTENNA__09030__C1 net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12802__A net1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_1887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout929 net932 vssd1 vssd1 vccd1 vccd1 net929 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_74_1898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14997__Q team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[16\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08821_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[513\] net1006
+ _04762_ net1076 vssd1 vssd1 vccd1 vccd1 _04763_ sky130_fd_sc_hd__o211a_1
XFILLER_0_29_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_146_3368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1105 team_03_WB.instance_to_wrap.core.register_file.registers_state\[142\] vssd1
+ vssd1 vccd1 vccd1 net2598 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_146_3379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1116 team_03_WB.instance_to_wrap.core.register_file.registers_state\[586\] vssd1
+ vssd1 vccd1 vccd1 net2609 sky130_fd_sc_hd__dlygate4sd3_1
X_08752_ net1239 team_03_WB.instance_to_wrap.core.register_file.registers_state\[675\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[643\] net980 vssd1
+ vssd1 vccd1 vccd1 _04694_ sky130_fd_sc_hd__a22o_1
Xhold1127 team_03_WB.instance_to_wrap.core.register_file.registers_state\[201\] vssd1
+ vssd1 vccd1 vccd1 net2620 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1138 team_03_WB.instance_to_wrap.core.register_file.registers_state\[196\] vssd1
+ vssd1 vccd1 vccd1 net2631 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1149 team_03_WB.instance_to_wrap.core.register_file.registers_state\[720\] vssd1
+ vssd1 vccd1 vccd1 net2642 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_174_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07703_ net1197 team_03_WB.instance_to_wrap.core.register_file.registers_state\[173\]
+ net899 net1133 vssd1 vssd1 vccd1 vccd1 _03645_ sky130_fd_sc_hd__a211o_1
XFILLER_0_135_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_124_2921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08683_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[616\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[584\]
+ net975 vssd1 vssd1 vccd1 vccd1 _04625_ sky130_fd_sc_hd__mux2_1
XANTENNA__07344__C1 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11852__S net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07634_ net746 _03574_ net815 vssd1 vssd1 vccd1 vccd1 _03576_ sky130_fd_sc_hd__o21a_1
XANTENNA__10494__A2 net1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07631__A net1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07565_ net1200 team_03_WB.instance_to_wrap.core.register_file.registers_state\[600\]
+ net781 team_03_WB.instance_to_wrap.core.register_file.registers_state\[632\] net734
+ vssd1 vssd1 vccd1 vccd1 _03507_ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout342_A _06805_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09304_ _05244_ _05245_ vssd1 vssd1 vccd1 vccd1 _05246_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout1084_A net1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_172_3907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_480 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09100__A3 _05041_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07496_ net1109 team_03_WB.instance_to_wrap.core.register_file.registers_state\[711\]
+ net803 team_03_WB.instance_to_wrap.core.register_file.registers_state\[743\] net735
+ vssd1 vssd1 vccd1 vccd1 _03438_ sky130_fd_sc_hd__a221o_1
XFILLER_0_48_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09235_ _04235_ _05175_ vssd1 vssd1 vccd1 vccd1 _05177_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10992__A net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout607_A net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1349_A net1358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_11_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09166_ net436 net428 _04893_ net546 vssd1 vssd1 vccd1 vccd1 _05108_ sky130_fd_sc_hd__o31a_1
XFILLER_0_161_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08117_ net1087 team_03_WB.instance_to_wrap.core.register_file.registers_state\[890\]
+ net892 _04058_ net1124 vssd1 vssd1 vccd1 vccd1 _04059_ sky130_fd_sc_hd__o311a_1
XANTENNA__11746__A2 net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09097_ _05035_ _05036_ _05038_ _05037_ net941 net863 vssd1 vssd1 vccd1 vccd1 _05039_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__08611__A2 net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_1__f_wb_clk_i_A clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1137_X net1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09992__S net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_792 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08048_ _03945_ _03946_ _03986_ _03987_ vssd1 vssd1 vccd1 vccd1 _03990_ sky130_fd_sc_hd__o22a_1
Xhold950 team_03_WB.instance_to_wrap.core.register_file.registers_state\[176\] vssd1
+ vssd1 vccd1 vccd1 net2443 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10216__B _03206_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout976_A net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout597_X net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold961 team_03_WB.instance_to_wrap.core.register_file.registers_state\[496\] vssd1
+ vssd1 vccd1 vccd1 net2454 sky130_fd_sc_hd__dlygate4sd3_1
Xhold972 team_03_WB.instance_to_wrap.core.register_file.registers_state\[847\] vssd1
+ vssd1 vccd1 vccd1 net2465 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09167__A3 _04953_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold983 team_03_WB.instance_to_wrap.core.register_file.registers_state\[340\] vssd1
+ vssd1 vccd1 vccd1 net2476 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09021__C1 net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold994 team_03_WB.instance_to_wrap.core.register_file.registers_state\[795\] vssd1
+ vssd1 vccd1 vccd1 net2487 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10010_ net593 net1653 net287 vssd1 vssd1 vccd1 vccd1 _02704_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout764_X net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09999_ _05884_ net1701 net287 vssd1 vssd1 vccd1 vccd1 _02715_ sky130_fd_sc_hd__mux2_1
XANTENNA__07583__C1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08127__A1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11961_ net635 _06738_ net468 net365 net2669 vssd1 vssd1 vccd1 vccd1 _01582_ sky130_fd_sc_hd__a32o_1
XFILLER_0_153_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout931_X net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13543__A net1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10912_ net314 net309 _05928_ team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[11\]
+ vssd1 vssd1 vccd1 vccd1 _06502_ sky130_fd_sc_hd__or4b_1
X_13700_ clknet_leaf_30_wb_clk_i _01464_ _00065_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[54\]
+ sky130_fd_sc_hd__dfrtp_1
X_14680_ clknet_leaf_82_wb_clk_i _02444_ _01045_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.ADR_I\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_11892_ net630 _06701_ net462 net372 net2162 vssd1 vssd1 vccd1 vccd1 _01649_ sky130_fd_sc_hd__a32o_1
XFILLER_0_168_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_80_2014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13631_ net1421 vssd1 vssd1 vccd1 vccd1 _01395_ sky130_fd_sc_hd__inv_2
X_10843_ team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[21\] net305 vssd1
+ vssd1 vccd1 vccd1 _06443_ sky130_fd_sc_hd__and2_1
XANTENNA_clkbuf_leaf_50_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_2025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_434 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11063__A net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13562_ net1427 vssd1 vssd1 vccd1 vccd1 _01326_ sky130_fd_sc_hd__inv_2
XFILLER_0_165_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_491 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10774_ _02831_ _02838_ vssd1 vssd1 vccd1 vccd1 _06384_ sky130_fd_sc_hd__nand2_1
XFILLER_0_82_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15051__1492 vssd1 vssd1 vccd1 vccd1 net1492 _15051__1492/LO sky130_fd_sc_hd__conb_1
X_12513_ net1262 vssd1 vssd1 vccd1 vccd1 _00277_ sky130_fd_sc_hd__inv_2
XFILLER_0_136_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13493_ net1327 vssd1 vssd1 vccd1 vccd1 _01257_ sky130_fd_sc_hd__inv_2
XFILLER_0_82_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_256 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12444_ net1421 vssd1 vssd1 vccd1 vccd1 _00208_ sky130_fd_sc_hd__inv_2
XFILLER_0_48_1019 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12375_ net1385 vssd1 vssd1 vccd1 vccd1 _00139_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14114_ clknet_leaf_175_wb_clk_i _01878_ _00479_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[468\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09755__X _05697_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11326_ _06630_ net2726 net407 vssd1 vssd1 vccd1 vccd1 _02119_ sky130_fd_sc_hd__mux2_1
X_15094_ net1480 vssd1 vssd1 vccd1 vccd1 la_data_out[30] sky130_fd_sc_hd__buf_2
XFILLER_0_120_542 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07623__A_N _03278_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11937__S net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14045_ clknet_leaf_165_wb_clk_i _01809_ _00410_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[399\]
+ sky130_fd_sc_hd__dfrtp_1
X_11257_ net274 net709 net827 vssd1 vssd1 vccd1 vccd1 _06696_ sky130_fd_sc_hd__and3_1
XANTENNA__09915__B _05676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_3010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12622__A net1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08366__A1 net1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10208_ _06047_ _06048_ _06046_ vssd1 vssd1 vccd1 vccd1 _06050_ sky130_fd_sc_hd__a21o_1
XFILLER_0_98_1120 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11188_ net1043 net838 _06536_ net669 vssd1 vssd1 vccd1 vccd1 _06675_ sky130_fd_sc_hd__and4_2
XANTENNA__11370__B1 net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10139_ _03390_ _05980_ vssd1 vssd1 vccd1 vccd1 _05981_ sky130_fd_sc_hd__or2_1
XFILLER_0_89_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09931__A _03312_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14947_ clknet_leaf_55_wb_clk_i _00009_ _01312_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.wb.curr_state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_141_3265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11672__S net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_141_3276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11673__A1 net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14878_ clknet_leaf_88_wb_clk_i _02641_ _01243_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.pc.current_pc\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09142__S net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07341__A2 net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07451__A net1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09618__A1 net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13829_ clknet_leaf_14_wb_clk_i _01593_ _00194_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[183\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_159_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07629__B1 net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07350_ net1170 team_03_WB.instance_to_wrap.core.register_file.registers_state\[476\]
+ net757 team_03_WB.instance_to_wrap.core.register_file.registers_state\[508\] net1149
+ vssd1 vssd1 vccd1 vccd1 _03292_ sky130_fd_sc_hd__o221a_1
XFILLER_0_70_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11425__B2 net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08826__C1 net1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_426 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07281_ net751 _03220_ _03221_ net808 vssd1 vssd1 vccd1 vccd1 _03223_ sky130_fd_sc_hd__o211a_1
XFILLER_0_31_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09020_ net1244 team_03_WB.instance_to_wrap.core.register_file.registers_state\[80\]
+ net984 team_03_WB.instance_to_wrap.core.register_file.registers_state\[112\] net928
+ vssd1 vssd1 vccd1 vccd1 _04962_ sky130_fd_sc_hd__o221a_1
XFILLER_0_14_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11189__B1 net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_144 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11420__B _06751_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08054__B1 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold202 net227 vssd1 vssd1 vccd1 vccd1 net1695 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_117_2780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_1938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold213 net182 vssd1 vssd1 vccd1 vccd1 net1706 sky130_fd_sc_hd__dlygate4sd3_1
Xhold224 _02595_ vssd1 vssd1 vccd1 vccd1 net1717 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_339 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold235 net216 vssd1 vssd1 vccd1 vccd1 net1728 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07801__B1 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold246 net134 vssd1 vssd1 vccd1 vccd1 net1739 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_148_3408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_740 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_148_3419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07329__C net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold257 net194 vssd1 vssd1 vccd1 vccd1 net1750 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold268 team_03_WB.instance_to_wrap.ADR_I\[2\] vssd1 vssd1 vccd1 vccd1 net1761 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_113_2688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11847__S net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09922_ _05517_ _05541_ _05563_ vssd1 vssd1 vccd1 vccd1 _05864_ sky130_fd_sc_hd__or3_1
Xhold279 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1\] vssd1
+ vssd1 vccd1 vccd1 net1772 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_113_2699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09003__C1 net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout704 net708 vssd1 vssd1 vccd1 vccd1 net704 sky130_fd_sc_hd__clkbuf_8
Xfanout715 net716 vssd1 vssd1 vccd1 vccd1 net715 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08357__A1 net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout726 net727 vssd1 vssd1 vccd1 vccd1 net726 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_165_3755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09853_ net565 _05738_ vssd1 vssd1 vccd1 vccd1 _05795_ sky130_fd_sc_hd__nand2_1
XANTENNA__07626__A net1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout737 net738 vssd1 vssd1 vccd1 vccd1 net737 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_165_3766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08221__S net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout748 net749 vssd1 vssd1 vccd1 vccd1 net748 sky130_fd_sc_hd__buf_4
XANTENNA_fanout292_A net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout759 net760 vssd1 vssd1 vccd1 vccd1 net759 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07565__C1 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11148__A net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08804_ net1053 team_03_WB.instance_to_wrap.core.register_file.registers_state\[193\]
+ net1006 team_03_WB.instance_to_wrap.core.register_file.registers_state\[225\] net927
+ vssd1 vssd1 vccd1 vccd1 _04746_ sky130_fd_sc_hd__a221o_1
X_09784_ _03459_ _04619_ _05725_ _02945_ vssd1 vssd1 vccd1 vccd1 _05726_ sky130_fd_sc_hd__o22a_1
X_06996_ _02925_ _02927_ _02932_ _02934_ _02926_ vssd1 vssd1 vccd1 vccd1 _02938_ sky130_fd_sc_hd__o2111ai_4
XANTENNA__08109__A1 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08735_ _04674_ _04676_ net1208 vssd1 vssd1 vccd1 vccd1 _04677_ sky130_fd_sc_hd__o21a_1
XANTENNA__10987__A net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11582__S net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13363__A net1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout557_A net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1299_A net1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07868__B1 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11664__A1 _06505_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08666_ net1058 team_03_WB.instance_to_wrap.core.register_file.registers_state\[839\]
+ net1011 team_03_WB.instance_to_wrap.core.register_file.registers_state\[871\] team_03_WB.instance_to_wrap.core.decoder.inst\[17\]
+ vssd1 vssd1 vccd1 vccd1 _04608_ sky130_fd_sc_hd__a221o_1
XFILLER_0_163_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07617_ net1112 team_03_WB.instance_to_wrap.core.register_file.registers_state\[665\]
+ net735 _03547_ vssd1 vssd1 vccd1 vccd1 _03559_ sky130_fd_sc_hd__a211o_1
X_08597_ net1058 team_03_WB.instance_to_wrap.core.register_file.registers_state\[581\]
+ net1011 team_03_WB.instance_to_wrap.core.register_file.registers_state\[613\] net947
+ vssd1 vssd1 vccd1 vccd1 _04539_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout724_A _02863_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout345_X net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1087_X net1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09987__S net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07548_ _03489_ vssd1 vssd1 vccd1 vccd1 _03490_ sky130_fd_sc_hd__inv_2
XANTENNA__08817__C1 net1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_962 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_165_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07096__A1 net1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_134_wb_clk_i_A clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_63_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10926__S net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07479_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[789\] net793
+ _03420_ vssd1 vssd1 vccd1 vccd1 _03421_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout512_X net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_146_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09218_ _03823_ _05143_ _05159_ vssd1 vssd1 vccd1 vccd1 _05160_ sky130_fd_sc_hd__and3_1
XFILLER_0_134_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09288__A _04646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10490_ net110 net1029 net906 net1743 vssd1 vssd1 vccd1 vccd1 _02619_ sky130_fd_sc_hd__a22o_1
XFILLER_0_17_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_144 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_101_Left_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09149_ net543 _04296_ _05090_ vssd1 vssd1 vccd1 vccd1 _05091_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_16_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_20_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_952 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10927__B1 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12160_ net1523 vssd1 vssd1 vccd1 vccd1 _02393_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__08920__A net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout881_X net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09749__B1_N net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11111_ _06630_ net2679 net419 vssd1 vssd1 vccd1 vccd1 _02247_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout979_X net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10661__S net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12091_ net632 _06659_ net465 net441 net1756 vssd1 vssd1 vccd1 vccd1 _01456_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_9_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold780 team_03_WB.instance_to_wrap.core.register_file.registers_state\[777\] vssd1
+ vssd1 vccd1 vccd1 net2273 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold791 team_03_WB.instance_to_wrap.core.register_file.registers_state\[260\] vssd1
+ vssd1 vccd1 vccd1 net2284 sky130_fd_sc_hd__dlygate4sd3_1
X_11042_ net2198 net423 _06597_ net512 vssd1 vssd1 vccd1 vccd1 _02283_ sky130_fd_sc_hd__a22o_1
XANTENNA__11352__B1 net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07556__C1 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_110_Left_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14801_ clknet_leaf_85_wb_clk_i _02565_ _01166_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_I\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input20_A DAT_I[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09848__A1 net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07308__C1 net1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12993_ net1263 vssd1 vssd1 vccd1 vccd1 _00757_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11492__S net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1108 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14732_ clknet_leaf_61_wb_clk_i _02496_ _01097_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.decoder.inst\[29\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__11655__A1 _06454_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11944_ net627 _06721_ net458 net364 net2126 vssd1 vssd1 vccd1 vccd1 _01599_ sky130_fd_sc_hd__a32o_1
XANTENNA_clkbuf_leaf_173_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_99_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14663_ clknet_leaf_97_wb_clk_i _02427_ _01028_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1017\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_52_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11875_ net1043 net654 net701 net466 vssd1 vssd1 vccd1 vccd1 _06813_ sky130_fd_sc_hd__or4b_4
XFILLER_0_28_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10826_ _06427_ _06429_ net586 vssd1 vssd1 vccd1 vccd1 _06430_ sky130_fd_sc_hd__o21a_2
X_13614_ net1421 vssd1 vssd1 vccd1 vccd1 _01378_ sky130_fd_sc_hd__inv_2
XFILLER_0_139_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08808__C1 net1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14594_ clknet_leaf_176_wb_clk_i _02358_ _00959_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[948\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_28_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10757_ team_03_WB.instance_to_wrap.core.pc.current_pc\[4\] _05769_ net605 vssd1
+ vssd1 vccd1 vccd1 _06372_ sky130_fd_sc_hd__mux2_1
X_13545_ net1306 vssd1 vssd1 vccd1 vccd1 _01309_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_45_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_483 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_164_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13476_ net1430 vssd1 vssd1 vccd1 vccd1 _01240_ sky130_fd_sc_hd__inv_2
XFILLER_0_125_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10688_ net522 _06327_ _06328_ net527 net1848 vssd1 vssd1 vccd1 vccd1 _02464_ sky130_fd_sc_hd__a32o_1
XFILLER_0_54_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_2363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07210__S net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_987 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_2374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12427_ net1281 vssd1 vssd1 vccd1 vccd1 _00191_ sky130_fd_sc_hd__inv_2
XFILLER_0_51_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08036__B1 net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10137__A _03528_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_1114 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12358_ net1293 vssd1 vssd1 vccd1 vccd1 _00122_ sky130_fd_sc_hd__inv_2
XANTENNA__11591__A0 net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11667__S net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10933__A3 _06519_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11309_ _06619_ net2623 net405 vssd1 vssd1 vccd1 vccd1 _02136_ sky130_fd_sc_hd__mux2_1
X_15077_ net1463 vssd1 vssd1 vccd1 vccd1 la_data_out[13] sky130_fd_sc_hd__buf_2
XFILLER_0_121_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12289_ net1272 vssd1 vssd1 vccd1 vccd1 _00053_ sky130_fd_sc_hd__inv_2
XFILLER_0_10_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_71_1835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14028_ clknet_leaf_22_wb_clk_i _01792_ _00393_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[382\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_4_0__f_wb_clk_i_X clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_143_3305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_3316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06850_ net1249 vssd1 vssd1 vccd1 vccd1 _02793_ sky130_fd_sc_hd__inv_2
XANTENNA__08976__S net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11894__A1 net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10303__C _06144_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_160_3652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_160_3663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09839__A1 net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08520_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[63\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[31\]
+ net959 vssd1 vssd1 vccd1 vccd1 _04462_ sky130_fd_sc_hd__mux2_1
XANTENNA__13183__A net1347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07314__A2 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08511__A1 net1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08451_ _04391_ _04392_ net867 vssd1 vssd1 vccd1 vccd1 _04393_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_69_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07402_ net1171 team_03_WB.instance_to_wrap.core.register_file.registers_state\[991\]
+ vssd1 vssd1 vccd1 vccd1 _03344_ sky130_fd_sc_hd__or2_1
XFILLER_0_86_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_147_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08382_ _04323_ vssd1 vssd1 vccd1 vccd1 _04324_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_940 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11134__C net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_189_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_189_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_133_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07078__A1 net1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07333_ net1162 _03273_ _03274_ _03270_ vssd1 vssd1 vccd1 vccd1 _03275_ sky130_fd_sc_hd__o22a_1
XFILLER_0_129_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_162_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_119_2820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10973__C net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_118_wb_clk_i clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_118_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_144_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07264_ team_03_WB.instance_to_wrap.core.decoder.inst\[28\] net826 vssd1 vssd1 vccd1
+ vccd1 _03206_ sky130_fd_sc_hd__nand2_1
XANTENNA__09539__C _05125_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09003_ net1046 team_03_WB.instance_to_wrap.core.register_file.registers_state\[586\]
+ net995 team_03_WB.instance_to_wrap.core.register_file.registers_state\[618\] net933
+ vssd1 vssd1 vccd1 vccd1 _04945_ sky130_fd_sc_hd__a221o_1
XFILLER_0_170_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_115_2728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11150__B _06468_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_2739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07195_ _03108_ _03136_ net613 vssd1 vssd1 vccd1 vccd1 _03137_ sky130_fd_sc_hd__mux2_2
XFILLER_0_14_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10909__A0 net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout305_A net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08578__A1 net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1047_A net1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_167_3806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10385__A1 _06213_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11582__A0 _06430_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11577__S net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1214_A net1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout501 net502 vssd1 vssd1 vccd1 vccd1 net501 sky130_fd_sc_hd__clkbuf_4
X_09905_ net315 _05623_ _05632_ _05812_ vssd1 vssd1 vccd1 vccd1 _05847_ sky130_fd_sc_hd__nand4_1
Xfanout512 net513 vssd1 vssd1 vccd1 vccd1 net512 sky130_fd_sc_hd__buf_4
XFILLER_0_6_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout523 _06322_ vssd1 vssd1 vccd1 vccd1 net523 sky130_fd_sc_hd__buf_2
Xfanout534 _06298_ vssd1 vssd1 vccd1 vccd1 net534 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout674_A _05948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout545 _03106_ vssd1 vssd1 vccd1 vccd1 net545 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__11334__B1 net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout556 net557 vssd1 vssd1 vccd1 vccd1 net556 sky130_fd_sc_hd__buf_2
X_15050__1491 vssd1 vssd1 vccd1 vccd1 net1491 _15050__1491/LO sky130_fd_sc_hd__conb_1
X_09836_ net557 _04713_ _05777_ net566 vssd1 vssd1 vccd1 vccd1 _05778_ sky130_fd_sc_hd__a211o_1
Xfanout567 _03025_ vssd1 vssd1 vccd1 vccd1 net567 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11885__A1 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout578 _02993_ vssd1 vssd1 vccd1 vccd1 net578 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout1002_X net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08750__A1 net1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07553__A2 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout841_A _06304_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09767_ _05707_ _05708_ vssd1 vssd1 vccd1 vccd1 _05709_ sky130_fd_sc_hd__nor2_1
X_06979_ net724 _02906_ _02913_ _02920_ vssd1 vssd1 vccd1 vccd1 _02921_ sky130_fd_sc_hd__o22a_2
XANTENNA_fanout462_X net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08189__S0 net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout939_A net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08718_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[420\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[388\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[292\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[260\]
+ net985 net1079 vssd1 vssd1 vccd1 vccd1 _04660_ sky130_fd_sc_hd__mux4_1
X_09698_ _02804_ _03864_ _04820_ _05639_ vssd1 vssd1 vccd1 vccd1 _05640_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__07091__A net1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_139_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08649_ _04579_ _04590_ net852 vssd1 vssd1 vccd1 vccd1 _04591_ sky130_fd_sc_hd__mux2_4
XANTENNA_fanout727_X net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07710__C1 net1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11660_ net2054 _06623_ net343 vssd1 vssd1 vccd1 vccd1 _01873_ sky130_fd_sc_hd__mux2_1
X_10611_ net1809 team_03_WB.instance_to_wrap.CPU_DAT_O\[18\] net841 vssd1 vssd1 vccd1
+ vccd1 _02517_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_25_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_206 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10656__S net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11591_ net272 net2504 net450 vssd1 vssd1 vccd1 vccd1 _01938_ sky130_fd_sc_hd__mux2_1
XFILLER_0_147_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13330_ net1319 vssd1 vssd1 vccd1 vccd1 _01094_ sky130_fd_sc_hd__inv_2
XANTENNA__11341__A net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10542_ net1 _06284_ vssd1 vssd1 vccd1 vccd1 _06287_ sky130_fd_sc_hd__nand2_1
XFILLER_0_18_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1147 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13261_ net1292 vssd1 vssd1 vccd1 vccd1 _01025_ sky130_fd_sc_hd__inv_2
X_10473_ team_03_WB.instance_to_wrap.wb.curr_state\[2\] team_03_WB.instance_to_wrap.wb.curr_state\[1\]
+ vssd1 vssd1 vccd1 vccd1 _06284_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_40_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15000_ clknet_leaf_44_wb_clk_i net48 _01365_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_12212_ net1508 vssd1 vssd1 vccd1 vccd1 _02341_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__09766__B1 net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13192_ net1298 vssd1 vssd1 vccd1 vccd1 _00956_ sky130_fd_sc_hd__inv_2
XANTENNA__08650__A _04591_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input68_A wbs_adr_i[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_92_2260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12143_ net1585 vssd1 vssd1 vccd1 vccd1 _02410_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_92_2271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10244__X _06086_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_4_4__f_wb_clk_i clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_4__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
X_12074_ _06780_ net454 net439 net2045 vssd1 vssd1 vccd1 vccd1 _01473_ sky130_fd_sc_hd__a22o_1
XANTENNA__11325__A0 net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11025_ net651 _06586_ vssd1 vssd1 vccd1 vccd1 _06587_ sky130_fd_sc_hd__and2_1
XANTENNA__11876__A1 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08649__X _04591_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08741__A1 net1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input23_X net23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1099 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09912__C net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_99_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12976_ net1410 vssd1 vssd1 vccd1 vccd1 _00740_ sky130_fd_sc_hd__inv_2
X_14715_ clknet_leaf_48_wb_clk_i _02479_ _01080_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.decoder.inst\[12\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__11235__B net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11927_ _06625_ net2498 net369 vssd1 vssd1 vccd1 vccd1 _01615_ sky130_fd_sc_hd__mux2_1
XANTENNA__07432__C net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_157_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14646_ clknet_leaf_151_wb_clk_i _02410_ _01011_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1000\]
+ sky130_fd_sc_hd__dfstp_1
X_11858_ _06483_ net2376 net377 vssd1 vssd1 vccd1 vccd1 _01682_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_99_2403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_99_2414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_64_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10809_ team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[28\] net307 net685 vssd1
+ vssd1 vccd1 vccd1 _06416_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_28_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11789_ net2381 _06469_ net327 vssd1 vssd1 vccd1 vccd1 _01749_ sky130_fd_sc_hd__mux2_1
X_14577_ clknet_leaf_140_wb_clk_i _02341_ _00942_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[931\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__11251__A net1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_136_3164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_3175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13528_ net1316 vssd1 vssd1 vccd1 vccd1 _01292_ sky130_fd_sc_hd__inv_2
XANTENNA__11800__A1 _06519_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09927__Y _05868_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13459_ net1327 vssd1 vssd1 vccd1 vccd1 _01223_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_140_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09757__B1 net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput104 net104 vssd1 vssd1 vccd1 vccd1 ADR_O[10] sky130_fd_sc_hd__clkbuf_4
Xoutput115 net115 vssd1 vssd1 vccd1 vccd1 ADR_O[20] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_2_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput126 net126 vssd1 vssd1 vccd1 vccd1 ADR_O[30] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_100_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput137 net137 vssd1 vssd1 vccd1 vccd1 DAT_O[10] sky130_fd_sc_hd__clkbuf_4
XANTENNA__10906__A3 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13178__A net1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput148 net148 vssd1 vssd1 vccd1 vccd1 DAT_O[20] sky130_fd_sc_hd__buf_2
XFILLER_0_121_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_110_2625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10017__D net72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput159 net159 vssd1 vssd1 vccd1 vccd1 DAT_O[30] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_142_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_110_2636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12108__A2 net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08980__A1 net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07951_ net1128 _03888_ _03889_ _03891_ net1141 vssd1 vssd1 vccd1 vccd1 _03893_ sky130_fd_sc_hd__a311o_1
XANTENNA__11316__A0 _06623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_162_3703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06902_ net1017 net1015 net1018 vssd1 vssd1 vccd1 vccd1 _02844_ sky130_fd_sc_hd__o21a_1
XFILLER_0_128_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07882_ net1090 team_03_WB.instance_to_wrap.core.register_file.registers_state\[47\]
+ net894 vssd1 vssd1 vccd1 vccd1 _03824_ sky130_fd_sc_hd__or3_1
XFILLER_0_128_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11129__C net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08193__C1 net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08732__A1 net1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06833_ team_03_WB.instance_to_wrap.WRITE_I vssd1 vssd1 vccd1 vccd1 _02776_ sky130_fd_sc_hd__inv_2
X_09621_ net581 _05543_ _05544_ _05562_ vssd1 vssd1 vccd1 vccd1 _05563_ sky130_fd_sc_hd__a31oi_4
X_09552_ _05391_ _05395_ net562 vssd1 vssd1 vccd1 vccd1 _05494_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_108_2587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08503_ _04444_ vssd1 vssd1 vccd1 vccd1 _04445_ sky130_fd_sc_hd__inv_2
X_09483_ _03641_ _04503_ net535 _05424_ _03639_ vssd1 vssd1 vccd1 vccd1 _05425_ sky130_fd_sc_hd__o311a_1
XANTENNA__08496__B1 net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11860__S net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08434_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[826\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[794\]
+ net964 vssd1 vssd1 vccd1 vccd1 _04376_ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06954__S net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10984__B net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_22_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_392 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08365_ net1063 _04304_ _04305_ vssd1 vssd1 vccd1 vccd1 _04307_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_22_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout422_A _06560_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1164_A net1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07316_ _03256_ _03257_ net812 vssd1 vssd1 vccd1 vccd1 _03258_ sky130_fd_sc_hd__a21o_1
XFILLER_0_163_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_72 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08296_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[56\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[24\]
+ net987 vssd1 vssd1 vccd1 vccd1 _04238_ sky130_fd_sc_hd__mux2_1
XFILLER_0_144_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07247_ net1191 team_03_WB.instance_to_wrap.core.register_file.registers_state\[40\]
+ net881 vssd1 vssd1 vccd1 vccd1 _03189_ sky130_fd_sc_hd__and3_1
XFILLER_0_5_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_171_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1012 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1331_A net1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07178_ net1115 _03117_ _03118_ vssd1 vssd1 vccd1 vccd1 _03120_ sky130_fd_sc_hd__or3_1
XANTENNA__10358__A1 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09212__A2 _03428_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout791_A net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08470__A net1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout889_A net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13088__A net1402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_86_wb_clk_i clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_86_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__11100__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1217_X net1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07774__A2 net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1307 net1309 vssd1 vssd1 vccd1 vccd1 net1307 sky130_fd_sc_hd__buf_4
Xfanout320 _05355_ vssd1 vssd1 vccd1 vccd1 net320 sky130_fd_sc_hd__clkbuf_4
Xfanout1318 net1320 vssd1 vssd1 vccd1 vccd1 net1318 sky130_fd_sc_hd__buf_4
XFILLER_0_79_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_15_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_15_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xfanout1329 net1330 vssd1 vssd1 vccd1 vccd1 net1329 sky130_fd_sc_hd__buf_4
Xfanout331 _06809_ vssd1 vssd1 vccd1 vccd1 net331 sky130_fd_sc_hd__buf_6
Xfanout342 _06805_ vssd1 vssd1 vccd1 vccd1 net342 sky130_fd_sc_hd__buf_8
Xfanout353 _04776_ vssd1 vssd1 vccd1 vccd1 net353 sky130_fd_sc_hd__clkbuf_2
Xfanout364 _06815_ vssd1 vssd1 vccd1 vccd1 net364 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12720__A net1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout375 _06812_ vssd1 vssd1 vccd1 vccd1 net375 sky130_fd_sc_hd__clkbuf_8
XANTENNA__08184__C1 net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout386 net387 vssd1 vssd1 vccd1 vccd1 net386 sky130_fd_sc_hd__buf_2
X_09819_ net583 _04679_ net537 _05760_ vssd1 vssd1 vccd1 vccd1 _05761_ sky130_fd_sc_hd__o31ai_1
Xfanout397 _06752_ vssd1 vssd1 vccd1 vccd1 net397 sky130_fd_sc_hd__buf_4
XANTENNA_fanout844_X net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12830_ net1414 vssd1 vssd1 vccd1 vccd1 _00594_ sky130_fd_sc_hd__inv_2
XANTENNA__10240__A _03944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_112 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11055__B net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12761_ net1359 vssd1 vssd1 vccd1 vccd1 _00525_ sky130_fd_sc_hd__inv_2
XFILLER_0_68_167 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14500_ clknet_leaf_22_wb_clk_i _02264_ _00865_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[854\]
+ sky130_fd_sc_hd__dfrtp_1
X_11712_ net2106 _06409_ net335 vssd1 vssd1 vccd1 vccd1 _01824_ sky130_fd_sc_hd__mux2_1
X_12692_ net1312 vssd1 vssd1 vccd1 vccd1 _00456_ sky130_fd_sc_hd__inv_2
XFILLER_0_90_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_154_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11643_ net1248 _06462_ net382 vssd1 vssd1 vccd1 vccd1 _06805_ sky130_fd_sc_hd__and3_4
X_14431_ clknet_leaf_166_wb_clk_i _02195_ _00796_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[785\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_65_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12035__A1 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_42_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09987__A0 _05872_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11574_ _06447_ _06394_ vssd1 vssd1 vccd1 vccd1 _06800_ sky130_fd_sc_hd__and2b_1
X_14362_ clknet_leaf_144_wb_clk_i _02126_ _00727_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[716\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_94_2300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput17 DAT_I[23] vssd1 vssd1 vccd1 vccd1 net17 sky130_fd_sc_hd__buf_1
Xinput28 DAT_I[4] vssd1 vssd1 vccd1 vccd1 net28 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08083__C net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10525_ net141 net1032 net1024 net1773 vssd1 vssd1 vccd1 vccd1 _02585_ sky130_fd_sc_hd__a22o_1
X_13313_ net1308 vssd1 vssd1 vccd1 vccd1 _01077_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_2311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput39 gpio_in[14] vssd1 vssd1 vccd1 vccd1 net39 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_134_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14293_ clknet_leaf_107_wb_clk_i _02057_ _00658_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[647\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_161_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13244_ net1422 vssd1 vssd1 vccd1 vccd1 _01008_ sky130_fd_sc_hd__inv_2
X_10456_ _06051_ _06052_ vssd1 vssd1 vccd1 vccd1 _06271_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_131_3061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_3072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11546__B1 net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_2219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13175_ net1385 vssd1 vssd1 vccd1 vccd1 _00939_ sky130_fd_sc_hd__inv_2
XANTENNA__11010__A2 net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10387_ team_03_WB.instance_to_wrap.core.pc.current_pc\[17\] _06143_ vssd1 vssd1
+ vccd1 vccd1 _06215_ sky130_fd_sc_hd__nor2_1
X_12126_ net1583 vssd1 vssd1 vccd1 vccd1 _02427_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__08962__A1 net1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06973__B1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12057_ _06623_ net2331 net356 vssd1 vssd1 vccd1 vccd1 _01489_ sky130_fd_sc_hd__mux2_1
XFILLER_0_165_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08714__A1 net1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07724__A net1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11008_ net711 net701 net300 vssd1 vssd1 vccd1 vccd1 _06577_ sky130_fd_sc_hd__or3b_1
XFILLER_0_133_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_66_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_1138 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12959_ net1347 vssd1 vssd1 vccd1 vccd1 _00723_ sky130_fd_sc_hd__inv_2
XFILLER_0_90_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_3204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08573__S0 net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10824__A2 net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_3215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07150__B1 net1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_2484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_103_2495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14629_ clknet_leaf_40_wb_clk_i _02393_ _00994_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[983\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_172_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_155_3551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_155_3562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09978__A0 _03023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08150_ net1230 team_03_WB.instance_to_wrap.core.register_file.registers_state\[84\]
+ net960 team_03_WB.instance_to_wrap.core.register_file.registers_state\[116\] net919
+ vssd1 vssd1 vccd1 vccd1 _04092_ sky130_fd_sc_hd__o221a_1
XFILLER_0_16_727 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_34 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07101_ team_03_WB.instance_to_wrap.core.decoder.inst\[23\] _03042_ _03036_ net718
+ vssd1 vssd1 vccd1 vccd1 _03043_ sky130_fd_sc_hd__a211o_2
XANTENNA__10588__B2 _03103_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07453__A1 net1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08081_ net1088 team_03_WB.instance_to_wrap.core.register_file.registers_state\[950\]
+ net894 vssd1 vssd1 vccd1 vccd1 _04023_ sky130_fd_sc_hd__or3_1
XFILLER_0_141_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09386__A _04267_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07032_ net1196 team_03_WB.instance_to_wrap.core.register_file.registers_state\[131\]
+ vssd1 vssd1 vccd1 vccd1 _02974_ sky130_fd_sc_hd__or2_1
XFILLER_0_140_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_218 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_140_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_3_0_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_0_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__07205__A1 net1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08402__B1 net1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08983_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[10\] net996
+ net918 _04924_ vssd1 vssd1 vccd1 vccd1 _04925_ sky130_fd_sc_hd__o211a_1
XANTENNA__11855__S net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07934_ net812 _03871_ _03872_ _03875_ vssd1 vssd1 vccd1 vccd1 _03876_ sky130_fd_sc_hd__o22a_1
XANTENNA__08166__C1 net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09053__S1 net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07865_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[443\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[411\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[315\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[283\]
+ net783 net1136 vssd1 vssd1 vccd1 vccd1 _03807_ sky130_fd_sc_hd__mux4_1
XANTENNA__07064__S0 net1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout372_A _06813_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_2974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09604_ _05545_ vssd1 vssd1 vccd1 vccd1 _05546_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_127_2985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07796_ _03733_ _03734_ net749 vssd1 vssd1 vccd1 vccd1 _03738_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09535_ _05371_ _05463_ _05468_ _05472_ _05476_ vssd1 vssd1 vccd1 vccd1 _05477_ sky130_fd_sc_hd__a221o_2
XTAP_TAPCELL_ROW_27_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09666__C1 _05607_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1281_A net1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_133_wb_clk_i clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_133_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout637_A net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11590__S net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1379_A net1380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09466_ net547 _04417_ _05094_ vssd1 vssd1 vccd1 vccd1 _05408_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_93_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_149_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08465__A net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_148_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_164_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08417_ net1228 team_03_WB.instance_to_wrap.core.register_file.registers_state\[90\]
+ net954 team_03_WB.instance_to_wrap.core.register_file.registers_state\[122\] net917
+ vssd1 vssd1 vccd1 vccd1 _04359_ sky130_fd_sc_hd__o221a_1
X_09397_ _05170_ _05174_ _05338_ _05172_ vssd1 vssd1 vccd1 vccd1 _05339_ sky130_fd_sc_hd__a31o_1
XFILLER_0_148_397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout804_A net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1167_X net1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09995__S net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08348_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[437\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[405\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[309\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[277\]
+ net972 net1074 vssd1 vssd1 vccd1 vccd1 _04290_ sky130_fd_sc_hd__mux4_1
XFILLER_0_11_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_163_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08279_ net1220 _04220_ vssd1 vssd1 vccd1 vccd1 _04221_ sky130_fd_sc_hd__or2_1
XANTENNA__11240__A2 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10310_ team_03_WB.instance_to_wrap.core.pc.current_pc\[29\] team_03_WB.instance_to_wrap.core.pc.current_pc\[28\]
+ _06151_ vssd1 vssd1 vccd1 vccd1 _06152_ sky130_fd_sc_hd__and3_1
XANTENNA__09296__A _03459_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11290_ net511 net639 _06712_ net411 net2145 vssd1 vssd1 vccd1 vccd1 _02150_ sky130_fd_sc_hd__a32o_1
XFILLER_0_21_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11528__B1 net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout794_X net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08619__S1 net1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10241_ _06082_ vssd1 vssd1 vccd1 vccd1 _06083_ sky130_fd_sc_hd__inv_2
XFILLER_0_104_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08944__A1 net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10172_ _06013_ vssd1 vssd1 vccd1 vccd1 _06014_ sky130_fd_sc_hd__inv_2
XFILLER_0_100_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07247__C net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout961_X net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10751__A1 net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06955__B1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1104 net1105 vssd1 vssd1 vccd1 vccd1 net1104 sky130_fd_sc_hd__clkbuf_4
Xfanout1115 net1117 vssd1 vssd1 vccd1 vccd1 net1115 sky130_fd_sc_hd__clkbuf_4
Xfanout1126 net1127 vssd1 vssd1 vccd1 vccd1 net1126 sky130_fd_sc_hd__buf_2
X_14980_ clknet_leaf_91_wb_clk_i _02732_ _01345_ vssd1 vssd1 vccd1 vccd1 net232 sky130_fd_sc_hd__dfrtp_1
Xfanout1137 _02785_ vssd1 vssd1 vccd1 vccd1 net1137 sky130_fd_sc_hd__buf_6
Xfanout1148 team_03_WB.instance_to_wrap.core.decoder.inst\[23\] vssd1 vssd1 vccd1
+ vccd1 net1148 sky130_fd_sc_hd__buf_12
XFILLER_0_22_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_156_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1159 team_03_WB.instance_to_wrap.core.decoder.inst\[22\] vssd1 vssd1 vccd1
+ vccd1 net1159 sky130_fd_sc_hd__buf_6
XANTENNA__08157__C1 net1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13931_ clknet_leaf_38_wb_clk_i _01695_ _00296_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[285\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10503__A1 net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11700__B1 net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07904__C1 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11066__A net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_87_2170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13862_ clknet_leaf_73_wb_clk_i _01626_ _00227_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[216\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_159_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12813_ net1311 vssd1 vssd1 vccd1 vccd1 _00577_ sky130_fd_sc_hd__inv_2
XFILLER_0_69_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13793_ clknet_leaf_181_wb_clk_i _01557_ _00158_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[147\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08555__S0 net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_2078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_2089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12744_ net1297 vssd1 vssd1 vccd1 vccd1 _00508_ sky130_fd_sc_hd__inv_2
XFILLER_0_69_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12675_ net1356 vssd1 vssd1 vccd1 vccd1 _00439_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_61_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14414_ clknet_leaf_125_wb_clk_i _02178_ _00779_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[768\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_133_3101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11626_ _06700_ net385 net348 net2454 vssd1 vssd1 vccd1 vccd1 _01906_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_133_3112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11767__B1 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_710 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14345_ clknet_leaf_70_wb_clk_i _02109_ _00710_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[699\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09918__B _02837_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11557_ net658 _06667_ vssd1 vssd1 vccd1 vccd1 _06793_ sky130_fd_sc_hd__nor2_1
XFILLER_0_8_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08632__B1 net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10508_ net160 net1031 net1023 net1758 vssd1 vssd1 vccd1 vccd1 _02602_ sky130_fd_sc_hd__a22o_1
XFILLER_0_12_218 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold609 team_03_WB.instance_to_wrap.core.register_file.registers_state\[48\] vssd1
+ vssd1 vccd1 vccd1 net2102 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11488_ net1248 _06449_ net650 _06463_ vssd1 vssd1 vccd1 vccd1 _06778_ sky130_fd_sc_hd__or4_4
X_14276_ clknet_leaf_24_wb_clk_i _02040_ _00641_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[630\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_100_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10990__B2 net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10439_ net285 _06137_ _06257_ net682 vssd1 vssd1 vccd1 vccd1 _06258_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_111_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13227_ net1287 vssd1 vssd1 vccd1 vccd1 _00991_ sky130_fd_sc_hd__inv_2
XANTENNA__10145__A _03109_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13158_ net1301 vssd1 vssd1 vccd1 vccd1 _00922_ sky130_fd_sc_hd__inv_2
XANTENNA__10742__A1 _05686_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11675__S net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12109_ net1142 team_03_WB.instance_to_wrap.core.ru.state\[0\] team_03_WB.instance_to_wrap.core.ru.state\[5\]
+ _06281_ net840 vssd1 vssd1 vccd1 vccd1 _06821_ sky130_fd_sc_hd__a221o_1
X_13089_ net1262 vssd1 vssd1 vccd1 vccd1 _00853_ sky130_fd_sc_hd__inv_2
XANTENNA__12360__A net1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08148__C1 net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08699__B1 net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11298__A2 net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_98 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09360__A1 _05278_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08163__A2 net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07650_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[654\] net777
+ net730 _03591_ vssd1 vssd1 vccd1 vccd1 _03592_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_105_2524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07371__B1 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_2535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07581_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[792\] net794
+ net1041 _03522_ vssd1 vssd1 vccd1 vccd1 _03523_ sky130_fd_sc_hd__o211a_1
XFILLER_0_125_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11126__D net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_240 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_157_3602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09320_ _05259_ _05261_ vssd1 vssd1 vccd1 vccd1 _05262_ sky130_fd_sc_hd__nand2b_1
XANTENNA__09112__A1 net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_122_2871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_122_2882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09251_ _05183_ _05187_ _05192_ vssd1 vssd1 vccd1 vccd1 _05193_ sky130_fd_sc_hd__or3_1
XANTENNA__07674__A1 net1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_735 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11470__A2 net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_174_3960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08202_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[1011\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[979\]
+ net957 vssd1 vssd1 vccd1 vccd1 _04144_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_174_3971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09182_ _03061_ _03062_ _03066_ _03104_ vssd1 vssd1 vccd1 vccd1 _05124_ sky130_fd_sc_hd__and4b_1
XFILLER_0_90_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11758__B1 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_170_3857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08133_ _03137_ _03170_ _04073_ _04074_ vssd1 vssd1 vccd1 vccd1 _04075_ sky130_fd_sc_hd__nand4_1
XFILLER_0_161_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_170_3868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_952 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_540 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08064_ net1163 _04004_ _04005_ vssd1 vssd1 vccd1 vccd1 _04006_ sky130_fd_sc_hd__o21a_1
XFILLER_0_70_173 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09179__A1 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07015_ net1196 team_03_WB.instance_to_wrap.core.register_file.registers_state\[867\]
+ net883 vssd1 vssd1 vccd1 vccd1 _02957_ sky130_fd_sc_hd__and3_1
XANTENNA__09179__B2 net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08387__C1 net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1127_A _02785_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08926__A1 net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09844__A net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10194__C1 _02893_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07067__C net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11585__S net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08966_ _04902_ _04907_ net874 vssd1 vssd1 vccd1 vccd1 _04908_ sky130_fd_sc_hd__mux2_1
X_07917_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[911\] net781
+ _03858_ vssd1 vssd1 vccd1 vccd1 _03859_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout754_A net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08897_ net1239 team_03_WB.instance_to_wrap.core.register_file.registers_state\[204\]
+ net979 team_03_WB.instance_to_wrap.core.register_file.registers_state\[236\] net942
+ vssd1 vssd1 vccd1 vccd1 _04839_ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout375_X net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10497__B1 net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07848_ _03788_ _03789_ net611 vssd1 vssd1 vccd1 vccd1 _03790_ sky130_fd_sc_hd__mux2_2
XFILLER_0_168_404 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_162_Right_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_40_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout921_A net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07779_ net815 _03719_ _03720_ net818 vssd1 vssd1 vccd1 vccd1 _03721_ sky130_fd_sc_hd__o211ai_1
XANTENNA__09103__A1 net1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09518_ _05379_ _05382_ net561 vssd1 vssd1 vccd1 vccd1 _05460_ sky130_fd_sc_hd__mux2_1
XFILLER_0_116_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10790_ _02829_ net688 _06399_ vssd1 vssd1 vccd1 vccd1 _06400_ sky130_fd_sc_hd__o21a_1
XANTENNA__11997__A0 net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07114__B1 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08311__C1 net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11333__B net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07665__A1 net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09449_ net546 net350 _05108_ vssd1 vssd1 vccd1 vccd1 _05391_ sky130_fd_sc_hd__o21ba_1
XANTENNA__07530__C net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout807_X net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_164_654 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12460_ net1314 vssd1 vssd1 vccd1 vccd1 _00224_ sky130_fd_sc_hd__inv_2
XANTENNA__11749__B1 net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11411_ _06468_ net2643 net396 vssd1 vssd1 vccd1 vccd1 _02069_ sky130_fd_sc_hd__mux2_1
XANTENNA__08614__B1 net1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12391_ net1368 vssd1 vssd1 vccd1 vccd1 _00155_ sky130_fd_sc_hd__inv_2
XFILLER_0_34_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11342_ net502 net629 _06723_ net401 net1907 vssd1 vssd1 vccd1 vccd1 _02109_ sky130_fd_sc_hd__a32o_1
XFILLER_0_105_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14130_ clknet_leaf_165_wb_clk_i _01894_ _00495_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[484\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07512__S1 net1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_387 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_30_wb_clk_i clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_30_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_104_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11273_ net712 net297 net829 vssd1 vssd1 vccd1 vccd1 _06704_ sky130_fd_sc_hd__and3_1
X_14061_ clknet_leaf_186_wb_clk_i _01825_ _00426_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[415\]
+ sky130_fd_sc_hd__dfrtp_1
X_10224_ _06012_ _06065_ vssd1 vssd1 vccd1 vccd1 _06066_ sky130_fd_sc_hd__nand2_1
XANTENNA_input50_A gpio_in[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13012_ net1304 vssd1 vssd1 vccd1 vccd1 _00776_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_37_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11495__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10155_ team_03_WB.instance_to_wrap.core.pc.current_pc\[16\] net674 vssd1 vssd1 vccd1
+ vccd1 _05997_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_89_2210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_54_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10086_ _05718_ _05730_ net319 _05929_ vssd1 vssd1 vccd1 vccd1 _05930_ sky130_fd_sc_hd__and4b_1
Xhold6 team_03_WB.instance_to_wrap.core.register_file.registers_state\[953\] vssd1
+ vssd1 vccd1 vccd1 net1499 sky130_fd_sc_hd__dlygate4sd3_1
X_14963_ clknet_leaf_103_wb_clk_i _02715_ _01328_ vssd1 vssd1 vccd1 vccd1 net215 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_85_2118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10488__B1 net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13914_ clknet_leaf_146_wb_clk_i _01678_ _00279_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[268\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_85_2129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14894_ clknet_leaf_63_wb_clk_i _02657_ _01259_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.pc.current_pc\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_50_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09893__A2 _04323_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13845_ clknet_leaf_129_wb_clk_i _01609_ _00210_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[199\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_162_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11524__A net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13776_ clknet_leaf_160_wb_clk_i _01540_ _00141_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[130\]
+ sky130_fd_sc_hd__dfrtp_1
X_10988_ net2361 net420 _06565_ net490 vssd1 vssd1 vccd1 vccd1 _02305_ sky130_fd_sc_hd__a22o_1
XFILLER_0_128_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_100_2421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_2432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11243__B net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07656__A1 net1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12727_ net1392 vssd1 vssd1 vccd1 vccd1 _00491_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08853__B1 net1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09929__A _03277_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12658_ net1396 vssd1 vssd1 vccd1 vccd1 _00422_ sky130_fd_sc_hd__inv_2
XFILLER_0_154_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_378 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11609_ net650 net461 vssd1 vssd1 vccd1 vccd1 _06803_ sky130_fd_sc_hd__nand2_2
XFILLER_0_4_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12589_ net1331 vssd1 vssd1 vccd1 vccd1 _00353_ sky130_fd_sc_hd__inv_2
XFILLER_0_68_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_170_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07959__A2 net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11755__A3 net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14328_ clknet_leaf_19_wb_clk_i _02092_ _00693_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[682\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_871 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold406 team_03_WB.instance_to_wrap.core.register_file.registers_state\[267\] vssd1
+ vssd1 vccd1 vccd1 net1899 sky130_fd_sc_hd__dlygate4sd3_1
Xhold417 team_03_WB.instance_to_wrap.core.register_file.registers_state\[396\] vssd1
+ vssd1 vccd1 vccd1 net1910 sky130_fd_sc_hd__dlygate4sd3_1
Xhold428 team_03_WB.instance_to_wrap.core.register_file.registers_state\[406\] vssd1
+ vssd1 vccd1 vccd1 net1921 sky130_fd_sc_hd__dlygate4sd3_1
Xhold439 team_03_WB.instance_to_wrap.core.register_file.registers_state\[61\] vssd1
+ vssd1 vccd1 vccd1 net1932 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_78_1980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09935__Y _05872_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14259_ clknet_leaf_99_wb_clk_i _02023_ _00624_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[613\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_111_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08369__C1 net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07736__X _03678_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09030__B1 net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout908 _06285_ vssd1 vssd1 vccd1 vccd1 net908 sky130_fd_sc_hd__clkbuf_2
Xfanout919 net923 vssd1 vssd1 vccd1 vccd1 net919 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_29_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_74_1888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07041__C1 net1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08820_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[545\] net983
+ vssd1 vssd1 vccd1 vccd1 _04762_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_74_1899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_146_3369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07592__B1 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1106 team_03_WB.instance_to_wrap.core.register_file.registers_state\[94\] vssd1
+ vssd1 vccd1 vccd1 net2599 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1117 team_03_WB.instance_to_wrap.core.register_file.registers_state\[922\] vssd1
+ vssd1 vccd1 vccd1 net2610 sky130_fd_sc_hd__dlygate4sd3_1
X_08751_ _04687_ _04692_ net873 vssd1 vssd1 vccd1 vccd1 _04693_ sky130_fd_sc_hd__mux2_1
Xhold1128 team_03_WB.instance_to_wrap.core.register_file.registers_state\[664\] vssd1
+ vssd1 vccd1 vccd1 net2621 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07615__C net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1139 team_03_WB.instance_to_wrap.core.register_file.registers_state\[355\] vssd1
+ vssd1 vccd1 vccd1 net2632 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10479__B1 net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07702_ net1104 net899 team_03_WB.instance_to_wrap.core.register_file.registers_state\[141\]
+ vssd1 vssd1 vccd1 vccd1 _03644_ sky130_fd_sc_hd__o21a_1
XFILLER_0_75_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_124_2922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08682_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[552\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[520\]
+ net975 vssd1 vssd1 vccd1 vccd1 _04624_ sky130_fd_sc_hd__mux2_1
XFILLER_0_174_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07344__B1 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09603__S net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07633_ net1094 team_03_WB.instance_to_wrap.core.register_file.registers_state\[206\]
+ net798 team_03_WB.instance_to_wrap.core.register_file.registers_state\[238\] net730
+ vssd1 vssd1 vccd1 vccd1 _03575_ sky130_fd_sc_hd__a221o_1
XFILLER_0_71_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07895__A1 net1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11691__A2 net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07564_ _03504_ _03505_ net822 vssd1 vssd1 vccd1 vccd1 _03506_ sky130_fd_sc_hd__o21a_1
XANTENNA__11979__A0 net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09303_ _04591_ _05243_ vssd1 vssd1 vccd1 vccd1 _05245_ sky130_fd_sc_hd__nor2_1
XFILLER_0_76_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_172_3908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07647__A1 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_254 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07495_ net1110 team_03_WB.instance_to_wrap.core.register_file.registers_state\[583\]
+ net803 team_03_WB.instance_to_wrap.core.register_file.registers_state\[615\] net752
+ vssd1 vssd1 vccd1 vccd1 _03437_ sky130_fd_sc_hd__a221o_1
XFILLER_0_158_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_124_wb_clk_i_A clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout335_A net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10651__A0 team_03_WB.instance_to_wrap.core.decoder.inst\[10\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1077_A net1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09234_ _04235_ _05175_ vssd1 vssd1 vccd1 vccd1 _05176_ sky130_fd_sc_hd__nor2_1
XFILLER_0_119_879 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_3_Right_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_173_451 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_490 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09165_ net576 _05106_ _05093_ vssd1 vssd1 vccd1 vccd1 _05107_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_173_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout502_A net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12265__A net1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1244_A net1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08116_ net1181 team_03_WB.instance_to_wrap.core.register_file.registers_state\[858\]
+ vssd1 vssd1 vccd1 vccd1 _04058_ sky130_fd_sc_hd__or2_1
XFILLER_0_161_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_142_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09096_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[877\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[845\]
+ net989 vssd1 vssd1 vccd1 vccd1 _05038_ sky130_fd_sc_hd__mux2_1
XFILLER_0_142_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08047_ _03988_ vssd1 vssd1 vccd1 vccd1 _03989_ sky130_fd_sc_hd__inv_2
XFILLER_0_101_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_7_wb_clk_i_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout1032_X net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold940 team_03_WB.instance_to_wrap.core.register_file.registers_state\[416\] vssd1
+ vssd1 vccd1 vccd1 net2433 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold951 team_03_WB.instance_to_wrap.core.register_file.registers_state\[555\] vssd1
+ vssd1 vccd1 vccd1 net2444 sky130_fd_sc_hd__dlygate4sd3_1
Xhold962 team_03_WB.instance_to_wrap.core.register_file.registers_state\[278\] vssd1
+ vssd1 vccd1 vccd1 net2455 sky130_fd_sc_hd__dlygate4sd3_1
Xhold973 team_03_WB.instance_to_wrap.core.register_file.registers_state\[853\] vssd1
+ vssd1 vccd1 vccd1 net2466 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09021__B1 net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold984 team_03_WB.instance_to_wrap.core.register_file.registers_state\[533\] vssd1
+ vssd1 vccd1 vccd1 net2477 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout871_A net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout492_X net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold995 team_03_WB.instance_to_wrap.core.register_file.registers_state\[88\] vssd1
+ vssd1 vccd1 vccd1 net2488 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout969_A net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11903__B1 net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15115__1486 vssd1 vssd1 vccd1 vccd1 _15115__1486/HI net1486 sky130_fd_sc_hd__conb_1
XANTENNA__11609__A net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09998_ net587 net1728 net287 vssd1 vssd1 vccd1 vccd1 _02716_ sky130_fd_sc_hd__mux2_1
XANTENNA__08780__C1 net1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08949_ net873 _04889_ _04890_ vssd1 vssd1 vccd1 vccd1 _04891_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_4_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10800__X _06409_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11960_ net637 _06737_ net469 net365 net2025 vssd1 vssd1 vccd1 vccd1 _01583_ sky130_fd_sc_hd__a32o_1
XFILLER_0_98_324 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_163_wb_clk_i_A clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09875__A2 _04820_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_174_Left_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10911_ net312 _05845_ net318 _02780_ vssd1 vssd1 vccd1 vccd1 _06501_ sky130_fd_sc_hd__a31o_1
XANTENNA__10659__S net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07886__A1 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout924_X net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11682__A2 net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11891_ net642 _06700_ net473 net374 net2105 vssd1 vssd1 vccd1 vccd1 _01650_ sky130_fd_sc_hd__a32o_1
XFILLER_0_98_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_169_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13630_ net1421 vssd1 vssd1 vccd1 vccd1 _01394_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_80_2015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10890__B1 net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09088__B1 net1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_2026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10842_ net300 net2452 net519 vssd1 vssd1 vccd1 vccd1 _02328_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11063__B net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13561_ net1430 vssd1 vssd1 vccd1 vccd1 _01325_ sky130_fd_sc_hd__inv_2
X_10773_ _02802_ _02807_ _02822_ _02827_ vssd1 vssd1 vccd1 vccd1 _06383_ sky130_fd_sc_hd__or4_1
XFILLER_0_54_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10642__A0 team_03_WB.instance_to_wrap.core.decoder.inst\[19\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12512_ net1395 vssd1 vssd1 vccd1 vccd1 _00276_ sky130_fd_sc_hd__inv_2
X_13492_ net1327 vssd1 vssd1 vccd1 vccd1 _01256_ sky130_fd_sc_hd__inv_2
XANTENNA_input98_A wbs_adr_i[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12443_ net1362 vssd1 vssd1 vccd1 vccd1 _00207_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_268 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07269__A net1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08063__A1 net1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_860 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12374_ net1258 vssd1 vssd1 vccd1 vccd1 _00138_ sky130_fd_sc_hd__inv_2
XFILLER_0_62_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08091__C net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14113_ clknet_leaf_177_wb_clk_i _01877_ _00478_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[467\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07271__C1 net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11325_ net265 net2741 net406 vssd1 vssd1 vccd1 vccd1 _02120_ sky130_fd_sc_hd__mux2_1
X_15093_ net1479 vssd1 vssd1 vccd1 vccd1 la_data_out[29] sky130_fd_sc_hd__buf_2
XANTENNA__12903__A net1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_554 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14044_ clknet_leaf_157_wb_clk_i _01808_ _00409_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[398\]
+ sky130_fd_sc_hd__dfrtp_1
X_11256_ net499 net627 _06695_ net409 net2239 vssd1 vssd1 vccd1 vccd1 _02167_ sky130_fd_sc_hd__a32o_1
XFILLER_0_63_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06901__A net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_3000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_3011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10207_ _06046_ _06048_ vssd1 vssd1 vccd1 vccd1 _06049_ sky130_fd_sc_hd__nand2b_1
X_11187_ net516 net657 _06674_ net415 net1881 vssd1 vssd1 vccd1 vccd1 _02215_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_52_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1132 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11370__A1 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10138_ _04119_ _02772_ net673 vssd1 vssd1 vccd1 vccd1 _05980_ sky130_fd_sc_hd__mux2_1
XANTENNA__09931__B net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14946_ clknet_leaf_55_wb_clk_i _00008_ _01311_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.wb.curr_state\[1\]
+ sky130_fd_sc_hd__dfrtp_2
X_10069_ _02825_ _05910_ _05911_ _05912_ vssd1 vssd1 vccd1 vccd1 _05913_ sky130_fd_sc_hd__or4_1
XANTENNA__09866__A2 _05126_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08523__C1 net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_141_3266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_141_3277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07877__A1 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14877_ clknet_leaf_88_wb_clk_i _02640_ _01242_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.pc.current_pc\[6\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_159_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13828_ clknet_leaf_35_wb_clk_i _01592_ _00193_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[182\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_106_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08266__C _04207_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11425__A2 net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13759_ clknet_leaf_171_wb_clk_i _01523_ _00124_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[113\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10633__A0 team_03_WB.instance_to_wrap.core.decoder.inst\[28\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07280_ _03218_ _03219_ net813 vssd1 vssd1 vccd1 vccd1 _03222_ sky130_fd_sc_hd__o21a_1
XFILLER_0_45_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08563__A net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09011__X _04953_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_170_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11189__A1 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08054__A1 net1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_2770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold203 team_03_WB.instance_to_wrap.CPU_DAT_I\[20\] vssd1 vssd1 vccd1 vccd1 net1696
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_117_2781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_1928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_1939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold214 net188 vssd1 vssd1 vccd1 vccd1 net1707 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09665__Y _05607_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold225 team_03_WB.instance_to_wrap.CPU_DAT_I\[13\] vssd1 vssd1 vccd1 vccd1 net1718
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold236 team_03_WB.instance_to_wrap.CPU_DAT_I\[30\] vssd1 vssd1 vccd1 vccd1 net1729
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_148_3409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold247 net206 vssd1 vssd1 vccd1 vccd1 net1740 sky130_fd_sc_hd__dlygate4sd3_1
Xhold258 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[28\] vssd1 vssd1 vccd1
+ vccd1 net1751 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_752 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09394__A _04415_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09921_ _05435_ _05453_ _05500_ _05843_ _05862_ vssd1 vssd1 vccd1 vccd1 _05863_ sky130_fd_sc_hd__o2111ai_1
Xhold269 team_03_WB.instance_to_wrap.core.register_file.registers_state\[0\] vssd1
+ vssd1 vccd1 vccd1 net1762 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07907__A net1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_2689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09003__B1 net995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08502__S net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout705 net706 vssd1 vssd1 vccd1 vccd1 net705 sky130_fd_sc_hd__clkbuf_4
Xfanout716 _06460_ vssd1 vssd1 vccd1 vccd1 net716 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_165_3756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09852_ net578 _05683_ vssd1 vssd1 vccd1 vccd1 _05794_ sky130_fd_sc_hd__nor2_1
Xfanout727 net738 vssd1 vssd1 vccd1 vccd1 net727 sky130_fd_sc_hd__clkbuf_4
Xfanout738 _02853_ vssd1 vssd1 vccd1 vccd1 net738 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_165_3767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout749 net754 vssd1 vssd1 vccd1 vccd1 net749 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07565__B1 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09681__X _05623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08803_ net1053 team_03_WB.instance_to_wrap.core.register_file.registers_state\[65\]
+ net1006 team_03_WB.instance_to_wrap.core.register_file.registers_state\[97\] net942
+ vssd1 vssd1 vccd1 vccd1 _04745_ sky130_fd_sc_hd__a221o_1
XANTENNA__11148__B net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11900__A3 net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09783_ _03459_ _04619_ _04816_ vssd1 vssd1 vccd1 vccd1 _05725_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07345__C net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06995_ _02925_ _02927_ _02932_ _02934_ _02926_ vssd1 vssd1 vccd1 vccd1 _02937_ sky130_fd_sc_hd__o2111a_4
XANTENNA_fanout285_A net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08734_ net1222 _04672_ _04675_ net1075 vssd1 vssd1 vccd1 vccd1 _04676_ sky130_fd_sc_hd__o211a_1
XANTENNA__10987__B net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07868__A1 net1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08665_ _04601_ _04606_ net874 vssd1 vssd1 vccd1 vccd1 _04607_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout452_A net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1194_A net1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11164__A net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07616_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[537\] net787
+ net753 _03557_ vssd1 vssd1 vccd1 vccd1 _03558_ sky130_fd_sc_hd__a211o_1
XANTENNA__10872__B1 net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08596_ _02954_ _04537_ vssd1 vssd1 vccd1 vccd1 _04538_ sky130_fd_sc_hd__and2_1
XFILLER_0_49_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_70 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_165_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07547_ _03460_ _03488_ net615 vssd1 vssd1 vccd1 vccd1 _03489_ sky130_fd_sc_hd__mux2_4
XFILLER_0_36_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1361_A net1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout717_A net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout338_X net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_147_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07478_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[821\] net770
+ net1041 vssd1 vssd1 vccd1 vccd1 _03420_ sky130_fd_sc_hd__o21a_1
XANTENNA__11967__A3 net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09217_ _03567_ _03904_ _05155_ _02937_ vssd1 vssd1 vccd1 vccd1 _05159_ sky130_fd_sc_hd__o31ai_2
XFILLER_0_173_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout505_X net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1247_X net1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11103__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09856__X _05798_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07089__A net1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08045__A1 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09148_ net433 net427 _04119_ net548 vssd1 vssd1 vccd1 vccd1 _05090_ sky130_fd_sc_hd__o31a_1
XFILLER_0_133_156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10927__A1 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_370 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07253__C1 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09079_ net863 _05017_ _05020_ vssd1 vssd1 vccd1 vccd1 _05021_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_130_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11110_ net834 net269 vssd1 vssd1 vccd1 vccd1 _06630_ sky130_fd_sc_hd__and2_1
XFILLER_0_32_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_4_3__f_wb_clk_i clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_3__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
X_12090_ _06789_ net462 net440 net1859 vssd1 vssd1 vccd1 vccd1 _01457_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_9_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout874_X net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold770 team_03_WB.instance_to_wrap.core.register_file.registers_state\[891\] vssd1
+ vssd1 vccd1 vccd1 net2263 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold781 team_03_WB.instance_to_wrap.core.register_file.registers_state\[363\] vssd1
+ vssd1 vccd1 vccd1 net2274 sky130_fd_sc_hd__dlygate4sd3_1
Xhold792 team_03_WB.instance_to_wrap.core.register_file.registers_state\[376\] vssd1
+ vssd1 vccd1 vccd1 net2285 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11339__A net1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11041_ net640 _06596_ vssd1 vssd1 vccd1 vccd1 _06597_ sky130_fd_sc_hd__nor2_1
XANTENNA__11352__A1 net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07556__B1 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14800_ clknet_leaf_87_wb_clk_i _02564_ _01165_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_I\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08919__Y _04861_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07308__B1 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12992_ net1400 vssd1 vssd1 vccd1 vccd1 _00756_ sky130_fd_sc_hd__inv_2
XANTENNA__10897__B _05821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07552__A net1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14731_ clknet_leaf_54_wb_clk_i _02495_ _01096_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.decoder.inst\[28\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA_input13_A DAT_I[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11943_ net620 _06720_ net453 net363 net2159 vssd1 vssd1 vccd1 vccd1 _01600_ sky130_fd_sc_hd__a32o_1
XANTENNA__08000__X _03942_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11074__A net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14662_ clknet_leaf_71_wb_clk_i _02426_ _01027_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1016\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_54_1057 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11874_ net266 net2354 net378 vssd1 vssd1 vccd1 vccd1 _01666_ sky130_fd_sc_hd__mux2_1
XFILLER_0_157_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_204 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13613_ net1269 vssd1 vssd1 vccd1 vccd1 _01377_ sky130_fd_sc_hd__inv_2
X_10825_ team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[25\] net305 _06428_ net691
+ vssd1 vssd1 vccd1 vccd1 _06429_ sky130_fd_sc_hd__o211a_1
X_14593_ clknet_leaf_179_wb_clk_i _02357_ _00958_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[947\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_82_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10076__D1 _02937_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_900 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09479__A net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13544_ net1316 vssd1 vssd1 vccd1 vccd1 _01308_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11958__A3 net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10756_ net1863 net530 net525 _06371_ vssd1 vssd1 vccd1 vccd1 _02439_ sky130_fd_sc_hd__a22o_1
XANTENNA__09481__B1 net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12080__A2 net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_165_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_45_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11521__B net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13475_ net1430 vssd1 vssd1 vccd1 vccd1 _01239_ sky130_fd_sc_hd__inv_2
X_10687_ _06314_ _06325_ net606 vssd1 vssd1 vccd1 vccd1 _06328_ sky130_fd_sc_hd__a21o_1
XFILLER_0_125_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_97_2364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_97_2375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12426_ net1279 vssd1 vssd1 vccd1 vccd1 _00190_ sky130_fd_sc_hd__inv_2
XANTENNA__08036__A1 net1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_964 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09784__A1 _03459_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_1078 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09784__B2 _02945_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12357_ net1353 vssd1 vssd1 vccd1 vccd1 _00121_ sky130_fd_sc_hd__inv_2
XFILLER_0_51_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_1126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11308_ _06618_ net2561 net405 vssd1 vssd1 vccd1 vccd1 _02137_ sky130_fd_sc_hd__mux2_1
X_15076_ net1462 vssd1 vssd1 vccd1 vccd1 la_data_out[12] sky130_fd_sc_hd__buf_2
X_12288_ net1402 vssd1 vssd1 vccd1 vccd1 _00052_ sky130_fd_sc_hd__inv_2
XANTENNA__11249__A net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14027_ clknet_leaf_41_wb_clk_i _01791_ _00392_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[381\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10153__A _03985_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_1836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11239_ net1247 net837 _06413_ net670 vssd1 vssd1 vccd1 vccd1 _06687_ sky130_fd_sc_hd__and4_1
XANTENNA__07547__A0 _03460_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_143_3306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08744__C1 net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_143_3317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13464__A net1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_160_3653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_160_3664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14929_ clknet_leaf_43_wb_clk_i _02684_ _01294_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_O\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_69_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08450_ _04387_ _04388_ net859 vssd1 vssd1 vccd1 vccd1 _04392_ sky130_fd_sc_hd__o21a_1
XFILLER_0_33_1108 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07401_ net1171 team_03_WB.instance_to_wrap.core.register_file.registers_state\[863\]
+ vssd1 vssd1 vccd1 vccd1 _03343_ sky130_fd_sc_hd__or2_1
XFILLER_0_19_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08381_ net851 _04309_ _04322_ vssd1 vssd1 vccd1 vccd1 _04323_ sky130_fd_sc_hd__o21a_4
XANTENNA__11134__D net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07332_ net1152 _03271_ _03272_ net1116 vssd1 vssd1 vccd1 vccd1 _03274_ sky130_fd_sc_hd__a31o_1
XANTENNA__08275__A1 net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11949__A3 net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_900 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_2810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_2821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07263_ net723 _03188_ _03197_ _03204_ vssd1 vssd1 vccd1 vccd1 _03205_ sky130_fd_sc_hd__o2bb2a_4
XFILLER_0_61_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09002_ _04940_ _04943_ net1207 vssd1 vssd1 vccd1 vccd1 _04944_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_143_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_115_2729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11150__C net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07194_ _03122_ _03135_ net721 vssd1 vssd1 vccd1 vccd1 _03136_ sky130_fd_sc_hd__mux2_8
XFILLER_0_171_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11858__S net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09775__A1 net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_158_wb_clk_i clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_158_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_42_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_167_3807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07196__X _03138_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07250__A2 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09904_ _05844_ _05454_ _05429_ _05542_ vssd1 vssd1 vccd1 vccd1 _05846_ sky130_fd_sc_hd__or4bb_2
Xfanout502 net517 vssd1 vssd1 vccd1 vccd1 net502 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_6_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11159__A net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout513 net517 vssd1 vssd1 vccd1 vccd1 net513 sky130_fd_sc_hd__clkbuf_4
Xfanout524 _06322_ vssd1 vssd1 vccd1 vccd1 net524 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11334__A1 net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07538__B1 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout535 net536 vssd1 vssd1 vccd1 vccd1 net535 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout1207_A net1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout546 _03106_ vssd1 vssd1 vccd1 vccd1 net546 sky130_fd_sc_hd__buf_2
XANTENNA__09852__A net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09835_ _04566_ _04593_ net561 vssd1 vssd1 vccd1 vccd1 _05777_ sky130_fd_sc_hd__o21a_1
Xfanout557 net558 vssd1 vssd1 vccd1 vccd1 net557 sky130_fd_sc_hd__buf_2
XANTENNA_input5_A DAT_I[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout568 net569 vssd1 vssd1 vccd1 vccd1 net568 sky130_fd_sc_hd__clkbuf_4
Xfanout579 _02993_ vssd1 vssd1 vccd1 vccd1 net579 sky130_fd_sc_hd__buf_1
XANTENNA_fanout288_X net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout667_A _04818_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11593__S net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09766_ _05239_ _05271_ _05273_ net595 vssd1 vssd1 vccd1 vccd1 _05708_ sky130_fd_sc_hd__a31o_1
X_06978_ net814 _02916_ _02918_ _02919_ net819 vssd1 vssd1 vccd1 vccd1 _02920_ sky130_fd_sc_hd__o311a_1
XANTENNA__08189__S1 net1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08717_ net1048 team_03_WB.instance_to_wrap.core.register_file.registers_state\[452\]
+ net999 team_03_WB.instance_to_wrap.core.register_file.registers_state\[484\] net1079
+ vssd1 vssd1 vccd1 vccd1 _04659_ sky130_fd_sc_hd__a221o_1
XANTENNA__11637__A2 net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09697_ _03866_ net589 vssd1 vssd1 vccd1 vccd1 _05639_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout834_A _06387_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout455_X net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1197_X net1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10002__S net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08648_ _04582_ _04583_ _04589_ _04586_ net1066 net1081 vssd1 vssd1 vccd1 vccd1 _04590_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_96_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07710__B1 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08579_ _04519_ _04520_ net1220 vssd1 vssd1 vccd1 vccd1 _04521_ sky130_fd_sc_hd__o21a_1
XFILLER_0_3_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout622_X net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1364_X net1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09299__A _04619_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10610_ net1556 team_03_WB.instance_to_wrap.CPU_DAT_O\[19\] net841 vssd1 vssd1 vccd1
+ vccd1 _02518_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_1039 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08407__S net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11590_ _06477_ net2076 net447 vssd1 vssd1 vccd1 vccd1 _01939_ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_148_1018 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11341__B net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10541_ net1621 net1031 net1023 vssd1 vssd1 vccd1 vccd1 _02569_ sky130_fd_sc_hd__a21o_1
XFILLER_0_134_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11270__B1 net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_920 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08018__A1 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13260_ net1315 vssd1 vssd1 vccd1 vccd1 _01024_ sky130_fd_sc_hd__inv_2
X_10472_ team_03_WB.instance_to_wrap.wb.curr_state\[2\] team_03_WB.instance_to_wrap.wb.curr_state\[1\]
+ vssd1 vssd1 vccd1 vccd1 _06283_ sky130_fd_sc_hd__nor2_1
XFILLER_0_162_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09215__B1 _02937_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout991_X net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_161_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_40_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12211_ net1519 vssd1 vssd1 vccd1 vccd1 _02342_ sky130_fd_sc_hd__clkbuf_1
X_13191_ net1399 vssd1 vssd1 vccd1 vccd1 _00955_ sky130_fd_sc_hd__inv_2
XANTENNA__10376__A2 _06144_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11573__B2 net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_2261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12142_ net1516 vssd1 vssd1 vccd1 vccd1 _02411_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_92_2272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12073_ _05908_ _06394_ vssd1 vssd1 vccd1 vccd1 _06819_ sky130_fd_sc_hd__nand2b_4
XANTENNA__08726__C1 net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11024_ net1043 net838 net299 net671 vssd1 vssd1 vccd1 vccd1 _06586_ sky130_fd_sc_hd__and4_1
XANTENNA__07282__A net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_17 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input16_X net16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11628__A2 net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07713__C net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12975_ net1336 vssd1 vssd1 vccd1 vccd1 _00739_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14714_ clknet_leaf_31_wb_clk_i _02478_ _01079_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.decoder.inst\[11\]
+ sky130_fd_sc_hd__dfrtp_4
X_11926_ _06624_ net2601 net369 vssd1 vssd1 vccd1 vccd1 _01616_ sky130_fd_sc_hd__mux2_1
XANTENNA__11235__C net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_7 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14645_ clknet_leaf_106_wb_clk_i _02409_ _01010_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[999\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__10847__S net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11857_ _06681_ net456 net375 net2005 vssd1 vssd1 vccd1 vccd1 _01683_ sky130_fd_sc_hd__a22o_1
XFILLER_0_170_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_248 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12628__A net1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_99_2404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11532__A _06430_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_2415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10808_ team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[28\] net305 vssd1
+ vssd1 vccd1 vccd1 _06415_ sky130_fd_sc_hd__nand2_1
XANTENNA__08257__A1 net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14576_ clknet_leaf_159_wb_clk_i _02340_ _00941_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[930\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_64_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11788_ net2476 _06454_ net327 vssd1 vssd1 vccd1 vccd1 _01750_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_64_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13527_ net1329 vssd1 vssd1 vccd1 vccd1 _01291_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_136_3165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11251__B net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10739_ net1526 net529 net524 _06361_ vssd1 vssd1 vccd1 vccd1 _02446_ sky130_fd_sc_hd__a22o_1
XFILLER_0_82_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_3176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_780 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09937__A _03563_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13458_ net1323 vssd1 vssd1 vccd1 vccd1 _01222_ sky130_fd_sc_hd__inv_2
XANTENNA__07480__A2 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_402 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12409_ net1365 vssd1 vssd1 vccd1 vccd1 _00173_ sky130_fd_sc_hd__inv_2
XFILLER_0_140_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput105 net105 vssd1 vssd1 vccd1 vccd1 ADR_O[11] sky130_fd_sc_hd__clkbuf_4
X_13389_ net1421 vssd1 vssd1 vccd1 vccd1 _01153_ sky130_fd_sc_hd__inv_2
Xoutput116 net116 vssd1 vssd1 vccd1 vccd1 ADR_O[21] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_2_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput127 net127 vssd1 vssd1 vccd1 vccd1 ADR_O[31] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_50_271 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11564__B2 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07457__A net1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput138 net138 vssd1 vssd1 vccd1 vccd1 DAT_O[11] sky130_fd_sc_hd__buf_2
Xoutput149 net149 vssd1 vssd1 vccd1 vccd1 DAT_O[21] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_110_2626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_2637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15059_ net1445 vssd1 vssd1 vccd1 vccd1 gpio_out[36] sky130_fd_sc_hd__buf_2
XANTENNA__09943__Y _05876_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07950_ net1088 team_03_WB.instance_to_wrap.core.register_file.registers_state\[951\]
+ net893 vssd1 vssd1 vccd1 vccd1 _03892_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_162_3704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08717__C1 net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06901_ net1019 _02834_ _02838_ _02841_ vssd1 vssd1 vccd1 vccd1 _02843_ sky130_fd_sc_hd__or4_1
X_07881_ _03821_ _03822_ net610 vssd1 vssd1 vccd1 vccd1 _03823_ sky130_fd_sc_hd__mux2_1
XANTENNA__11129__D net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08193__B1 net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09620_ _05549_ _05561_ vssd1 vssd1 vccd1 vccd1 _05562_ sky130_fd_sc_hd__or2_2
X_06832_ team_03_WB.instance_to_wrap.core.pc.current_pc\[2\] vssd1 vssd1 vccd1 vccd1
+ _02775_ sky130_fd_sc_hd__inv_2
XANTENNA__07940__B1 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09551_ _05392_ _05416_ net555 vssd1 vssd1 vccd1 vccd1 _05493_ sky130_fd_sc_hd__mux2_1
XANTENNA__11619__A2 net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_2588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10827__A0 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08502_ _04430_ _04443_ net848 vssd1 vssd1 vccd1 vccd1 _04444_ sky130_fd_sc_hd__mux2_4
X_09482_ _03641_ _04503_ net664 _05423_ vssd1 vssd1 vccd1 vccd1 _05424_ sky130_fd_sc_hd__a22o_1
XANTENNA__08496__A1 net1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_13__f_wb_clk_i_A clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08433_ net1207 _04371_ _04374_ vssd1 vssd1 vccd1 vccd1 _04375_ sky130_fd_sc_hd__or3_1
XANTENNA__10757__S net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_516 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_842 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08364_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[438\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[406\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[310\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[278\]
+ net965 net1073 vssd1 vssd1 vccd1 vccd1 _04306_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_22_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10055__B2 team_03_WB.instance_to_wrap.CPU_DAT_O\[8\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_07315_ net1089 team_03_WB.instance_to_wrap.core.register_file.registers_state\[669\]
+ net728 _03245_ vssd1 vssd1 vccd1 vccd1 _03257_ sky130_fd_sc_hd__a211o_1
XANTENNA__11252__B1 net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08295_ net432 net424 _04236_ vssd1 vssd1 vccd1 vccd1 _04237_ sky130_fd_sc_hd__or3_1
XFILLER_0_144_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout415_A _06635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1157_A net1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07246_ _03180_ _03187_ net1164 vssd1 vssd1 vccd1 vccd1 _03188_ sky130_fd_sc_hd__mux2_1
XANTENNA__07471__A2 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11588__S net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1024 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07177_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[435\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[403\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[307\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[275\]
+ net763 net1125 vssd1 vssd1 vccd1 vccd1 _03119_ sky130_fd_sc_hd__mux4_1
XFILLER_0_131_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1324_A net1330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07759__B1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11555__B2 net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08420__A1 net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout784_A net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout310 _05845_ vssd1 vssd1 vccd1 vccd1 net310 sky130_fd_sc_hd__clkbuf_4
Xfanout1308 net1309 vssd1 vssd1 vccd1 vccd1 net1308 sky130_fd_sc_hd__buf_4
XANTENNA_fanout1112_X net1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1319 net1320 vssd1 vssd1 vccd1 vccd1 net1319 sky130_fd_sc_hd__clkbuf_4
Xfanout321 _04833_ vssd1 vssd1 vccd1 vccd1 net321 sky130_fd_sc_hd__clkbuf_4
Xfanout332 _06809_ vssd1 vssd1 vccd1 vccd1 net332 sky130_fd_sc_hd__buf_4
Xfanout343 _06805_ vssd1 vssd1 vccd1 vccd1 net343 sky130_fd_sc_hd__buf_4
XANTENNA_input8_X net8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout572_X net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout951_A net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08184__B1 net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout365 _06815_ vssd1 vssd1 vccd1 vccd1 net365 sky130_fd_sc_hd__clkbuf_8
Xfanout376 _06812_ vssd1 vssd1 vccd1 vccd1 net376 sky130_fd_sc_hd__buf_4
X_09818_ _02892_ _04679_ net667 _05759_ vssd1 vssd1 vccd1 vccd1 _05760_ sky130_fd_sc_hd__a22o_1
Xfanout387 _06802_ vssd1 vssd1 vccd1 vccd1 net387 sky130_fd_sc_hd__clkbuf_8
Xfanout398 _06752_ vssd1 vssd1 vccd1 vccd1 net398 sky130_fd_sc_hd__clkbuf_8
Xclkbuf_leaf_55_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_55_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_154_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10530__A2 net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09749_ _04775_ _05570_ net352 vssd1 vssd1 vccd1 vccd1 _05691_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_97_934 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout837_X net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11055__C _06541_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12760_ net1376 vssd1 vssd1 vccd1 vccd1 _00524_ sky130_fd_sc_hd__inv_2
XFILLER_0_68_124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09684__B1 _04816_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_6_Left_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_154_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_1125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11711_ net1942 net281 net335 vssd1 vssd1 vccd1 vccd1 _01825_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12691_ net1261 vssd1 vssd1 vccd1 vccd1 _00455_ sky130_fd_sc_hd__inv_2
XFILLER_0_68_179 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14430_ clknet_leaf_119_wb_clk_i _02194_ _00795_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[784\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_166_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11642_ _06716_ net386 net349 net2562 vssd1 vssd1 vccd1 vccd1 _01890_ sky130_fd_sc_hd__a22o_1
XFILLER_0_83_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10046__A1 net10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10046__B2 team_03_WB.instance_to_wrap.CPU_DAT_O\[17\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14361_ clknet_leaf_155_wb_clk_i _02125_ _00726_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[715\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_42_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11573_ net2510 net484 _06799_ net514 vssd1 vssd1 vccd1 vccd1 _01954_ sky130_fd_sc_hd__a22o_1
XANTENNA__11794__A1 _06624_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput18 DAT_I[24] vssd1 vssd1 vccd1 vccd1 net18 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__07998__B1 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13312_ net1333 vssd1 vssd1 vccd1 vccd1 _01076_ sky130_fd_sc_hd__inv_2
XANTENNA_input80_A wbs_adr_i[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_2301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10524_ net142 net1034 net1026 net1746 vssd1 vssd1 vccd1 vccd1 _02586_ sky130_fd_sc_hd__a22o_1
Xinput29 DAT_I[5] vssd1 vssd1 vccd1 vccd1 net29 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_94_2312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14292_ clknet_leaf_124_wb_clk_i _02056_ _00657_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[646\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_761 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11498__S net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09739__B2 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13243_ net1367 vssd1 vssd1 vccd1 vccd1 _01007_ sky130_fd_sc_hd__inv_2
X_10455_ team_03_WB.instance_to_wrap.core.pc.current_pc\[5\] _06270_ net683 vssd1
+ vssd1 vccd1 vccd1 _02639_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_3062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_3073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11546__A1 net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08411__A1 net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13174_ net1257 vssd1 vssd1 vccd1 vccd1 _00938_ sky130_fd_sc_hd__inv_2
X_10386_ team_03_WB.instance_to_wrap.core.pc.current_pc\[18\] _06214_ net677 vssd1
+ vssd1 vccd1 vccd1 _02652_ sky130_fd_sc_hd__mux2_1
XANTENNA__07845__S0 net1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12125_ net1649 vssd1 vssd1 vccd1 vccd1 _02428_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__06973__A1 net1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08600__S net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12056_ _06622_ net2678 net358 vssd1 vssd1 vccd1 vccd1 _01490_ sky130_fd_sc_hd__mux2_1
XANTENNA__09923__C net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08175__B1 net1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_9__f_wb_clk_i_A clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11007_ net2060 net421 _06576_ net499 vssd1 vssd1 vccd1 vccd1 _02297_ sky130_fd_sc_hd__a22o_1
XFILLER_0_74_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10521__A2 net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07216__S net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10150__B _05990_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08478__A1 net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12958_ net1415 vssd1 vssd1 vccd1 vccd1 _00722_ sky130_fd_sc_hd__inv_2
XANTENNA__08836__A net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09675__B1 _02804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_3205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11909_ _06609_ net2593 net367 vssd1 vssd1 vccd1 vccd1 _01633_ sky130_fd_sc_hd__mux2_1
XANTENNA__08573__S1 net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_3216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10824__A3 net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12889_ net1359 vssd1 vssd1 vccd1 vccd1 _00653_ sky130_fd_sc_hd__inv_2
XANTENNA__07150__A1 net1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_103_2485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_2496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14628_ clknet_leaf_21_wb_clk_i _02392_ _00993_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[982\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__12026__A2 net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_155_3552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_155_3563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07438__C1 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14559_ clknet_leaf_167_wb_clk_i _02323_ _00924_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[913\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_16_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10588__A2 net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_903 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07100_ _03039_ _03040_ _03041_ net1118 vssd1 vssd1 vccd1 vccd1 _03042_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_55_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_99_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07739__X _03681_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08080_ _04019_ _04021_ net1163 vssd1 vssd1 vccd1 vccd1 _04022_ sky130_fd_sc_hd__o21a_1
XFILLER_0_99_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07031_ team_03_WB.instance_to_wrap.core.decoder.inst\[23\] _02961_ _02972_ net718
+ vssd1 vssd1 vccd1 vccd1 _02973_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_114_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11201__S net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08938__C1 net1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11537__B2 net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08402__A1 net1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07610__C1 net1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08982_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[42\] net960
+ vssd1 vssd1 vccd1 vccd1 _04924_ sky130_fd_sc_hd__or2_1
XANTENNA__12821__A net1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_143_Right_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07933_ net743 _03873_ _03874_ net807 vssd1 vssd1 vccd1 vccd1 _03875_ sky130_fd_sc_hd__a31o_1
XANTENNA__08166__B1 net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07864_ net820 _03804_ _03805_ _03797_ _03800_ vssd1 vssd1 vccd1 vccd1 _03806_ sky130_fd_sc_hd__a32o_1
XANTENNA__07064__S1 net1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10512__A2 net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09603_ _04828_ _05460_ net572 vssd1 vssd1 vccd1 vccd1 _05545_ sky130_fd_sc_hd__mux2_2
XTAP_TAPCELL_ROW_127_2975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07795_ _03735_ _03736_ vssd1 vssd1 vccd1 vccd1 _03737_ sky130_fd_sc_hd__and2_1
XANTENNA__11871__S net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09115__C1 net1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout365_A _06815_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_30_wb_clk_i_A clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09534_ _04536_ _04777_ _05475_ vssd1 vssd1 vccd1 vccd1 _05476_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_27_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09465_ _05405_ _05406_ net554 vssd1 vssd1 vccd1 vccd1 _05407_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout532_A net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07141__A1 net1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_171_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_148_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08416_ net933 _04356_ _04357_ vssd1 vssd1 vccd1 vccd1 _04358_ sky130_fd_sc_hd__o21a_1
XFILLER_0_164_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12017__A2 net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09396_ _05331_ _05335_ _05337_ vssd1 vssd1 vccd1 vccd1 _05338_ sky130_fd_sc_hd__o21ai_4
XANTENNA__07692__A2 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_173_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_173_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_164_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout320_X net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08347_ net1234 team_03_WB.instance_to_wrap.core.register_file.registers_state\[469\]
+ net968 team_03_WB.instance_to_wrap.core.register_file.registers_state\[501\] net1212
+ vssd1 vssd1 vccd1 vccd1 _04289_ sky130_fd_sc_hd__o221a_1
XFILLER_0_163_357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1062_X net1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout418_X net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10579__A2 net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07796__S net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_102_wb_clk_i clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_102_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_08278_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[439\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[407\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[311\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[279\]
+ net963 net1072 vssd1 vssd1 vccd1 vccd1 _04220_ sky130_fd_sc_hd__mux4_1
XFILLER_0_85_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout999_A net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07229_ net1096 team_03_WB.instance_to_wrap.core.register_file.registers_state\[936\]
+ net896 vssd1 vssd1 vccd1 vccd1 _03171_ sky130_fd_sc_hd__or3_1
XFILLER_0_46_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11528__A1 net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11111__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_720 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10240_ _03944_ _05998_ vssd1 vssd1 vccd1 vccd1 _06082_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_132_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout787_X net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10171_ _06010_ _06011_ _03758_ vssd1 vssd1 vccd1 vccd1 _06013_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_121_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06955__A1 net1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_110_Right_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1105 _02787_ vssd1 vssd1 vccd1 vccd1 net1105 sky130_fd_sc_hd__buf_2
XANTENNA__07825__A net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1116 net1117 vssd1 vssd1 vccd1 vccd1 net1116 sky130_fd_sc_hd__buf_4
Xfanout1127 _02785_ vssd1 vssd1 vccd1 vccd1 net1127 sky130_fd_sc_hd__clkbuf_4
Xfanout1138 net1141 vssd1 vssd1 vccd1 vccd1 net1138 sky130_fd_sc_hd__buf_6
XANTENNA__08157__B1 net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1149 net1151 vssd1 vssd1 vccd1 vccd1 net1149 sky130_fd_sc_hd__buf_4
X_13930_ clknet_leaf_2_wb_clk_i _01694_ _00295_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[284\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11347__A net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07904__B1 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11066__B net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13861_ clknet_leaf_10_wb_clk_i _01625_ _00226_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[215\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_87_2160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09106__C1 net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11781__S net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12812_ net1333 vssd1 vssd1 vccd1 vccd1 _00576_ sky130_fd_sc_hd__inv_2
X_13792_ clknet_leaf_190_wb_clk_i _01556_ _00157_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[146\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_466 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07668__C1 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08555__S1 net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12743_ net1369 vssd1 vssd1 vccd1 vccd1 _00507_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_83_2079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_319 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07132__A1 net1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11082__A net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12008__A2 net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12674_ net1360 vssd1 vssd1 vccd1 vccd1 _00438_ sky130_fd_sc_hd__inv_2
XFILLER_0_60_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_61_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_398 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11216__A0 net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14413_ clknet_leaf_188_wb_clk_i _02177_ _00778_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[767\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_166_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11625_ _06699_ net379 net346 net2345 vssd1 vssd1 vccd1 vccd1 _01907_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_133_3102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_4_12__f_wb_clk_i_X clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_108_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12906__A net1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_3113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_536 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14344_ clknet_leaf_17_wb_clk_i _02108_ _00709_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[698\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07435__A2 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11556_ net491 net620 _06666_ net482 net1720 vssd1 vssd1 vccd1 vccd1 _01964_ sky130_fd_sc_hd__a32o_1
XANTENNA__08632__A1 net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06904__A net1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08391__A net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10507_ team_03_WB.instance_to_wrap.wb.curr_state\[1\] _02797_ team_03_WB.instance_to_wrap.wb.curr_state\[2\]
+ vssd1 vssd1 vccd1 vccd1 _06286_ sky130_fd_sc_hd__and3b_4
XFILLER_0_122_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_150_3460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14275_ clknet_leaf_34_wb_clk_i _02039_ _00640_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[629\]
+ sky130_fd_sc_hd__dfrtp_1
X_11487_ net2591 net394 _06777_ net514 vssd1 vssd1 vccd1 vccd1 _02018_ sky130_fd_sc_hd__a22o_1
XANTENNA__10990__A2 net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13226_ net1284 vssd1 vssd1 vccd1 vccd1 _00990_ sky130_fd_sc_hd__inv_2
X_10438_ team_03_WB.instance_to_wrap.core.pc.current_pc\[8\] _06136_ vssd1 vssd1 vccd1
+ vccd1 _06257_ sky130_fd_sc_hd__nor2_1
XFILLER_0_123_799 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_59_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11809__X _06811_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13157_ net1348 vssd1 vssd1 vccd1 vccd1 _00921_ sky130_fd_sc_hd__inv_2
X_10369_ net282 _06146_ _06197_ net677 vssd1 vssd1 vccd1 vccd1 _06201_ sky130_fd_sc_hd__o31a_1
XFILLER_0_0_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06946__B2 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12108_ net1145 net606 _06300_ net1578 _02765_ vssd1 vssd1 vccd1 vccd1 _00001_ sky130_fd_sc_hd__a32o_1
XANTENNA__08330__S net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13088_ net1402 vssd1 vssd1 vccd1 vccd1 _00852_ sky130_fd_sc_hd__inv_2
XFILLER_0_109_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11257__A net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12039_ _06777_ net480 net361 net2428 vssd1 vssd1 vccd1 vccd1 _01506_ sky130_fd_sc_hd__a22o_1
XANTENNA__08699__A1 net1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_69_Left_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09360__A2 _05281_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07371__A1 team_03_WB.instance_to_wrap.core.decoder.inst\[28\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_2525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07580_ net1092 team_03_WB.instance_to_wrap.core.register_file.registers_state\[824\]
+ net895 vssd1 vssd1 vccd1 vccd1 _03522_ sky130_fd_sc_hd__or3_1
XFILLER_0_88_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_157_3603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07470__A net1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11455__B1 net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_2872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07123__A1 net1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_2883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_0_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_47_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_114_wb_clk_i_A clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_29_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09250_ _05190_ _05191_ vssd1 vssd1 vccd1 vccd1 _05192_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_174_3950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_174_3961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08201_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[947\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[915\]
+ net957 vssd1 vssd1 vccd1 vccd1 _04143_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11207__A0 _06438_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_174_3972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_145_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_146_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09668__Y _05610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09181_ net552 _04807_ _05121_ _05122_ vssd1 vssd1 vccd1 vccd1 _05123_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_56_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_173_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08132_ _03208_ _03243_ _03759_ _03790_ vssd1 vssd1 vccd1 vccd1 _04074_ sky130_fd_sc_hd__and4b_1
XPHY_EDGE_ROW_78_Left_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_170_3858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08623__A1 net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_wire588_X net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_170_3869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_95 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08063_ net1130 _04000_ _04001_ _04003_ net1116 vssd1 vssd1 vccd1 vccd1 _04005_ sky130_fd_sc_hd__a311o_1
XFILLER_0_144_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_964 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_141_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09179__A2 _04807_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07014_ net1196 team_03_WB.instance_to_wrap.core.register_file.registers_state\[995\]
+ net883 _02955_ vssd1 vssd1 vccd1 vccd1 _02956_ sky130_fd_sc_hd__a31o_1
XFILLER_0_101_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10733__A2 net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08965_ net1223 _04905_ _04906_ vssd1 vssd1 vccd1 vccd1 _04907_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout482_A _06779_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11167__A _06562_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07916_ net1200 team_03_WB.instance_to_wrap.core.register_file.registers_state\[943\]
+ net878 _02870_ vssd1 vssd1 vccd1 vccd1 _03858_ sky130_fd_sc_hd__a31o_1
XPHY_EDGE_ROW_87_Left_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08896_ _04836_ _04837_ net863 vssd1 vssd1 vccd1 vccd1 _04838_ sky130_fd_sc_hd__a21o_1
XANTENNA_clkbuf_leaf_153_wb_clk_i_A clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09860__A _05706_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07847_ team_03_WB.instance_to_wrap.core.decoder.inst\[30\] net826 vssd1 vssd1 vccd1
+ vccd1 _03789_ sky130_fd_sc_hd__nand2_1
XANTENNA__11694__B1 net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout747_A net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout368_X net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_4_8__f_wb_clk_i_X clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_07778_ net731 _03708_ _03709_ _03707_ net809 vssd1 vssd1 vccd1 vccd1 _03720_ sky130_fd_sc_hd__a311o_1
XANTENNA__07380__A net1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09517_ net561 _05380_ _05458_ vssd1 vssd1 vccd1 vccd1 _05459_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_39_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout914_A net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11106__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08311__B1 net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09448_ net594 _05340_ vssd1 vssd1 vccd1 vccd1 _05390_ sky130_fd_sc_hd__nor2_1
XANTENNA__11333__C net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07665__A2 net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_163_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_163_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_96_Left_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_163_132 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09379_ _05315_ _05320_ vssd1 vssd1 vccd1 vccd1 _05321_ sky130_fd_sc_hd__and2_1
XFILLER_0_34_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout702_X net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11749__A1 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11410_ net274 net2473 net396 vssd1 vssd1 vccd1 vccd1 _02070_ sky130_fd_sc_hd__mux2_1
XFILLER_0_164_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_176 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08614__A1 net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12390_ net1337 vssd1 vssd1 vccd1 vccd1 _00154_ sky130_fd_sc_hd__inv_2
X_11341_ net302 net711 net696 vssd1 vssd1 vccd1 vccd1 _06723_ sky130_fd_sc_hd__and3_1
XFILLER_0_34_399 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14060_ clknet_leaf_16_wb_clk_i _01824_ _00425_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[414\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_160_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11272_ net508 net637 _06703_ net410 net2188 vssd1 vssd1 vccd1 vccd1 _02159_ sky130_fd_sc_hd__a32o_1
X_13011_ net1255 vssd1 vssd1 vccd1 vccd1 _00775_ sky130_fd_sc_hd__inv_2
X_10223_ _06017_ _06021_ _06062_ _06016_ _06013_ vssd1 vssd1 vccd1 vccd1 _06065_ sky130_fd_sc_hd__a311o_2
XANTENNA_clkbuf_leaf_192_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_70_wb_clk_i clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_70_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_input43_A gpio_in[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10154_ _05995_ vssd1 vssd1 vccd1 vccd1 _05996_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_89_2200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_2211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14962_ clknet_leaf_95_wb_clk_i _02714_ _01327_ vssd1 vssd1 vccd1 vccd1 net214 sky130_fd_sc_hd__dfrtp_1
X_10085_ _05757_ _05926_ net318 vssd1 vssd1 vccd1 vccd1 _05929_ sky130_fd_sc_hd__and3b_1
Xhold7 team_03_WB.instance_to_wrap.core.register_file.registers_state\[27\] vssd1
+ vssd1 vccd1 vccd1 net1500 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10488__A1 net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13913_ clknet_leaf_169_wb_clk_i _01677_ _00278_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[267\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11685__B1 net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07889__C1 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14893_ clknet_leaf_60_wb_clk_i _02656_ _01258_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.pc.current_pc\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_50_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13844_ clknet_leaf_132_wb_clk_i _01608_ _00209_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[198\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_71_17 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07290__A net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_18_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11524__B net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13775_ clknet_leaf_144_wb_clk_i _01539_ _00140_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[129\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10987_ net281 net646 net703 net827 vssd1 vssd1 vccd1 vccd1 _06565_ sky130_fd_sc_hd__and4_1
XANTENNA__07105__A1 net1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_100_2422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12726_ net1258 vssd1 vssd1 vccd1 vccd1 _00490_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_100_2433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11243__C net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10660__A1 team_03_WB.instance_to_wrap.CPU_DAT_O\[1\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_66_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_152_3500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12657_ net1273 vssd1 vssd1 vccd1 vccd1 _00421_ sky130_fd_sc_hd__inv_2
XANTENNA__09929__B net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_142_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11608_ net653 net464 vssd1 vssd1 vccd1 vccd1 _06802_ sky130_fd_sc_hd__and2_1
XFILLER_0_81_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_167_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12588_ net1310 vssd1 vssd1 vccd1 vccd1 _00352_ sky130_fd_sc_hd__inv_2
XFILLER_0_25_355 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09010__A net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10412__A1 net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14327_ clknet_leaf_79_wb_clk_i _02091_ _00692_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[681\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08700__S1 net1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11539_ net2093 net483 _06787_ net498 vssd1 vssd1 vccd1 vccd1 _01976_ sky130_fd_sc_hd__a22o_1
Xhold407 team_03_WB.instance_to_wrap.core.register_file.registers_state\[563\] vssd1
+ vssd1 vccd1 vccd1 net1900 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold418 team_03_WB.instance_to_wrap.core.register_file.registers_state\[744\] vssd1
+ vssd1 vccd1 vccd1 net1911 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_151_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09945__A _03425_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_347 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold429 net198 vssd1 vssd1 vccd1 vccd1 net1922 sky130_fd_sc_hd__dlygate4sd3_1
X_14258_ clknet_leaf_168_wb_clk_i _02022_ _00623_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[612\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_78_1970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06921__X _02863_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_1981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13209_ net1355 vssd1 vssd1 vccd1 vccd1 _00973_ sky130_fd_sc_hd__inv_2
XANTENNA__09030__A1 net1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14189_ clknet_leaf_182_wb_clk_i _01953_ _00554_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[543\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout909 net910 vssd1 vssd1 vccd1 vccd1 net909 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_0_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07041__B1 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_1889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08750_ net1065 _04690_ _04691_ vssd1 vssd1 vccd1 vccd1 _04692_ sky130_fd_sc_hd__a21o_1
Xhold1107 team_03_WB.instance_to_wrap.core.register_file.registers_state\[467\] vssd1
+ vssd1 vccd1 vccd1 net2600 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1118 team_03_WB.instance_to_wrap.core.register_file.registers_state\[118\] vssd1
+ vssd1 vccd1 vccd1 net2611 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1129 team_03_WB.instance_to_wrap.core.register_file.registers_state\[670\] vssd1
+ vssd1 vccd1 vccd1 net2622 sky130_fd_sc_hd__dlygate4sd3_1
X_07701_ net1195 team_03_WB.instance_to_wrap.core.register_file.registers_state\[45\]
+ net882 vssd1 vssd1 vccd1 vccd1 _03643_ sky130_fd_sc_hd__and3_1
XFILLER_0_136_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_124_2912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08681_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[744\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[712\]
+ net975 vssd1 vssd1 vccd1 vccd1 _04623_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_124_2923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07344__A1 net1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07632_ net1192 team_03_WB.instance_to_wrap.core.register_file.registers_state\[110\]
+ net881 _03573_ vssd1 vssd1 vccd1 vccd1 _03574_ sky130_fd_sc_hd__a31o_1
XFILLER_0_136_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11428__B1 net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07563_ net1130 _03501_ _03502_ net1117 vssd1 vssd1 vccd1 vccd1 _03505_ sky130_fd_sc_hd__a211oi_1
X_09302_ _04591_ _05243_ vssd1 vssd1 vccd1 vccd1 _05244_ sky130_fd_sc_hd__and2_1
XFILLER_0_152_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_447 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_172_3909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07494_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[679\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[647\]
+ net785 vssd1 vssd1 vccd1 vccd1 _03436_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_266 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09233_ _03904_ _05156_ vssd1 vssd1 vccd1 vccd1 _05175_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10651__A1 team_03_WB.instance_to_wrap.CPU_DAT_O\[10\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10765__S net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12546__A net1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_146_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout328_A _06810_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11450__A net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_161_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09164_ net563 _05105_ _05100_ vssd1 vssd1 vccd1 vccd1 _05106_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_160_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_161_647 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_675 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08115_ _04050_ _04051_ _04056_ net1160 vssd1 vssd1 vccd1 vccd1 _04057_ sky130_fd_sc_hd__o22a_1
XANTENNA__10403__B2 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07804__C1 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10066__A team_03_WB.instance_to_wrap.core.decoder.inst\[31\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09095_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[1005\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[973\]
+ net989 vssd1 vssd1 vccd1 vccd1 _05037_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout1237_A net1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08046_ _03986_ _03987_ vssd1 vssd1 vccd1 vccd1 _03988_ sky130_fd_sc_hd__nor2_2
Xclkbuf_4_2__f_wb_clk_i clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_2__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__07280__B1 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold930 team_03_WB.instance_to_wrap.core.register_file.registers_state\[102\] vssd1
+ vssd1 vccd1 vccd1 net2423 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold941 team_03_WB.instance_to_wrap.core.register_file.registers_state\[799\] vssd1
+ vssd1 vccd1 vccd1 net2434 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11596__S net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout697_A net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold952 team_03_WB.instance_to_wrap.core.register_file.registers_state\[207\] vssd1
+ vssd1 vccd1 vccd1 net2445 sky130_fd_sc_hd__dlygate4sd3_1
Xhold963 team_03_WB.instance_to_wrap.core.register_file.registers_state\[150\] vssd1
+ vssd1 vccd1 vccd1 net2456 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09021__A1 net1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1404_A net1408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold974 team_03_WB.instance_to_wrap.core.register_file.registers_state\[222\] vssd1
+ vssd1 vccd1 vccd1 net2467 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1025_X net1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11903__A1 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold985 team_03_WB.instance_to_wrap.core.register_file.registers_state\[815\] vssd1
+ vssd1 vccd1 vccd1 net2478 sky130_fd_sc_hd__dlygate4sd3_1
Xhold996 team_03_WB.instance_to_wrap.core.register_file.registers_state\[501\] vssd1
+ vssd1 vccd1 vccd1 net2489 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11609__B net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09997_ _05882_ net1786 net287 vssd1 vssd1 vccd1 vccd1 _02717_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout485_X net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout864_A net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07583__A1 net1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08780__B1 net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08948_ net924 _04887_ _04888_ net862 vssd1 vssd1 vccd1 vccd1 _04890_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_32_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08879_ _02944_ _02947_ vssd1 vssd1 vccd1 vccd1 _04821_ sky130_fd_sc_hd__nand2b_1
XANTENNA_fanout652_X net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10910_ net692 _05676_ net586 vssd1 vssd1 vccd1 vccd1 _06500_ sky130_fd_sc_hd__o21ai_1
X_11890_ net624 _06699_ net455 net371 net1923 vssd1 vssd1 vccd1 vccd1 _01651_ sky130_fd_sc_hd__a32o_1
XANTENNA__11419__A0 _06499_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10841_ _06439_ _06440_ _06441_ net586 vssd1 vssd1 vccd1 vccd1 _06442_ sky130_fd_sc_hd__o211a_2
XANTENNA__10890__A1 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_2016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout917_X net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_2027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13560_ net1407 vssd1 vssd1 vccd1 vccd1 _01324_ sky130_fd_sc_hd__inv_2
XANTENNA__12092__B1 net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10772_ team_03_WB.instance_to_wrap.core.decoder.inst\[10\] net1248 vssd1 vssd1 vccd1
+ vccd1 _06382_ sky130_fd_sc_hd__nand2_1
XANTENNA__08934__A net1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12511_ net1287 vssd1 vssd1 vccd1 vccd1 _00275_ sky130_fd_sc_hd__inv_2
XFILLER_0_66_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13491_ net1327 vssd1 vssd1 vccd1 vccd1 _01255_ sky130_fd_sc_hd__inv_2
XFILLER_0_152_603 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08653__B net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12442_ net1378 vssd1 vssd1 vccd1 vccd1 _00206_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08599__B1 net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12373_ net1272 vssd1 vssd1 vccd1 vccd1 _00137_ sky130_fd_sc_hd__inv_2
XFILLER_0_133_872 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14112_ clknet_leaf_192_wb_clk_i _01876_ _00477_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[466\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_50_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11324_ _06629_ net2686 net407 vssd1 vssd1 vccd1 vccd1 _02121_ sky130_fd_sc_hd__mux2_1
X_15092_ net1478 vssd1 vssd1 vccd1 vccd1 la_data_out[28] sky130_fd_sc_hd__buf_2
XFILLER_0_22_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14043_ clknet_leaf_159_wb_clk_i _01807_ _00408_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[397\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_56_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11255_ net275 net711 net828 vssd1 vssd1 vccd1 vccd1 _06695_ sky130_fd_sc_hd__and3_1
XFILLER_0_120_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_128_3001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10206_ net592 net676 _06044_ _02994_ vssd1 vssd1 vccd1 vccd1 _06048_ sky130_fd_sc_hd__o211ai_1
XTAP_TAPCELL_ROW_128_3012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07285__A net1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11186_ net707 net269 net700 vssd1 vssd1 vccd1 vccd1 _06674_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_52_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11370__A2 net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10137_ _03528_ _05978_ vssd1 vssd1 vccd1 vccd1 _05979_ sky130_fd_sc_hd__nor2_1
X_14945_ clknet_leaf_56_wb_clk_i _00007_ _01310_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.wb.curr_state\[0\]
+ sky130_fd_sc_hd__dfstp_1
X_10068_ team_03_WB.instance_to_wrap.core.decoder.inst\[14\] team_03_WB.instance_to_wrap.core.decoder.inst\[13\]
+ team_03_WB.instance_to_wrap.core.decoder.inst\[12\] team_03_WB.instance_to_wrap.core.decoder.inst\[7\]
+ vssd1 vssd1 vccd1 vccd1 _05912_ sky130_fd_sc_hd__or4_1
XPHY_EDGE_ROW_13_Right_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_314 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08523__B1 net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_141_3267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_141_3278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14876_ clknet_leaf_89_wb_clk_i _02639_ _01241_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.pc.current_pc\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_77_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07451__C net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09079__A1 net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13827_ clknet_leaf_30_wb_clk_i _01591_ _00192_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[181\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_134_1097 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08826__A1 net1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13758_ clknet_leaf_118_wb_clk_i _01522_ _00123_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[112\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12083__B1 net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08844__A net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12709_ net1354 vssd1 vssd1 vccd1 vccd1 _00473_ sky130_fd_sc_hd__inv_2
XFILLER_0_17_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11830__B1 net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13689_ clknet_leaf_168_wb_clk_i _01453_ _00054_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[43\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08563__B net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_142_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_22_Right_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_984 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_117_2771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_2782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold204 _02591_ vssd1 vssd1 vccd1 vccd1 net1697 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_360 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_1929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold215 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[31\] vssd1 vssd1 vccd1
+ vccd1 net1708 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07262__B1 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07801__A2 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold226 _02584_ vssd1 vssd1 vccd1 vccd1 net1719 sky130_fd_sc_hd__dlygate4sd3_1
Xhold237 _02601_ vssd1 vssd1 vccd1 vccd1 net1730 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold248 net187 vssd1 vssd1 vccd1 vccd1 net1741 sky130_fd_sc_hd__dlygate4sd3_1
X_09920_ _05847_ _05596_ _05583_ vssd1 vssd1 vccd1 vccd1 _05862_ sky130_fd_sc_hd__nor3b_1
XFILLER_0_150_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold259 _02527_ vssd1 vssd1 vccd1 vccd1 net1752 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09003__A1 net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_764 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout706 net708 vssd1 vssd1 vccd1 vccd1 net706 sky130_fd_sc_hd__buf_2
X_09851_ net561 _05136_ vssd1 vssd1 vccd1 vccd1 _05793_ sky130_fd_sc_hd__nor2_1
Xfanout717 net720 vssd1 vssd1 vccd1 vccd1 net717 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_1_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08211__C1 net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11897__B1 net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout728 net729 vssd1 vssd1 vccd1 vccd1 net728 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_165_3757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07626__C net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_165_3768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout739 net740 vssd1 vssd1 vccd1 vccd1 net739 sky130_fd_sc_hd__buf_4
XANTENNA__07565__A1 net1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08802_ _04742_ _04743_ net857 vssd1 vssd1 vccd1 vccd1 _04744_ sky130_fd_sc_hd__o21a_1
X_09782_ net578 _05638_ _05723_ net353 vssd1 vssd1 vccd1 vccd1 _05724_ sky130_fd_sc_hd__o211a_1
X_06994_ team_03_WB.instance_to_wrap.core.decoder.inst\[13\] _02832_ _02925_ _02927_
+ vssd1 vssd1 vccd1 vccd1 _02936_ sky130_fd_sc_hd__nor4_1
XPHY_EDGE_ROW_31_Right_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11148__C net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08733_ net1050 team_03_WB.instance_to_wrap.core.register_file.registers_state\[836\]
+ net1002 team_03_WB.instance_to_wrap.core.register_file.registers_state\[868\] net1067
+ vssd1 vssd1 vccd1 vccd1 _04675_ sky130_fd_sc_hd__a221o_1
XANTENNA__07923__A net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10987__C net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout278_A _06426_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08664_ net1068 _04604_ _04605_ vssd1 vssd1 vccd1 vccd1 _04606_ sky130_fd_sc_hd__a21o_1
XFILLER_0_163_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_152_1131 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07615_ net1205 team_03_WB.instance_to_wrap.core.register_file.registers_state\[569\]
+ net886 vssd1 vssd1 vccd1 vccd1 _03557_ sky130_fd_sc_hd__and3_1
XANTENNA__11164__B net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10872__A1 net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08595_ _04327_ _04536_ _02992_ vssd1 vssd1 vccd1 vccd1 _04537_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout445_A net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1187_A net1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12074__B1 net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07546_ net718 _03471_ _03480_ _03487_ vssd1 vssd1 vccd1 vccd1 _03488_ sky130_fd_sc_hd__o22a_4
XFILLER_0_76_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08817__A1 net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_290 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09202__X _05144_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10624__A1 team_03_WB.instance_to_wrap.CPU_DAT_O\[5\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11821__B1 net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07477_ _03417_ _03418_ net1162 vssd1 vssd1 vccd1 vccd1 _03419_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_5_1070 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07096__A3 net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_40_Right_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1354_A net1358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_631 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_162_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09216_ net607 _03529_ _05157_ vssd1 vssd1 vccd1 vccd1 _05158_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_8_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_176 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_945 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_173_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_984 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09147_ _05087_ _05088_ vssd1 vssd1 vccd1 vccd1 _05089_ sky130_fd_sc_hd__nor2_1
XFILLER_0_72_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout400_X net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08676__S0 net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10927__A2 _05718_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07253__B1 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09078_ net857 _05018_ _05019_ vssd1 vssd1 vccd1 vccd1 _05020_ sky130_fd_sc_hd__or3_1
XFILLER_0_114_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout981_A net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08029_ net742 _03969_ _03970_ net806 vssd1 vssd1 vccd1 vccd1 _03971_ sky130_fd_sc_hd__a31o_1
Xhold760 team_03_WB.instance_to_wrap.core.register_file.registers_state\[244\] vssd1
+ vssd1 vccd1 vccd1 net2253 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold771 team_03_WB.instance_to_wrap.core.register_file.registers_state\[801\] vssd1
+ vssd1 vccd1 vccd1 net2264 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold782 team_03_WB.instance_to_wrap.core.register_file.registers_state\[598\] vssd1
+ vssd1 vccd1 vccd1 net2275 sky130_fd_sc_hd__dlygate4sd3_1
X_11040_ net702 net714 net296 vssd1 vssd1 vccd1 vccd1 _06596_ sky130_fd_sc_hd__or3b_1
XANTENNA__11888__B1 net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold793 team_03_WB.instance_to_wrap.core.register_file.registers_state\[700\] vssd1
+ vssd1 vccd1 vccd1 net2286 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11339__B net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout867_X net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07556__A1 net1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11352__A2 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10560__B1 net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12991_ net1349 vssd1 vssd1 vccd1 vccd1 _00755_ sky130_fd_sc_hd__inv_2
XANTENNA__07308__A1 net1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11355__A net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14730_ clknet_leaf_61_wb_clk_i _02494_ _01095_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.decoder.inst\[27\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_118_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11942_ net622 _06719_ net454 net363 net2687 vssd1 vssd1 vccd1 vccd1 _01601_ sky130_fd_sc_hd__a32o_1
XFILLER_0_19_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_1074 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_24_Left_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11074__B net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14661_ clknet_leaf_40_wb_clk_i _02425_ _01026_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1015\]
+ sky130_fd_sc_hd__dfstp_1
X_11873_ net267 net2078 net377 vssd1 vssd1 vccd1 vccd1 _01667_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_419 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13612_ net1303 vssd1 vssd1 vccd1 vccd1 _01376_ sky130_fd_sc_hd__inv_2
XFILLER_0_156_216 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10824_ net311 net310 net317 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[25\]
+ vssd1 vssd1 vccd1 vccd1 _06428_ sky130_fd_sc_hd__a31o_1
X_14592_ clknet_leaf_192_wb_clk_i _02356_ _00957_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[946\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__08808__A1 net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10076__C1 net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10615__A1 team_03_WB.instance_to_wrap.CPU_DAT_O\[14\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13543_ net1326 vssd1 vssd1 vccd1 vccd1 _01307_ sky130_fd_sc_hd__inv_2
XFILLER_0_138_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10755_ team_03_WB.instance_to_wrap.core.pc.current_pc\[5\] _05757_ net605 vssd1
+ vssd1 vccd1 vccd1 _06371_ sky130_fd_sc_hd__mux2_1
XANTENNA__11812__B1 net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_912 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13474_ net1431 vssd1 vssd1 vccd1 vccd1 _01238_ sky130_fd_sc_hd__inv_2
XFILLER_0_168_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10686_ _06319_ _06326_ net602 vssd1 vssd1 vccd1 vccd1 _06327_ sky130_fd_sc_hd__a21o_1
XANTENNA__08951__X _04893_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12425_ net1257 vssd1 vssd1 vccd1 vccd1 _00189_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_97_2365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_146 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_2376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12914__A net1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1132 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07244__B1 net1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09784__A2 _04619_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12356_ net1382 vssd1 vssd1 vccd1 vccd1 _00120_ sky130_fd_sc_hd__inv_2
XANTENNA__08603__S net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06912__A net1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11307_ _06617_ net2589 net404 vssd1 vssd1 vccd1 vccd1 _02138_ sky130_fd_sc_hd__mux2_1
X_15075_ net1461 vssd1 vssd1 vccd1 vccd1 la_data_out[11] sky130_fd_sc_hd__buf_2
XFILLER_0_26_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12287_ net1348 vssd1 vssd1 vccd1 vccd1 _00051_ sky130_fd_sc_hd__inv_2
XFILLER_0_22_199 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14026_ clknet_leaf_0_wb_clk_i _01790_ _00391_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[380\]
+ sky130_fd_sc_hd__dfrtp_1
X_11238_ net495 net630 _06686_ net408 net2363 vssd1 vssd1 vccd1 vccd1 _02176_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_71_1826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11249__B net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11879__B1 net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_1837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07547__A1 _03488_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08744__B1 net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_143_3307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_3318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11169_ net2288 net414 _06663_ net507 vssd1 vssd1 vccd1 vccd1 _02222_ sky130_fd_sc_hd__a22o_1
XFILLER_0_93_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11894__A3 net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_160_3654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_160_3665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11265__A net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14928_ clknet_leaf_50_wb_clk_i _02683_ _01293_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_O\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_117_77 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_69_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14859_ clknet_leaf_57_wb_clk_i net1565 _01224_ vssd1 vssd1 vccd1 vccd1 net115 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_69_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07400_ net1082 team_03_WB.instance_to_wrap.core.register_file.registers_state\[895\]
+ net888 vssd1 vssd1 vccd1 vccd1 _03342_ sky130_fd_sc_hd__or3_1
X_08380_ net867 _04321_ _04316_ vssd1 vssd1 vccd1 vccd1 _04322_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_92_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08574__A net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07331_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[445\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[413\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[317\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[285\]
+ net768 net1128 vssd1 vssd1 vccd1 vccd1 _03273_ sky130_fd_sc_hd__mux4_1
XFILLER_0_156_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_964 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_119_2811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_2822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11204__S net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07262_ net818 _03203_ net718 vssd1 vssd1 vccd1 vccd1 _03204_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_143_422 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09001_ net1218 _04941_ _04942_ net1070 vssd1 vssd1 vccd1 vccd1 _04943_ sky130_fd_sc_hd__o211a_1
XFILLER_0_42_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07193_ net1146 _03129_ _03134_ net817 vssd1 vssd1 vccd1 vccd1 _03135_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_14_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07235__B1 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11031__B2 net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08432__C1 net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_167_3808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07786__B2 _03726_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08983__B1 net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09903_ _05844_ _05455_ _05429_ _05542_ vssd1 vssd1 vccd1 vccd1 _05845_ sky130_fd_sc_hd__and4b_2
XFILLER_0_111_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_6_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout503 net504 vssd1 vssd1 vccd1 vccd1 net503 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11159__B net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout514 net516 vssd1 vssd1 vccd1 vccd1 net514 sky130_fd_sc_hd__buf_4
Xfanout525 _06322_ vssd1 vssd1 vccd1 vccd1 net525 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_6_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout536 net537 vssd1 vssd1 vccd1 vccd1 net536 sky130_fd_sc_hd__clkbuf_2
XANTENNA__11334__A2 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08735__B1 net1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11874__S net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout547 net548 vssd1 vssd1 vccd1 vccd1 net547 sky130_fd_sc_hd__clkbuf_4
X_09834_ net322 _05436_ _05775_ vssd1 vssd1 vccd1 vccd1 _05776_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_67_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_127_wb_clk_i clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_127_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xfanout558 _03064_ vssd1 vssd1 vccd1 vccd1 net558 sky130_fd_sc_hd__buf_2
XANTENNA__06968__S net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1102_A net1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout569 _03024_ vssd1 vssd1 vccd1 vccd1 net569 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08749__A net1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11885__A3 net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09765_ _05239_ _05271_ _05273_ vssd1 vssd1 vccd1 vccd1 _05707_ sky130_fd_sc_hd__a21oi_1
X_06977_ _02914_ _02915_ net808 vssd1 vssd1 vccd1 vccd1 _02919_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout562_A _03063_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11175__A net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08716_ net1047 team_03_WB.instance_to_wrap.core.register_file.registers_state\[324\]
+ net999 team_03_WB.instance_to_wrap.core.register_file.registers_state\[356\] net1216
+ vssd1 vssd1 vccd1 vccd1 _04658_ sky130_fd_sc_hd__a221o_1
X_09696_ _04150_ _04326_ _05014_ _04210_ net562 net571 vssd1 vssd1 vccd1 vccd1 _05638_
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_68_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08647_ _04587_ _04588_ vssd1 vssd1 vccd1 vccd1 _04589_ sky130_fd_sc_hd__and2_1
XANTENNA__07171__C1 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07710__A1 net1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1092_X net1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout448_X net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout827_A net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12047__A0 _06616_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08578_ net1235 team_03_WB.instance_to_wrap.core.register_file.registers_state\[733\]
+ net966 team_03_WB.instance_to_wrap.core.register_file.registers_state\[765\] net937
+ vssd1 vssd1 vccd1 vccd1 _04520_ sky130_fd_sc_hd__o221a_1
XFILLER_0_7_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_166_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07529_ _03463_ _03464_ _03469_ _03470_ net1122 net1139 vssd1 vssd1 vccd1 vccd1 _03471_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_76_383 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout615_X net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11114__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10540_ net171 net1027 net905 net1495 vssd1 vssd1 vccd1 vccd1 _02570_ sky130_fd_sc_hd__a22o_1
XANTENNA__07474__B1 net1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11270__A1 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11341__C net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08671__C1 net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10471_ net1143 net2154 _06282_ vssd1 vssd1 vccd1 vccd1 _02635_ sky130_fd_sc_hd__o21a_1
XPHY_EDGE_ROW_157_Right_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10806__X _06414_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_168 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12210_ net1525 vssd1 vssd1 vccd1 vccd1 _02343_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_40_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13190_ net1301 vssd1 vssd1 vccd1 vccd1 _00954_ sky130_fd_sc_hd__inv_2
XANTENNA__07777__A1 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout984_X net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11573__A2 net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14722__Q team_03_WB.instance_to_wrap.core.decoder.inst\[19\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12141_ net1597 vssd1 vssd1 vccd1 vccd1 _02412_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_103_864 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_2262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10254__A _03901_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_2273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12072_ _06633_ net2682 net357 vssd1 vssd1 vccd1 vccd1 _01474_ sky130_fd_sc_hd__mux2_1
Xhold590 team_03_WB.instance_to_wrap.core.register_file.registers_state\[758\] vssd1
+ vssd1 vccd1 vccd1 net2083 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11784__S net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08726__B1 net999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11023_ net511 net656 _06585_ net423 net1847 vssd1 vssd1 vccd1 vccd1 _02290_ sky130_fd_sc_hd__a32o_1
XANTENNA__10533__B1 net1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11876__A3 net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_32_Left_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12974_ net1303 vssd1 vssd1 vccd1 vccd1 _00738_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1290 team_03_WB.instance_to_wrap.CPU_DAT_O\[26\] vssd1 vssd1 vccd1 vccd1 net2783
+ sky130_fd_sc_hd__dlygate4sd3_1
X_14713_ clknet_leaf_47_wb_clk_i _02477_ _01078_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.decoder.inst\[10\]
+ sky130_fd_sc_hd__dfrtp_4
X_11925_ _06623_ net2445 net368 vssd1 vssd1 vccd1 vccd1 _01617_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_339 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07162__C1 net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output112_A net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12038__B1 net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11856_ net273 net2173 net375 vssd1 vssd1 vccd1 vccd1 _01684_ sky130_fd_sc_hd__mux2_1
X_14644_ clknet_leaf_132_wb_clk_i _02408_ _01009_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[998\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_170_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_1034 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06907__A net1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_2405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10807_ _06413_ net2206 net519 vssd1 vssd1 vccd1 vccd1 _02335_ sky130_fd_sc_hd__mux2_1
XANTENNA__11532__B net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_2416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14575_ clknet_leaf_135_wb_clk_i _02339_ _00940_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[929\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11787_ net2495 _06620_ net327 vssd1 vssd1 vccd1 vccd1 _01751_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_219 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10738_ team_03_WB.instance_to_wrap.core.pc.current_pc\[12\] _05697_ net605 vssd1
+ vssd1 vccd1 vccd1 _06361_ sky130_fd_sc_hd__mux2_1
X_13526_ net1316 vssd1 vssd1 vccd1 vccd1 _01290_ sky130_fd_sc_hd__inv_2
XANTENNA__07465__B1 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11251__C net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_136_3166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_504 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_3177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_41_Left_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13457_ net1341 vssd1 vssd1 vccd1 vccd1 _01221_ sky130_fd_sc_hd__inv_2
XFILLER_0_36_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09937__B net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10669_ _05455_ _06310_ vssd1 vssd1 vccd1 vccd1 _06311_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_124_Right_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_140_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_274 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12408_ net1374 vssd1 vssd1 vccd1 vccd1 _00172_ sky130_fd_sc_hd__inv_2
XANTENNA__09757__A2 _04922_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07738__A net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08333__S net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13388_ net1421 vssd1 vssd1 vccd1 vccd1 _01152_ sky130_fd_sc_hd__inv_2
Xoutput106 net106 vssd1 vssd1 vccd1 vccd1 ADR_O[12] sky130_fd_sc_hd__clkbuf_4
Xoutput117 net117 vssd1 vssd1 vccd1 vccd1 ADR_O[22] sky130_fd_sc_hd__clkbuf_4
XANTENNA__11564__A2 net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput128 net128 vssd1 vssd1 vccd1 vccd1 ADR_O[3] sky130_fd_sc_hd__clkbuf_4
X_12339_ net1255 vssd1 vssd1 vccd1 vccd1 _00103_ sky130_fd_sc_hd__inv_2
XANTENNA__10164__A _03724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput139 net139 vssd1 vssd1 vccd1 vccd1 DAT_O[12] sky130_fd_sc_hd__buf_2
XFILLER_0_50_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_110_2627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_2638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15058_ net1444 vssd1 vssd1 vccd1 vccd1 gpio_out[4] sky130_fd_sc_hd__buf_2
XANTENNA__09953__A _03984_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08717__B1 net999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_162_3705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06900_ net1022 _02834_ _02838_ _02841_ vssd1 vssd1 vccd1 vccd1 _02842_ sky130_fd_sc_hd__nor4_1
X_14009_ clknet_leaf_155_wb_clk_i _01773_ _00374_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[363\]
+ sky130_fd_sc_hd__dfrtp_1
X_07880_ team_03_WB.instance_to_wrap.core.decoder.inst\[27\] net1019 net684 vssd1
+ vssd1 vccd1 vccd1 _03822_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_49_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10524__B1 net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08569__A net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_50_Left_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06831_ team_03_WB.instance_to_wrap.core.pc.current_pc\[3\] vssd1 vssd1 vccd1 vccd1
+ _02774_ sky130_fd_sc_hd__inv_2
X_09550_ _03529_ _04267_ net535 _05491_ _03527_ vssd1 vssd1 vccd1 vccd1 _05492_ sky130_fd_sc_hd__o311a_1
XANTENNA_clkbuf_leaf_20_wb_clk_i_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09142__A0 net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08501_ _04437_ _04442_ net874 vssd1 vssd1 vccd1 vccd1 _04443_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_108_2589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09481_ _03641_ _04503_ net538 vssd1 vssd1 vccd1 vccd1 _05423_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_53_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07153__C1 net1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08432_ net937 _04373_ _04372_ net1063 vssd1 vssd1 vccd1 vccd1 _04374_ sky130_fd_sc_hd__o211a_1
XFILLER_0_77_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12029__B1 net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08363_ net1236 team_03_WB.instance_to_wrap.core.register_file.registers_state\[470\]
+ net970 team_03_WB.instance_to_wrap.core.register_file.registers_state\[502\] net1212
+ vssd1 vssd1 vccd1 vccd1 _04305_ sky130_fd_sc_hd__o221a_1
XFILLER_0_92_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_528 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_160_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_260 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07314_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[541\] net768
+ net743 _03255_ vssd1 vssd1 vccd1 vccd1 _03256_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_22_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11252__A1 net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08294_ _04235_ vssd1 vssd1 vccd1 vccd1 _04236_ sky130_fd_sc_hd__inv_2
XFILLER_0_73_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_160_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11869__S net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07245_ net1139 _03181_ _03182_ _03185_ _03186_ vssd1 vssd1 vccd1 vccd1 _03187_ sky130_fd_sc_hd__o32a_1
XANTENNA_fanout310_A _05845_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1052_A net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout408_A _06684_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11004__B2 net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07176_ net1176 team_03_WB.instance_to_wrap.core.register_file.registers_state\[467\]
+ net762 team_03_WB.instance_to_wrap.core.register_file.registers_state\[499\] net1150
+ vssd1 vssd1 vccd1 vccd1 _03118_ sky130_fd_sc_hd__o221a_1
XFILLER_0_14_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07759__A1 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11555__A2 net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout300 _06442_ vssd1 vssd1 vccd1 vccd1 net300 sky130_fd_sc_hd__buf_2
Xfanout311 _05388_ vssd1 vssd1 vccd1 vccd1 net311 sky130_fd_sc_hd__buf_2
XFILLER_0_1_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout777_A _02851_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout398_X net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1309 net1330 vssd1 vssd1 vccd1 vccd1 net1309 sky130_fd_sc_hd__buf_2
Xfanout322 _04833_ vssd1 vssd1 vccd1 vccd1 net322 sky130_fd_sc_hd__clkbuf_2
Xfanout333 _06809_ vssd1 vssd1 vccd1 vccd1 net333 sky130_fd_sc_hd__buf_6
XANTENNA__10515__B1 net1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout344 _06805_ vssd1 vssd1 vccd1 vccd1 net344 sky130_fd_sc_hd__buf_6
XANTENNA_fanout1105_X net1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout355 _06818_ vssd1 vssd1 vccd1 vccd1 net355 sky130_fd_sc_hd__buf_8
Xfanout366 _06815_ vssd1 vssd1 vccd1 vccd1 net366 sky130_fd_sc_hd__clkbuf_4
X_09817_ _02892_ _04679_ net540 vssd1 vssd1 vccd1 vccd1 _05759_ sky130_fd_sc_hd__o21ai_1
Xfanout377 _06812_ vssd1 vssd1 vccd1 vccd1 net377 sky130_fd_sc_hd__clkbuf_8
Xfanout388 _06778_ vssd1 vssd1 vccd1 vccd1 net388 sky130_fd_sc_hd__buf_8
XANTENNA_fanout944_A net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout399 _06752_ vssd1 vssd1 vccd1 vccd1 net399 sky130_fd_sc_hd__buf_4
XANTENNA__11109__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09748_ _02891_ _05689_ vssd1 vssd1 vccd1 vccd1 _05690_ sky130_fd_sc_hd__or2_1
XFILLER_0_97_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09679_ _05568_ _05514_ net320 _05565_ vssd1 vssd1 vccd1 vccd1 _05621_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA_fanout732_X net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_139_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11055__D net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_95_wb_clk_i clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_95_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_11710_ _06459_ _06803_ vssd1 vssd1 vccd1 vccd1 _06808_ sky130_fd_sc_hd__or2_4
XANTENNA__15105__A net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12690_ net1396 vssd1 vssd1 vccd1 vccd1 _00454_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07695__B1 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07790__S0 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_24_wb_clk_i clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_24_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__14717__Q team_03_WB.instance_to_wrap.core.decoder.inst\[14\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11641_ _06715_ net383 net348 net2276 vssd1 vssd1 vccd1 vccd1 _01891_ sky130_fd_sc_hd__a22o_1
XFILLER_0_77_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12035__A3 net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09597__X _05539_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14360_ clknet_leaf_186_wb_clk_i _02124_ _00725_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[714\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_42_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11572_ net642 net708 net266 net700 vssd1 vssd1 vccd1 vccd1 _06799_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_42_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13311_ net1335 vssd1 vssd1 vccd1 vccd1 _01075_ sky130_fd_sc_hd__inv_2
XANTENNA__11779__S net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput19 DAT_I[25] vssd1 vssd1 vccd1 vccd1 net19 sky130_fd_sc_hd__buf_1
X_10523_ net143 net1034 net1026 net1684 vssd1 vssd1 vccd1 vccd1 _02587_ sky130_fd_sc_hd__a22o_1
XFILLER_0_107_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14291_ clknet_leaf_97_wb_clk_i _02055_ _00656_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[645\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_94_2302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_162_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_94_2313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13242_ net1377 vssd1 vssd1 vccd1 vccd1 _01006_ sky130_fd_sc_hd__inv_2
X_10454_ net285 _06054_ _06269_ _06268_ vssd1 vssd1 vccd1 vccd1 _06270_ sky130_fd_sc_hd__a31o_1
XANTENNA__09739__A2 _04953_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input73_A wbs_adr_i[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_131_3063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_1027 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08947__B1 net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11546__A2 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_3074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_423 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13173_ net1276 vssd1 vssd1 vccd1 vccd1 _00937_ sky130_fd_sc_hd__inv_2
X_10385_ _06211_ _06213_ net282 vssd1 vssd1 vccd1 vccd1 _06214_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10754__B1 net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07845__S1 net1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_107_Left_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09773__A net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12124_ net1529 vssd1 vssd1 vccd1 vccd1 _02429_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_182 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13295__A net1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12055_ _06479_ net2702 net355 vssd1 vssd1 vccd1 vccd1 _01491_ sky130_fd_sc_hd__mux2_1
XANTENNA__10506__B1 net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09923__D _05429_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07293__A net1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11006_ net649 _06575_ vssd1 vssd1 vccd1 vccd1 _06576_ sky130_fd_sc_hd__and2_1
XANTENNA__07724__C net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07922__A1 net1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07383__C1 net1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09124__B1 net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09675__A1 _03391_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12957_ net1389 vssd1 vssd1 vccd1 vccd1 _00721_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_66_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09675__B2 net1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06908__Y _02850_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_116_Left_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_29_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_104_wb_clk_i_A clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__07740__B _03681_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07686__B1 net1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11908_ net1043 net656 _06463_ net473 vssd1 vssd1 vccd1 vccd1 _06814_ sky130_fd_sc_hd__or4b_4
XTAP_TAPCELL_ROW_138_3206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08328__S net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11482__B2 net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_478 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_3217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12888_ net1376 vssd1 vssd1 vccd1 vccd1 _00652_ sky130_fd_sc_hd__inv_2
XFILLER_0_158_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_103_2486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14627_ clknet_leaf_47_wb_clk_i _02391_ _00992_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[981\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_8_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_103_2497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10159__A _05041_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_406 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11839_ net654 _06677_ net467 net325 net1851 vssd1 vssd1 vccd1 vccd1 _01700_ sky130_fd_sc_hd__a32o_1
XFILLER_0_157_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_155_3553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07438__B1 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_155_3564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14558_ clknet_leaf_116_wb_clk_i _02322_ _00923_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[912\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13509_ net1317 vssd1 vssd1 vccd1 vccd1 _01273_ sky130_fd_sc_hd__inv_2
XFILLER_0_114_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14489_ clknet_leaf_176_wb_clk_i _02253_ _00854_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[843\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_99_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07030_ _02963_ _02966_ _02971_ net1118 net1139 vssd1 vssd1 vccd1 vccd1 _02972_ sky130_fd_sc_hd__o221a_1
XFILLER_0_141_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11537__A2 net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09060__C1 net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07610__B1 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08981_ net435 net428 _04922_ net551 vssd1 vssd1 vccd1 vccd1 _04923_ sky130_fd_sc_hd__o31a_1
X_07932_ net1181 team_03_WB.instance_to_wrap.core.register_file.registers_state\[215\]
+ vssd1 vssd1 vccd1 vccd1 _03874_ sky130_fd_sc_hd__or2_1
XANTENNA__08166__A1 net1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_143_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_07863_ net808 _03793_ _03794_ vssd1 vssd1 vccd1 vccd1 _03805_ sky130_fd_sc_hd__or3_1
XFILLER_0_78_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09602_ _05171_ _05172_ _05174_ _05338_ vssd1 vssd1 vccd1 vccd1 _05544_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_74_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_2976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07794_ net1097 team_03_WB.instance_to_wrap.core.register_file.registers_state\[715\]
+ net797 team_03_WB.instance_to_wrap.core.register_file.registers_state\[747\] net730
+ vssd1 vssd1 vccd1 vccd1 _03736_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_127_2987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09115__B1 net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09533_ _03566_ _04354_ net535 _05474_ _03564_ vssd1 vssd1 vccd1 vccd1 _05475_ sky130_fd_sc_hd__o311a_1
XANTENNA__07931__A net1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09666__B2 net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout358_A _06818_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_979 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09464_ net547 _04384_ _05096_ vssd1 vssd1 vccd1 vccd1 _05406_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07141__A2 net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08415_ net1228 team_03_WB.instance_to_wrap.core.register_file.registers_state\[186\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[154\] net954 net917
+ vssd1 vssd1 vccd1 vccd1 _04357_ sky130_fd_sc_hd__a221o_1
XFILLER_0_171_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09395_ _05174_ _05336_ vssd1 vssd1 vccd1 vccd1 _05337_ sky130_fd_sc_hd__and2_1
XFILLER_0_80_60 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout525_A _06322_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1267_A net1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09858__A _05768_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07429__B1 net1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08346_ net1235 team_03_WB.instance_to_wrap.core.register_file.registers_state\[341\]
+ net968 team_03_WB.instance_to_wrap.core.register_file.registers_state\[373\] net1072
+ vssd1 vssd1 vccd1 vccd1 _04288_ sky130_fd_sc_hd__o221a_1
XANTENNA__11225__B2 net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_151_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11599__S net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08277_ net1234 team_03_WB.instance_to_wrap.core.register_file.registers_state\[471\]
+ net963 team_03_WB.instance_to_wrap.core.register_file.registers_state\[503\] net1212
+ vssd1 vssd1 vccd1 vccd1 _04219_ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout313_X net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1434_A net1435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1055_X net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07228_ _03139_ _03169_ net613 vssd1 vssd1 vccd1 vccd1 _03170_ sky130_fd_sc_hd__mux2_2
XFILLER_0_85_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_171_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout894_A net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_767 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11528__A2 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08929__B1 net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_142_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_142_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_42_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10008__S net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07159_ net823 _03096_ _03098_ _03100_ net724 vssd1 vssd1 vccd1 vccd1 _03101_ sky130_fd_sc_hd__a41o_1
XANTENNA_clkbuf_leaf_182_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout1222_X net1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09051__C1 net1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10170_ _03758_ _06010_ _06011_ vssd1 vssd1 vccd1 vccd1 _06012_ sky130_fd_sc_hd__nand3_2
XANTENNA_fanout682_X net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_160_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1106 net1108 vssd1 vssd1 vccd1 vccd1 net1106 sky130_fd_sc_hd__clkbuf_4
Xfanout1117 _02786_ vssd1 vssd1 vccd1 vccd1 net1117 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08157__A1 net1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1128 net1129 vssd1 vssd1 vccd1 vccd1 net1128 sky130_fd_sc_hd__buf_4
Xfanout1139 net1141 vssd1 vssd1 vccd1 vccd1 net1139 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_121_1099 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11347__B net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08002__A _03943_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout947_X net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07904__A1 net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11700__A2 net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13860_ clknet_leaf_28_wb_clk_i _01624_ _00225_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[214\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_87_2161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09106__B1 net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_2172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12811_ net1282 vssd1 vssd1 vccd1 vccd1 _00575_ sky130_fd_sc_hd__inv_2
XANTENNA__12459__A net1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13791_ clknet_leaf_21_wb_clk_i _01555_ _00156_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[145\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12110__C1 net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11363__A net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07668__B1 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12742_ net1299 vssd1 vssd1 vccd1 vccd1 _00506_ sky130_fd_sc_hd__inv_2
XFILLER_0_96_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_69_Right_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11082__B _06442_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12673_ net1290 vssd1 vssd1 vccd1 vccd1 _00437_ sky130_fd_sc_hd__inv_2
XFILLER_0_60_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08880__A2 _04770_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_539 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11624_ _06698_ net379 net346 net2470 vssd1 vssd1 vccd1 vccd1 _01908_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_61_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14412_ clknet_leaf_19_wb_clk_i _02176_ _00777_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[766\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08617__C1 net1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_133_3103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_3114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11767__A2 net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14343_ clknet_leaf_109_wb_clk_i _02107_ _00708_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[697\]
+ sky130_fd_sc_hd__dfrtp_1
X_11555_ net2444 net482 _06792_ net496 vssd1 vssd1 vccd1 vccd1 _01965_ sky130_fd_sc_hd__a22o_1
XFILLER_0_25_548 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11302__S net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06904__B net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10506_ net103 net1030 net907 net1599 vssd1 vssd1 vccd1 vccd1 _02603_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_150_3450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14274_ clknet_leaf_174_wb_clk_i _02038_ _00639_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[628\]
+ sky130_fd_sc_hd__dfrtp_1
X_11486_ net642 net708 _06557_ net831 vssd1 vssd1 vccd1 vccd1 _06777_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_150_3461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xmax_cap319 _05746_ vssd1 vssd1 vccd1 vccd1 net319 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_100_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13225_ net1255 vssd1 vssd1 vccd1 vccd1 _00989_ sky130_fd_sc_hd__inv_2
X_10437_ _06057_ _06059_ _06255_ vssd1 vssd1 vccd1 vccd1 _06256_ sky130_fd_sc_hd__o21a_1
XFILLER_0_111_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10727__B1 net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_78_Right_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13156_ net1365 vssd1 vssd1 vccd1 vccd1 _00920_ sky130_fd_sc_hd__inv_2
X_10368_ net304 net303 _06198_ _06199_ vssd1 vssd1 vccd1 vccd1 _06200_ sky130_fd_sc_hd__a211o_1
XFILLER_0_27_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12107_ net1142 net1624 _06820_ vssd1 vssd1 vccd1 vccd1 _00002_ sky130_fd_sc_hd__a21o_1
XANTENNA__11538__A net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13087_ net1347 vssd1 vssd1 vccd1 vccd1 _00851_ sky130_fd_sc_hd__inv_2
X_10299_ team_03_WB.instance_to_wrap.core.pc.current_pc\[13\] _06140_ vssd1 vssd1
+ vccd1 vccd1 _06141_ sky130_fd_sc_hd__and2_1
XANTENNA__08148__A1 net1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1028 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08148__B2 net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12038_ _06776_ net470 net361 net2242 vssd1 vssd1 vccd1 vccd1 _01507_ sky130_fd_sc_hd__a22o_1
XANTENNA__11257__B net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09896__A1 net1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07356__C1 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07371__A2 net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_2526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07751__A net1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_2537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_33 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07108__C1 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13989_ clknet_leaf_11_wb_clk_i _01753_ _00354_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[343\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11273__A net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_87_Right_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_157_3604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11455__A1 net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_2873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_122_2884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09949__Y _05879_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_174_3940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_174_3951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08200_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[883\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[851\]
+ net957 vssd1 vssd1 vccd1 vccd1 _04142_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_174_3962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09180_ net552 _04807_ net537 net667 vssd1 vssd1 vccd1 vccd1 _05122_ sky130_fd_sc_hd__o31ai_1
XTAP_TAPCELL_ROW_174_3973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_247 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08131_ _03604_ _03728_ _03866_ _03990_ vssd1 vssd1 vccd1 vccd1 _04073_ sky130_fd_sc_hd__and4b_1
XFILLER_0_172_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08084__B1 net1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_170_3859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_712 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11212__S net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10966__B1 net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08062_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[438\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[406\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[310\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[278\]
+ net767 net1129 vssd1 vssd1 vccd1 vccd1 _04004_ sky130_fd_sc_hd__mux4_1
XFILLER_0_153_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_4_1__f_wb_clk_i clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_1__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_102_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_144_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07013_ net1099 team_03_WB.instance_to_wrap.core.register_file.registers_state\[963\]
+ vssd1 vssd1 vccd1 vccd1 _02955_ sky130_fd_sc_hd__and2_1
XFILLER_0_4_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_96_Right_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09033__C1 net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08387__A1 net1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_242 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08387__B2 net992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07926__A net1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10194__A1 _04565_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11448__A net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12043__S net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08964_ net1067 _04903_ _04904_ vssd1 vssd1 vccd1 vccd1 _04906_ sky130_fd_sc_hd__or3_1
XANTENNA__11167__B net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07915_ _03854_ _03856_ net1115 vssd1 vssd1 vccd1 vccd1 _03857_ sky130_fd_sc_hd__a21o_1
X_08895_ net1239 team_03_WB.instance_to_wrap.core.register_file.registers_state\[172\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[140\] net979 net926
+ vssd1 vssd1 vccd1 vccd1 _04837_ sky130_fd_sc_hd__a221o_1
XANTENNA__10071__B _05914_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout475_A net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10497__A2 net1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07846_ net717 _03787_ _03776_ _03768_ vssd1 vssd1 vccd1 vccd1 _03788_ sky130_fd_sc_hd__a2bb2o_4
XANTENNA__07661__A net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07777_ net748 _03716_ _03717_ _03718_ _03702_ vssd1 vssd1 vccd1 vccd1 _03719_ sky130_fd_sc_hd__o32a_1
XANTENNA_fanout263_X net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout642_A net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1384_A net1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09516_ net557 _05375_ vssd1 vssd1 vccd1 vccd1 _05458_ sky130_fd_sc_hd__and2_1
XANTENNA__08847__C1 net1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07114__A2 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08311__A1 net1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09447_ _05167_ _05339_ vssd1 vssd1 vccd1 vccd1 _05389_ sky130_fd_sc_hd__nand2_1
XFILLER_0_38_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1172_X net1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout907_A _06285_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout528_X net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09378_ _05318_ _05319_ vssd1 vssd1 vccd1 vccd1 _05320_ sky130_fd_sc_hd__nor2_1
XFILLER_0_47_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_163_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_930 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08329_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[757\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[725\]
+ net968 vssd1 vssd1 vccd1 vccd1 _04271_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1437_X net1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11340_ net491 net619 _06722_ net400 net2286 vssd1 vssd1 vccd1 vccd1 _02110_ sky130_fd_sc_hd__a32o_1
XANTENNA__07822__B1 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout897_X net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11271_ net712 net298 net829 vssd1 vssd1 vccd1 vccd1 _06703_ sky130_fd_sc_hd__and3_1
XANTENNA__09024__C1 net1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13010_ net1396 vssd1 vssd1 vccd1 vccd1 _00774_ sky130_fd_sc_hd__inv_2
X_10222_ _06016_ _06063_ vssd1 vssd1 vccd1 vccd1 _06064_ sky130_fd_sc_hd__or2_1
XANTENNA__09575__B1 _05516_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08431__S net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_37_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11382__B1 net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14730__Q team_03_WB.instance_to_wrap.core.decoder.inst\[27\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10153_ _03985_ _05993_ vssd1 vssd1 vccd1 vccd1 _05995_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_89_2201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_2212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input36_A gpio_in[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14961_ clknet_leaf_95_wb_clk_i _02713_ _01326_ vssd1 vssd1 vccd1 vccd1 net213 sky130_fd_sc_hd__dfrtp_1
X_10084_ _05082_ _05142_ vssd1 vssd1 vccd1 vccd1 _05928_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_54_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09878__A1 net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold8 team_03_WB.instance_to_wrap.core.register_file.registers_state\[948\] vssd1
+ vssd1 vccd1 vccd1 net1501 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11792__S net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13912_ clknet_leaf_4_wb_clk_i _01676_ _00277_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[266\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07889__B1 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14892_ clknet_leaf_61_wb_clk_i _02655_ _01257_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.pc.current_pc\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_13843_ clknet_leaf_102_wb_clk_i _01607_ _00208_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[197\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11093__A net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11437__B2 net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11524__C net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13774_ clknet_leaf_124_wb_clk_i _01538_ _00139_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[128\]
+ sky130_fd_sc_hd__dfrtp_1
X_10986_ _06463_ _06562_ vssd1 vssd1 vccd1 vccd1 _06564_ sky130_fd_sc_hd__nand2_2
XFILLER_0_139_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12725_ net1292 vssd1 vssd1 vccd1 vccd1 _00489_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_100_2423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_2434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_152_3501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08606__S net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12656_ net1410 vssd1 vssd1 vccd1 vccd1 _00420_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11607_ _06557_ net2526 net449 vssd1 vssd1 vccd1 vccd1 _01922_ sky130_fd_sc_hd__mux2_1
X_12587_ net1288 vssd1 vssd1 vccd1 vccd1 _00351_ sky130_fd_sc_hd__inv_2
XANTENNA__09802__A1 net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10412__A2 net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14326_ clknet_leaf_153_wb_clk_i _02090_ _00691_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[680\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07813__B1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11538_ net649 _06648_ vssd1 vssd1 vccd1 vccd1 _06787_ sky130_fd_sc_hd__nor2_1
Xhold408 team_03_WB.instance_to_wrap.BUSY_O vssd1 vssd1 vccd1 vccd1 net1901 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_704 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold419 net231 vssd1 vssd1 vccd1 vccd1 net1912 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_150_350 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09945__B net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14257_ clknet_leaf_139_wb_clk_i _02021_ _00622_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[611\]
+ sky130_fd_sc_hd__dfrtp_1
X_11469_ net2405 net393 _06770_ net505 vssd1 vssd1 vccd1 vccd1 _02029_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_78_1971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_78_1982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08369__A1 net1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13208_ net1380 vssd1 vssd1 vccd1 vccd1 _00972_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_979 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14188_ clknet_leaf_18_wb_clk_i _01952_ _00553_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[542\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13139_ net1265 vssd1 vssd1 vccd1 vccd1 _00903_ sky130_fd_sc_hd__inv_2
XANTENNA__09961__A _03678_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1108 team_03_WB.instance_to_wrap.core.register_file.registers_state\[206\] vssd1
+ vssd1 vccd1 vccd1 net2601 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09869__A1 net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1119 team_03_WB.instance_to_wrap.core.register_file.registers_state\[556\] vssd1
+ vssd1 vccd1 vccd1 net2612 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_174_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07700_ net1101 net899 team_03_WB.instance_to_wrap.core.register_file.registers_state\[13\]
+ vssd1 vssd1 vccd1 vccd1 _03642_ sky130_fd_sc_hd__o21a_1
XFILLER_0_40_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_174_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10479__A2 net1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08680_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[680\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[648\]
+ net975 vssd1 vssd1 vccd1 vccd1 _04622_ sky130_fd_sc_hd__mux2_1
XFILLER_0_174_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_124_2913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_54 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_124_2924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08541__A1 net1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07631_ net1094 team_03_WB.instance_to_wrap.core.register_file.registers_state\[78\]
+ vssd1 vssd1 vccd1 vccd1 _03573_ sky130_fd_sc_hd__and2_1
XFILLER_0_75_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07895__A3 net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11207__S net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11428__A1 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_562 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07562_ net1163 _03503_ vssd1 vssd1 vccd1 vccd1 _03504_ sky130_fd_sc_hd__nor2_1
X_09301_ _03489_ _05242_ vssd1 vssd1 vccd1 vccd1 _05243_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_152_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07493_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[551\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[519\]
+ net785 vssd1 vssd1 vccd1 vccd1 _03435_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_459 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12827__A net1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09232_ _04415_ _05173_ vssd1 vssd1 vccd1 vccd1 _05174_ sky130_fd_sc_hd__or2_2
XFILLER_0_61_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_407 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08516__S net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09201__A net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09163_ _05102_ _05104_ vssd1 vssd1 vccd1 vccd1 _05105_ sky130_fd_sc_hd__nand2_1
XANTENNA__08057__B1 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08114_ net743 _04052_ _04053_ _04054_ _04055_ vssd1 vssd1 vccd1 vccd1 _04056_ sky130_fd_sc_hd__o32a_1
XFILLER_0_161_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_160_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07804__B1 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09094_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[941\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[909\]
+ net977 vssd1 vssd1 vccd1 vccd1 _05036_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10066__B team_03_WB.instance_to_wrap.core.decoder.inst\[30\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08045_ net717 _03962_ _03983_ net617 vssd1 vssd1 vccd1 vccd1 _03987_ sky130_fd_sc_hd__o211a_2
XFILLER_0_141_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09006__C1 net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold920 team_03_WB.instance_to_wrap.core.register_file.registers_state\[517\] vssd1
+ vssd1 vccd1 vccd1 net2413 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_82_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06831__Y _02774_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold931 team_03_WB.instance_to_wrap.core.register_file.registers_state\[797\] vssd1
+ vssd1 vccd1 vccd1 net2424 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1132_A net1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09557__B1 _05498_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold942 team_03_WB.instance_to_wrap.core.register_file.registers_state\[654\] vssd1
+ vssd1 vccd1 vccd1 net2435 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold953 team_03_WB.instance_to_wrap.core.register_file.registers_state\[456\] vssd1
+ vssd1 vccd1 vccd1 net2446 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08251__S net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold964 team_03_WB.instance_to_wrap.core.register_file.registers_state\[649\] vssd1
+ vssd1 vccd1 vccd1 net2457 sky130_fd_sc_hd__dlygate4sd3_1
Xhold975 team_03_WB.instance_to_wrap.core.register_file.registers_state\[137\] vssd1
+ vssd1 vccd1 vccd1 net2468 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11364__B1 net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold986 team_03_WB.instance_to_wrap.core.register_file.registers_state\[844\] vssd1
+ vssd1 vccd1 vccd1 net2479 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11178__A net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold997 team_03_WB.instance_to_wrap.core.register_file.registers_state\[73\] vssd1
+ vssd1 vccd1 vccd1 net2490 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10082__A _05768_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09996_ _05881_ net2073 net287 vssd1 vssd1 vccd1 vccd1 _02718_ sky130_fd_sc_hd__mux2_1
XANTENNA__08780__A1 net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout380_X net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08947_ _04885_ _04886_ net857 vssd1 vssd1 vccd1 vccd1 _04889_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout478_X net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout857_A net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11667__A1 _06519_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08878_ _02944_ _02947_ vssd1 vssd1 vccd1 vccd1 _04820_ sky130_fd_sc_hd__and2b_2
XTAP_TAPCELL_ROW_4_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07829_ net1084 team_03_WB.instance_to_wrap.core.register_file.registers_state\[458\]
+ vssd1 vssd1 vccd1 vccd1 _03771_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout645_X net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11117__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1387_X net1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10840_ net686 _05842_ vssd1 vssd1 vccd1 vccd1 _06441_ sky130_fd_sc_hd__nand2_1
XANTENNA__10890__A2 _05646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_2017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_2028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09924__D_N _05429_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10771_ team_03_WB.instance_to_wrap.core.decoder.inst\[11\] net1018 vssd1 vssd1 vccd1
+ vccd1 _06381_ sky130_fd_sc_hd__nand2_1
XFILLER_0_6_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout812_X net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12737__A net1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12510_ net1385 vssd1 vssd1 vccd1 vccd1 _00274_ sky130_fd_sc_hd__inv_2
X_13490_ net1327 vssd1 vssd1 vccd1 vccd1 _01254_ sky130_fd_sc_hd__inv_2
XANTENNA__08426__S net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_930 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09111__A net1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12441_ net1357 vssd1 vssd1 vccd1 vccd1 _00205_ sky130_fd_sc_hd__inv_2
XFILLER_0_164_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_615 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12372_ net1304 vssd1 vssd1 vccd1 vccd1 _00136_ sky130_fd_sc_hd__inv_2
XFILLER_0_34_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08950__A net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11323_ _06519_ net2067 net406 vssd1 vssd1 vccd1 vccd1 _02122_ sky130_fd_sc_hd__mux2_1
X_14111_ clknet_leaf_170_wb_clk_i _01875_ _00476_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[465\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11787__S net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15091_ net1477 vssd1 vssd1 vccd1 vccd1 la_data_out[27] sky130_fd_sc_hd__buf_2
XFILLER_0_133_884 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07271__A1 net1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12472__A net1380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09548__B1 net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1083 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14042_ clknet_leaf_145_wb_clk_i _01806_ _00407_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[396\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_56_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11254_ net501 net630 _06694_ net409 net2083 vssd1 vssd1 vccd1 vccd1 _02168_ sky130_fd_sc_hd__a32o_1
XANTENNA__08161__S net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10205_ _05953_ _05956_ _05952_ vssd1 vssd1 vccd1 vccd1 _06047_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_128_3002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11088__A net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_3013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11185_ net2272 net414 _06673_ net509 vssd1 vssd1 vccd1 vccd1 _02216_ sky130_fd_sc_hd__a22o_1
XFILLER_0_66_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10136_ _04267_ _02771_ net673 vssd1 vssd1 vccd1 vccd1 _05978_ sky130_fd_sc_hd__mux2_1
XANTENNA__09781__A _02992_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_145_3360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10067_ net1207 net1212 net1219 net1048 vssd1 vssd1 vccd1 vccd1 _05911_ sky130_fd_sc_hd__or4_1
X_14944_ clknet_leaf_43_wb_clk_i _02699_ _01309_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_O\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11658__A1 _06479_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08523__A1 net1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_167_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_159_203 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14875_ clknet_leaf_96_wb_clk_i _02638_ _01240_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.pc.current_pc\[4\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_141_3268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_141_3279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkload1_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13826_ clknet_leaf_172_wb_clk_i _01590_ _00191_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[180\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13757_ clknet_leaf_25_wb_clk_i _01521_ _00122_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[111\]
+ sky130_fd_sc_hd__dfrtp_1
X_10969_ net693 _05082_ _06399_ vssd1 vssd1 vccd1 vccd1 _06549_ sky130_fd_sc_hd__o21ai_1
XANTENNA__12647__A net1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12708_ net1382 vssd1 vssd1 vccd1 vccd1 _00472_ sky130_fd_sc_hd__inv_2
XANTENNA__08336__S net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13688_ clknet_leaf_4_wb_clk_i _01452_ _00053_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[42\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08563__C _04503_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_475 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12639_ net1350 vssd1 vssd1 vccd1 vccd1 _00403_ sky130_fd_sc_hd__inv_2
XFILLER_0_143_637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11189__A3 _06675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11594__A0 net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10397__B2 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_2772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_2783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold205 team_03_WB.instance_to_wrap.core.register_file.registers_state\[558\] vssd1
+ vssd1 vccd1 vccd1 net1698 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07262__A1 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14309_ clknet_leaf_36_wb_clk_i _02073_ _00674_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[663\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_106_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold216 _02530_ vssd1 vssd1 vccd1 vccd1 net1709 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_895 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold227 team_03_WB.instance_to_wrap.core.register_file.registers_state\[554\] vssd1
+ vssd1 vccd1 vccd1 net1720 sky130_fd_sc_hd__dlygate4sd3_1
Xhold238 net203 vssd1 vssd1 vccd1 vccd1 net1731 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_169_3850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold249 team_03_WB.instance_to_wrap.ADR_I\[18\] vssd1 vssd1 vccd1 vccd1 net1742 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11346__B1 net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07907__C net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07014__A1 net1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09850_ net556 _05133_ vssd1 vssd1 vccd1 vccd1 _05792_ sky130_fd_sc_hd__nor2_1
Xfanout707 net708 vssd1 vssd1 vccd1 vccd1 net707 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11897__A1 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout718 net720 vssd1 vssd1 vccd1 vccd1 net718 sky130_fd_sc_hd__buf_6
Xfanout729 net738 vssd1 vssd1 vccd1 vccd1 net729 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_165_3758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_165_3769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09691__A _05623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08801_ net1239 team_03_WB.instance_to_wrap.core.register_file.registers_state\[129\]
+ net983 team_03_WB.instance_to_wrap.core.register_file.registers_state\[161\] net941
+ vssd1 vssd1 vccd1 vccd1 _04743_ sky130_fd_sc_hd__o221a_1
X_09781_ _02992_ _05722_ vssd1 vssd1 vccd1 vccd1 _05723_ sky130_fd_sc_hd__or2_1
X_06993_ _02792_ _02927_ vssd1 vssd1 vccd1 vccd1 _02935_ sky130_fd_sc_hd__nor2_1
X_08732_ net1222 _04671_ _04673_ net1214 vssd1 vssd1 vccd1 vccd1 _04674_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_1_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09711__B1 _03679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10987__D net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08663_ net1224 _04602_ _04603_ vssd1 vssd1 vccd1 vccd1 _04605_ sky130_fd_sc_hd__and3_1
XFILLER_0_15_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07614_ net1158 _03554_ _03555_ net823 vssd1 vssd1 vccd1 vccd1 _03556_ sky130_fd_sc_hd__o31a_1
X_08594_ _04386_ _04448_ _04534_ _04478_ net559 net564 vssd1 vssd1 vccd1 vccd1 _04536_
+ sky130_fd_sc_hd__mux4_2
XANTENNA__10872__A2 net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07545_ net824 _03486_ net723 vssd1 vssd1 vccd1 vccd1 _03487_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_138_Right_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_810 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout340_A _06806_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1082_A net1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11461__A net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07476_ net1184 team_03_WB.instance_to_wrap.core.register_file.registers_state\[981\]
+ net769 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1013\] net1152
+ vssd1 vssd1 vccd1 vccd1 _03418_ sky130_fd_sc_hd__o221a_1
XANTENNA__11821__A1 net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07003__X _02945_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1082 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09215_ _03904_ _05155_ _02937_ vssd1 vssd1 vccd1 vccd1 _05157_ sky130_fd_sc_hd__o21a_1
XFILLER_0_9_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_146_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_hold1288_A team_03_WB.instance_to_wrap.CPU_DAT_O\[14\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout605_A _06295_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_162_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09146_ net432 net425 _04236_ net541 vssd1 vssd1 vccd1 vccd1 _05088_ sky130_fd_sc_hd__o31a_1
XFILLER_0_16_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_162_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11585__A0 net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1071 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08676__S1 _02788_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07253__A1 net1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09077_ net1240 team_03_WB.instance_to_wrap.core.register_file.registers_state\[205\]
+ net982 team_03_WB.instance_to_wrap.core.register_file.registers_state\[237\] net941
+ vssd1 vssd1 vccd1 vccd1 _05019_ sky130_fd_sc_hd__o221a_1
XFILLER_0_130_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_570 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08450__B1 net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1135_X net1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11400__S net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_49_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_49_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_08028_ net1177 team_03_WB.instance_to_wrap.core.register_file.registers_state\[209\]
+ vssd1 vssd1 vccd1 vccd1 _03970_ sky130_fd_sc_hd__or2_1
XANTENNA__10083__Y _05927_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold750 team_03_WB.instance_to_wrap.core.register_file.registers_state\[830\] vssd1
+ vssd1 vccd1 vccd1 net2243 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout974_A _04086_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout595_X net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold761 team_03_WB.instance_to_wrap.core.register_file.registers_state\[677\] vssd1
+ vssd1 vccd1 vccd1 net2254 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold772 team_03_WB.instance_to_wrap.core.register_file.registers_state\[452\] vssd1
+ vssd1 vccd1 vccd1 net2265 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold783 team_03_WB.instance_to_wrap.core.register_file.registers_state\[481\] vssd1
+ vssd1 vccd1 vccd1 net2276 sky130_fd_sc_hd__dlygate4sd3_1
Xhold794 team_03_WB.instance_to_wrap.core.register_file.registers_state\[181\] vssd1
+ vssd1 vccd1 vccd1 net2287 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1302_X net1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08769__X _04711_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11339__C net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09950__A0 _05879_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10811__Y _06418_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09979_ _03059_ net1692 net291 vssd1 vssd1 vccd1 vccd1 _02734_ sky130_fd_sc_hd__mux2_1
X_15069__1455 vssd1 vssd1 vccd1 vccd1 _15069__1455/HI net1455 sky130_fd_sc_hd__conb_1
XANTENNA__10560__B2 _05870_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_157_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12990_ net1414 vssd1 vssd1 vccd1 vccd1 _00754_ sky130_fd_sc_hd__inv_2
XFILLER_0_157_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09702__B1 _05638_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11355__B net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11941_ net1043 net654 net694 net466 vssd1 vssd1 vccd1 vccd1 _06815_ sky130_fd_sc_hd__or4b_4
XFILLER_0_118_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14660_ clknet_leaf_22_wb_clk_i _02424_ _01025_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1014\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_93_1086 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11872_ _06545_ net2418 net377 vssd1 vssd1 vccd1 vccd1 _01668_ sky130_fd_sc_hd__mux2_1
X_13611_ net1341 vssd1 vssd1 vccd1 vccd1 _01375_ sky130_fd_sc_hd__inv_2
XFILLER_0_157_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10823_ net692 _05479_ vssd1 vssd1 vccd1 vccd1 _06427_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_49_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_105_Right_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14591_ clknet_leaf_167_wb_clk_i _02355_ _00956_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[945\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_156_228 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11371__A net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08364__S0 net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_291 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13542_ net1320 vssd1 vssd1 vccd1 vccd1 _01306_ sky130_fd_sc_hd__inv_2
X_10754_ net525 _06369_ _06370_ net530 net1680 vssd1 vssd1 vccd1 vccd1 _02440_ sky130_fd_sc_hd__a32o_1
XANTENNA__09481__A2 _04503_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_153_924 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10685_ team_03_WB.instance_to_wrap.core.pc.current_pc\[30\] _06318_ vssd1 vssd1
+ vccd1 vccd1 _06326_ sky130_fd_sc_hd__or2_1
X_13473_ net1317 vssd1 vssd1 vccd1 vccd1 _01237_ sky130_fd_sc_hd__inv_2
XANTENNA__07995__S net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12424_ net1291 vssd1 vssd1 vccd1 vccd1 _00188_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_97_2366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_97_2377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11576__A0 net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08036__A3 net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_518 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07244__A1 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12355_ net1371 vssd1 vssd1 vccd1 vccd1 _00119_ sky130_fd_sc_hd__inv_2
XFILLER_0_65_1144 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11310__S net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11306_ _06616_ net2570 net407 vssd1 vssd1 vccd1 vccd1 _02139_ sky130_fd_sc_hd__mux2_1
X_15074_ net1460 vssd1 vssd1 vccd1 vccd1 la_data_out[10] sky130_fd_sc_hd__buf_2
X_12286_ net1385 vssd1 vssd1 vccd1 vccd1 _00050_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_147_3400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11237_ net280 net709 net828 vssd1 vssd1 vccd1 vccd1 _06686_ sky130_fd_sc_hd__and3_1
X_14025_ clknet_leaf_116_wb_clk_i _01789_ _00390_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[379\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_112_2680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11879__A1 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_1827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11249__C net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10000__A0 _05885_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_1838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08744__A1 net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_143_3308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11168_ net635 _06662_ vssd1 vssd1 vccd1 vccd1 _06663_ sky130_fd_sc_hd__nor2_1
XANTENNA__10551__A1 net1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_143_3319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07952__C1 net1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10119_ _04504_ team_03_WB.instance_to_wrap.core.pc.current_pc\[30\] net672 vssd1
+ vssd1 vccd1 vccd1 _05961_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_10_wb_clk_i_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_11099_ net835 net297 vssd1 vssd1 vccd1 vccd1 _06626_ sky130_fd_sc_hd__and2_2
XTAP_TAPCELL_ROW_160_3655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_160_3666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14927_ clknet_leaf_51_wb_clk_i _02682_ _01292_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_O\[14\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__11265__B net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11500__A0 _06454_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11980__S net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14858_ clknet_leaf_59_wb_clk_i _02622_ _01223_ vssd1 vssd1 vccd1 vccd1 net113 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_69_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13809_ clknet_leaf_140_wb_clk_i _01573_ _00174_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[163\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_129_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14789_ clknet_leaf_90_wb_clk_i _02553_ _01154_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_I\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_133_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11281__A net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07330_ net1182 team_03_WB.instance_to_wrap.core.register_file.registers_state\[477\]
+ vssd1 vssd1 vccd1 vccd1 _03272_ sky130_fd_sc_hd__or2_1
XFILLER_0_73_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_119_2812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_2823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07261_ net1164 _03201_ _03202_ _03200_ vssd1 vssd1 vccd1 vccd1 _03203_ sky130_fd_sc_hd__o22a_1
XANTENNA__09957__Y _05883_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_143_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_312 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09000_ net1045 team_03_WB.instance_to_wrap.core.register_file.registers_state\[842\]
+ net995 team_03_WB.instance_to_wrap.core.register_file.registers_state\[874\] net1062
+ vssd1 vssd1 vccd1 vccd1 _04942_ sky130_fd_sc_hd__a221o_1
XFILLER_0_143_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_462 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07192_ _03130_ _03131_ _03132_ _03133_ net811 net726 vssd1 vssd1 vccd1 vccd1 _03134_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_42_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_170_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_143_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11031__A2 net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_167_3809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07786__A2 _03681_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09902_ _05563_ _05824_ _05843_ _05583_ vssd1 vssd1 vccd1 vccd1 _05844_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_1_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout504 net506 vssd1 vssd1 vccd1 vccd1 net504 sky130_fd_sc_hd__buf_2
XANTENNA__12840__A net1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11159__C net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout515 net516 vssd1 vssd1 vccd1 vccd1 net515 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09932__A0 _05870_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout526 _02923_ vssd1 vssd1 vccd1 vccd1 net526 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_6_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09833_ net595 _05771_ _05774_ vssd1 vssd1 vccd1 vccd1 _05775_ sky130_fd_sc_hd__o21ai_1
Xfanout537 _04821_ vssd1 vssd1 vccd1 vccd1 net537 sky130_fd_sc_hd__clkbuf_4
Xfanout548 net549 vssd1 vssd1 vccd1 vccd1 net548 sky130_fd_sc_hd__clkbuf_4
Xfanout559 net560 vssd1 vssd1 vccd1 vccd1 net559 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07943__C1 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout388_A _06778_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12051__S net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09764_ net595 _05698_ _05705_ vssd1 vssd1 vccd1 vccd1 _05706_ sky130_fd_sc_hd__o21a_2
X_06976_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[549\] net788
+ net736 _02917_ vssd1 vssd1 vccd1 vccd1 _02918_ sky130_fd_sc_hd__o211a_1
XANTENNA__11175__B net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_167_wb_clk_i clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_167_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_08715_ net864 _04655_ _04656_ _04654_ vssd1 vssd1 vccd1 vccd1 _04657_ sky130_fd_sc_hd__a31o_1
X_09695_ _05196_ _05635_ _05203_ vssd1 vssd1 vccd1 vccd1 _05637_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout555_A net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_99_wb_clk_i_A clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout1297_A net1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11743__X _06809_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08646_ net1053 team_03_WB.instance_to_wrap.core.register_file.registers_state\[710\]
+ net1006 team_03_WB.instance_to_wrap.core.register_file.registers_state\[742\] net927
+ vssd1 vssd1 vccd1 vccd1 _04588_ sky130_fd_sc_hd__a221o_1
XFILLER_0_96_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_543 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08577_ net1235 team_03_WB.instance_to_wrap.core.register_file.registers_state\[605\]
+ net967 team_03_WB.instance_to_wrap.core.register_file.registers_state\[637\] net922
+ vssd1 vssd1 vccd1 vccd1 _04519_ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout722_A _02863_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout343_X net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1085_X net1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09999__A0 _05884_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07528_ _03465_ _03466_ net747 vssd1 vssd1 vccd1 vccd1 _03470_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_147_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_395 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07459_ net812 _03396_ _03397_ _03400_ vssd1 vssd1 vccd1 vccd1 _03401_ sky130_fd_sc_hd__o22a_1
XFILLER_0_36_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout510_X net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11270__A2 net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_568 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_1008 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10470_ net1142 team_03_WB.instance_to_wrap.BUSY_O vssd1 vssd1 vccd1 vccd1 _06282_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_161_242 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08704__S net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07226__A1 net1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09129_ _05042_ _05070_ vssd1 vssd1 vccd1 vccd1 _05071_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_40_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12140_ net1580 vssd1 vssd1 vccd1 vccd1 _02413_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_103_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_92_2263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_876 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout977_X net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_2274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12071_ _06632_ net2699 net357 vssd1 vssd1 vccd1 vccd1 _01475_ sky130_fd_sc_hd__mux2_1
Xhold580 net218 vssd1 vssd1 vccd1 vccd1 net2073 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12750__A net1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold591 team_03_WB.instance_to_wrap.core.register_file.registers_state\[824\] vssd1
+ vssd1 vccd1 vccd1 net2084 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08187__C1 net1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08726__A1 net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11022_ net707 net272 net830 vssd1 vssd1 vccd1 vccd1 _06585_ sky130_fd_sc_hd__and3_1
XFILLER_0_159_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12973_ net1294 vssd1 vssd1 vccd1 vccd1 _00737_ sky130_fd_sc_hd__inv_2
Xhold1280 team_03_WB.instance_to_wrap.core.register_file.registers_state\[199\] vssd1
+ vssd1 vccd1 vccd1 net2773 sky130_fd_sc_hd__dlygate4sd3_1
X_14712_ clknet_leaf_42_wb_clk_i _02476_ _01077_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.decoder.inst\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_11924_ _06622_ net2512 net370 vssd1 vssd1 vccd1 vccd1 _01618_ sky130_fd_sc_hd__mux2_1
X_14643_ clknet_leaf_100_wb_clk_i _02407_ _01008_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[997\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_47_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11855_ _06468_ net2075 net375 vssd1 vssd1 vccd1 vccd1 _01685_ sky130_fd_sc_hd__mux2_1
XANTENNA__06907__B net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11305__S net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08337__S0 net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10806_ _06410_ _06411_ _06412_ vssd1 vssd1 vccd1 vccd1 _06414_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_99_2406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11532__C net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14574_ clknet_leaf_124_wb_clk_i _02338_ _00939_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[928\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_99_2417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11786_ net2095 _06619_ net328 vssd1 vssd1 vccd1 vccd1 _01752_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_64_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13525_ net1306 vssd1 vssd1 vccd1 vccd1 _01289_ sky130_fd_sc_hd__inv_2
X_10737_ net1852 net529 net524 _06360_ vssd1 vssd1 vccd1 vccd1 _02447_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_24_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_343 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11251__D net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_136_3167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_3178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_968 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13456_ net1343 vssd1 vssd1 vccd1 vccd1 _01220_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10668_ _05541_ _05932_ vssd1 vssd1 vccd1 vccd1 _06310_ sky130_fd_sc_hd__nor2_1
XFILLER_0_70_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06923__A net1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11549__B1 net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14913__Q team_03_WB.instance_to_wrap.CPU_DAT_O\[0\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__07217__A1 net1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12407_ net1385 vssd1 vssd1 vccd1 vccd1 _00171_ sky130_fd_sc_hd__inv_2
XFILLER_0_152_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07738__B _03679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_114_2720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10599_ net1683 team_03_WB.instance_to_wrap.CPU_DAT_O\[30\] net841 vssd1 vssd1 vccd1
+ vccd1 _02529_ sky130_fd_sc_hd__mux2_1
X_13387_ net1420 vssd1 vssd1 vccd1 vccd1 _01151_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_11_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput107 net107 vssd1 vssd1 vccd1 vccd1 ADR_O[13] sky130_fd_sc_hd__clkbuf_4
XANTENNA__09793__X _05735_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08965__A1 net1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput118 net118 vssd1 vssd1 vccd1 vccd1 ADR_O[23] sky130_fd_sc_hd__clkbuf_4
Xoutput129 net129 vssd1 vssd1 vccd1 vccd1 ADR_O[4] sky130_fd_sc_hd__clkbuf_4
X_12338_ net1395 vssd1 vssd1 vccd1 vccd1 _00102_ sky130_fd_sc_hd__inv_2
XFILLER_0_142_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06976__B1 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_2628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11975__S net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_2639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15057_ net1443 vssd1 vssd1 vccd1 vccd1 gpio_out[3] sky130_fd_sc_hd__buf_2
XANTENNA__09953__B net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12269_ net1332 vssd1 vssd1 vccd1 vccd1 _00033_ sky130_fd_sc_hd__inv_2
XANTENNA__08717__A1 net1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14008_ clknet_leaf_186_wb_clk_i _01772_ _00373_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[362\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_162_3706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_133_wb_clk_i_A clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_06830_ team_03_WB.instance_to_wrap.core.pc.current_pc\[14\] vssd1 vssd1 vccd1 vccd1
+ _02773_ sky130_fd_sc_hd__inv_2
X_08500_ net1223 _04440_ _04441_ vssd1 vssd1 vccd1 vccd1 _04442_ sky130_fd_sc_hd__o21ai_1
X_09480_ _02953_ net573 _05421_ vssd1 vssd1 vccd1 vccd1 _05422_ sky130_fd_sc_hd__and3_1
XFILLER_0_77_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12029__A1 net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08431_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[570\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[538\]
+ net964 vssd1 vssd1 vccd1 vccd1 _04373_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11215__S net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08362_ net1236 team_03_WB.instance_to_wrap.core.register_file.registers_state\[342\]
+ net970 team_03_WB.instance_to_wrap.core.register_file.registers_state\[374\] net1072
+ vssd1 vssd1 vccd1 vccd1 _04304_ sky130_fd_sc_hd__o221a_1
XFILLER_0_46_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07313_ net1185 team_03_WB.instance_to_wrap.core.register_file.registers_state\[573\]
+ net879 vssd1 vssd1 vccd1 vccd1 _03255_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_22_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_22_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11252__A2 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08293_ _04223_ _04234_ net850 vssd1 vssd1 vccd1 vccd1 _04235_ sky130_fd_sc_hd__mux2_8
XFILLER_0_128_272 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15068__1454 vssd1 vssd1 vccd1 vccd1 _15068__1454/HI net1454 sky130_fd_sc_hd__conb_1
XANTENNA__07488__X _03430_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07244_ net746 _03183_ _03184_ net1148 vssd1 vssd1 vccd1 vccd1 _03186_ sky130_fd_sc_hd__a31o_1
XFILLER_0_6_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_376 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_144_776 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_927 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11004__A2 net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07175_ net1176 team_03_WB.instance_to_wrap.core.register_file.registers_state\[339\]
+ net762 team_03_WB.instance_to_wrap.core.register_file.registers_state\[371\] net1125
+ vssd1 vssd1 vccd1 vccd1 _03117_ sky130_fd_sc_hd__o221a_1
XFILLER_0_147_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12046__S net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout303_A _05945_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_172_wb_clk_i_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_48_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1045_A net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08956__A1 net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1048 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11960__B1 net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1212_A net1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout301 _06438_ vssd1 vssd1 vccd1 vccd1 net301 sky130_fd_sc_hd__buf_2
Xfanout312 _05388_ vssd1 vssd1 vccd1 vccd1 net312 sky130_fd_sc_hd__buf_2
XANTENNA__07664__A net1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout323 _06811_ vssd1 vssd1 vccd1 vccd1 net323 sky130_fd_sc_hd__clkbuf_8
Xfanout334 _06809_ vssd1 vssd1 vccd1 vccd1 net334 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout293_X net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout672_A net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout345 _06805_ vssd1 vssd1 vccd1 vccd1 net345 sky130_fd_sc_hd__buf_4
XANTENNA__11186__A net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout356 _06818_ vssd1 vssd1 vccd1 vccd1 net356 sky130_fd_sc_hd__buf_4
X_09816_ _05614_ _05615_ _02954_ vssd1 vssd1 vccd1 vccd1 _05758_ sky130_fd_sc_hd__o21ai_1
Xfanout367 _06814_ vssd1 vssd1 vccd1 vccd1 net367 sky130_fd_sc_hd__buf_8
XANTENNA__10090__A _05623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1000_X net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout378 _06812_ vssd1 vssd1 vccd1 vccd1 net378 sky130_fd_sc_hd__clkbuf_4
Xfanout389 _06778_ vssd1 vssd1 vccd1 vccd1 net389 sky130_fd_sc_hd__buf_4
X_09747_ _05613_ _05688_ net575 vssd1 vssd1 vccd1 vccd1 _05689_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout460_X net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06959_ net1112 team_03_WB.instance_to_wrap.core.register_file.registers_state\[325\]
+ net802 team_03_WB.instance_to_wrap.core.register_file.registers_state\[357\] net1158
+ vssd1 vssd1 vccd1 vccd1 _02901_ sky130_fd_sc_hd__a221o_1
XFILLER_0_20_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout558_X net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout937_A net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09678_ _04834_ _05577_ _05617_ _05619_ vssd1 vssd1 vccd1 vccd1 _05620_ sky130_fd_sc_hd__o211a_1
XANTENNA__09684__A2 _04178_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09090__S net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08629_ net1053 team_03_WB.instance_to_wrap.core.register_file.registers_state\[70\]
+ net1007 team_03_WB.instance_to_wrap.core.register_file.registers_state\[102\] net941
+ vssd1 vssd1 vccd1 vccd1 _04571_ sky130_fd_sc_hd__a221o_1
XANTENNA__07695__A1 net1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout725_X net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1029 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11640_ _06714_ net383 net348 net2205 vssd1 vssd1 vccd1 vccd1 _01892_ sky130_fd_sc_hd__a22o_1
XANTENNA__07790__S1 net1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07447__A1 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11571_ net2157 net484 _06798_ net509 vssd1 vssd1 vccd1 vccd1 _01955_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_42_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_64_wb_clk_i clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_64_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__15121__A net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13310_ net1314 vssd1 vssd1 vccd1 vccd1 _01074_ sky130_fd_sc_hd__inv_2
X_10522_ net144 net1034 net1026 net1711 vssd1 vssd1 vccd1 vccd1 _02588_ sky130_fd_sc_hd__a22o_1
XANTENNA__07542__S1 net1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14290_ clknet_leaf_164_wb_clk_i _02054_ _00655_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[644\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08434__S net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_2303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_2314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14733__Q team_03_WB.instance_to_wrap.core.decoder.inst\[30\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10453_ _06037_ _06053_ vssd1 vssd1 vccd1 vccd1 _06269_ sky130_fd_sc_hd__or2_1
X_13241_ net1351 vssd1 vssd1 vccd1 vccd1 _01005_ sky130_fd_sc_hd__inv_2
XFILLER_0_122_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_3064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_3075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_1039 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10384_ _06086_ _06212_ vssd1 vssd1 vccd1 vccd1 _06213_ sky130_fd_sc_hd__nor2_1
X_13172_ net1308 vssd1 vssd1 vccd1 vccd1 _00936_ sky130_fd_sc_hd__inv_2
XANTENNA_input66_A wb_rst_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10754__A1 net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_971 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_435 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1136 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11795__S net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11951__B1 net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12123_ net1608 vssd1 vssd1 vccd1 vccd1 _02430_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__10552__X _06295_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07574__A net1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12054_ _06621_ net2698 net355 vssd1 vssd1 vccd1 vccd1 _01492_ sky130_fd_sc_hd__mux2_1
XANTENNA__10506__A1 net103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11703__B1 net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11005_ net1044 net837 net301 net670 vssd1 vssd1 vccd1 vccd1 _06575_ sky130_fd_sc_hd__and4_1
XFILLER_0_99_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07383__B1 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08580__C1 net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout890 net891 vssd1 vssd1 vccd1 vccd1 net890 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_88_903 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09124__A1 net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10809__A2 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12956_ net1419 vssd1 vssd1 vccd1 vccd1 _00720_ sky130_fd_sc_hd__inv_2
XANTENNA__09675__A2 _04119_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11907_ net645 _06716_ net477 net373 net2144 vssd1 vssd1 vccd1 vccd1 _01634_ sky130_fd_sc_hd__a32o_1
XFILLER_0_158_835 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11482__A2 net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_3207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12887_ net1386 vssd1 vssd1 vccd1 vccd1 _00651_ sky130_fd_sc_hd__inv_2
XFILLER_0_157_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_138_3218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14626_ clknet_leaf_176_wb_clk_i _02390_ _00991_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[980\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_103_2487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11838_ _06676_ net468 net325 net1898 vssd1 vssd1 vccd1 vccd1 _01701_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_103_2498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10159__B net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_570 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07438__A1 net1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_155_3554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_88 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14557_ clknet_leaf_165_wb_clk_i _02321_ _00922_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[911\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_155_3565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11769_ _06602_ net470 net333 net2573 vssd1 vssd1 vccd1 vccd1 _01768_ sky130_fd_sc_hd__a22o_1
XFILLER_0_43_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13508_ net1322 vssd1 vssd1 vccd1 vccd1 _01272_ sky130_fd_sc_hd__inv_2
X_14488_ clknet_leaf_187_wb_clk_i _02252_ _00853_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[842\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10993__B2 net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_0__f_wb_clk_i clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_0__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_153_584 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13439_ net1432 vssd1 vssd1 vccd1 vccd1 _01203_ sky130_fd_sc_hd__inv_2
XANTENNA__10175__A _03789_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_646 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08938__A1 net1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08399__C1 net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11942__B1 net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15109_ net1484 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[14] sky130_fd_sc_hd__buf_2
XANTENNA__07071__C1 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07610__A1 net1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08980_ net853 _04908_ _04921_ vssd1 vssd1 vccd1 vccd1 _04922_ sky130_fd_sc_hd__o21a_4
XFILLER_0_139_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07931_ net1087 team_03_WB.instance_to_wrap.core.register_file.registers_state\[247\]
+ net892 vssd1 vssd1 vccd1 vccd1 _03873_ sky130_fd_sc_hd__or3_1
X_07862_ _03802_ _03803_ net813 vssd1 vssd1 vccd1 vccd1 _03804_ sky130_fd_sc_hd__a21o_1
X_09601_ _05174_ _05338_ _05171_ _05172_ vssd1 vssd1 vccd1 vccd1 _05543_ sky130_fd_sc_hd__a211o_1
XANTENNA__08571__C1 net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_2977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07793_ net1097 team_03_WB.instance_to_wrap.core.register_file.registers_state\[587\]
+ net797 team_03_WB.instance_to_wrap.core.register_file.registers_state\[619\] net746
+ vssd1 vssd1 vccd1 vccd1 _03735_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_127_2988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09115__A1 net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_155_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09532_ _03566_ _04354_ net664 _05473_ vssd1 vssd1 vccd1 vccd1 _05474_ sky130_fd_sc_hd__a22o_1
XANTENNA__07126__B1 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14818__Q net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09204__A net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09463_ _05088_ _05097_ vssd1 vssd1 vccd1 vccd1 _05405_ sky130_fd_sc_hd__nor2_1
XFILLER_0_149_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08414_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[58\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[26\]
+ net954 vssd1 vssd1 vccd1 vccd1 _04356_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09394_ _04415_ _05173_ vssd1 vssd1 vccd1 vccd1 _05336_ sky130_fd_sc_hd__nand2_1
XFILLER_0_19_535 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08345_ net861 _04283_ _04286_ vssd1 vssd1 vccd1 vccd1 _04287_ sky130_fd_sc_hd__o21a_1
XANTENNA__11225__A2 net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1013 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08626__B1 net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09858__B _05784_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout420_A _06560_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1162_A net1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout518_A _06395_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08276_ net1234 team_03_WB.instance_to_wrap.core.register_file.registers_state\[343\]
+ net963 team_03_WB.instance_to_wrap.core.register_file.registers_state\[375\] net1072
+ vssd1 vssd1 vccd1 vccd1 _04218_ sky130_fd_sc_hd__o221a_1
XFILLER_0_61_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07227_ net721 _03152_ _03168_ vssd1 vssd1 vccd1 vccd1 _03169_ sky130_fd_sc_hd__o21a_4
XANTENNA_fanout306_X net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1048_X net1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07158_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[256\] net785
+ _03099_ vssd1 vssd1 vccd1 vccd1 _03100_ sky130_fd_sc_hd__a21o_1
XANTENNA__09051__B1 net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10736__A1 _05659_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07089_ net1102 team_03_WB.instance_to_wrap.core.register_file.registers_state\[577\]
+ vssd1 vssd1 vccd1 vccd1 _03031_ sky130_fd_sc_hd__and2_1
XFILLER_0_160_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1215_X net1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09085__S net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_182_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_182_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xfanout1107 net1108 vssd1 vssd1 vccd1 vccd1 net1107 sky130_fd_sc_hd__clkbuf_2
Xfanout1118 net1119 vssd1 vssd1 vccd1 vccd1 net1118 sky130_fd_sc_hd__buf_4
XANTENNA_fanout675_X net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1129 net1130 vssd1 vssd1 vccd1 vccd1 net1129 sky130_fd_sc_hd__buf_2
Xclkbuf_leaf_111_wb_clk_i clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_111_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__11347__C net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11161__B2 net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout842_X net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_2162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09106__A1 net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12810_ net1279 vssd1 vssd1 vccd1 vccd1 _00574_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_87_2173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13790_ clknet_leaf_118_wb_clk_i _01554_ _00155_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[144\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08314__C1 net1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14728__Q team_03_WB.instance_to_wrap.core.decoder.inst\[25\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12741_ net1354 vssd1 vssd1 vccd1 vccd1 _00505_ sky130_fd_sc_hd__inv_2
XANTENNA__07668__A1 net1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11363__B net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12672_ net1402 vssd1 vssd1 vccd1 vccd1 _00436_ sky130_fd_sc_hd__inv_2
XFILLER_0_155_827 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08880__A3 net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14411_ clknet_leaf_41_wb_clk_i _02175_ _00776_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[765\]
+ sky130_fd_sc_hd__dfrtp_1
X_11623_ _06697_ net380 net346 net2281 vssd1 vssd1 vccd1 vccd1 _01909_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_61_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08617__B1 net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_154_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_3104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_133_3115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14342_ clknet_leaf_73_wb_clk_i _02106_ _00707_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[696\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_242 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08164__S net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11554_ net648 _06664_ vssd1 vssd1 vccd1 vccd1 _06792_ sky130_fd_sc_hd__nor2_1
X_10505_ net114 net1033 net908 net1552 vssd1 vssd1 vccd1 vccd1 _02604_ sky130_fd_sc_hd__a22o_1
X_14273_ clknet_leaf_180_wb_clk_i _02037_ _00638_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[627\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_150_3451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_746 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11485_ net2406 net393 _06776_ net509 vssd1 vssd1 vccd1 vccd1 _02019_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_150_3462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire587 _05883_ vssd1 vssd1 vccd1 vccd1 net587 sky130_fd_sc_hd__buf_2
XFILLER_0_150_543 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13224_ net1298 vssd1 vssd1 vccd1 vccd1 _00988_ sky130_fd_sc_hd__inv_2
X_10436_ _05925_ _05945_ _06060_ vssd1 vssd1 vccd1 vccd1 _06255_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_61_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input69_X net69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13155_ net1354 vssd1 vssd1 vccd1 vccd1 _00919_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_59_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10367_ _05981_ _06089_ _06094_ vssd1 vssd1 vccd1 vccd1 _06199_ sky130_fd_sc_hd__and3_1
X_12106_ net1143 net1145 _06293_ vssd1 vssd1 vccd1 vccd1 _06820_ sky130_fd_sc_hd__and3_1
X_10298_ team_03_WB.instance_to_wrap.core.pc.current_pc\[12\] team_03_WB.instance_to_wrap.core.pc.current_pc\[11\]
+ _06139_ vssd1 vssd1 vccd1 vccd1 _06140_ sky130_fd_sc_hd__and3_1
X_13086_ net1414 vssd1 vssd1 vccd1 vccd1 _00850_ sky130_fd_sc_hd__inv_2
X_12037_ net634 _06606_ net467 net361 net2094 vssd1 vssd1 vccd1 vccd1 _01508_ sky130_fd_sc_hd__a32o_1
XFILLER_0_109_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11257__C net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07356__B1 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09896__A2 _02804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15067__1453 vssd1 vssd1 vccd1 vccd1 _15067__1453/HI net1453 sky130_fd_sc_hd__conb_1
XANTENNA__11554__A net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_2527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08339__S net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07108__B1 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13988_ clknet_leaf_30_wb_clk_i _01752_ _00353_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[342\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_149_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12101__B1 net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08305__C1 net1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07659__A1 team_03_WB.instance_to_wrap.core.decoder.inst\[14\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11273__B net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07470__C net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11455__A2 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12939_ net1283 vssd1 vssd1 vccd1 vccd1 _00703_ sky130_fd_sc_hd__inv_2
XFILLER_0_158_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_157_3605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10112__C1 _03065_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_2874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_122_2885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09959__A _03600_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_174_3941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_174_3952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14609_ clknet_leaf_139_wb_clk_i _02373_ _00974_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[963\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_174_3963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08608__B1 _04097_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_174_3974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_151 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08130_ _03604_ _03728_ vssd1 vssd1 vccd1 vccd1 _04072_ sky130_fd_sc_hd__and2b_1
XFILLER_0_7_259 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10966__A1 net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_724 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08061_ net1090 team_03_WB.instance_to_wrap.core.register_file.registers_state\[502\]
+ net895 _04002_ net1153 vssd1 vssd1 vccd1 vccd1 _04003_ sky130_fd_sc_hd__o311a_1
XFILLER_0_109_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07292__C1 net1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07831__B2 net1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07012_ net584 _02953_ vssd1 vssd1 vccd1 vccd1 _02954_ sky130_fd_sc_hd__and2_4
XFILLER_0_71_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09033__B1 net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11915__A0 _06616_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_1153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08963_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[425\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[393\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[297\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[265\]
+ net986 net1079 vssd1 vssd1 vccd1 vccd1 _04905_ sky130_fd_sc_hd__mux4_1
XANTENNA__11448__B net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08103__A net1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07914_ net1178 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1007\]
+ net878 _03855_ net1126 vssd1 vssd1 vccd1 vccd1 _03856_ sky130_fd_sc_hd__a311o_1
X_08894_ net926 _04835_ vssd1 vssd1 vccd1 vccd1 _04836_ sky130_fd_sc_hd__nand2_1
XANTENNA__07347__B1 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09887__A2 _04148_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1008_A _04085_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07845_ _03779_ _03780_ _03785_ _03786_ net1114 net1138 vssd1 vssd1 vccd1 vccd1 _03787_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__11694__A2 net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout370_A _06814_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout468_A net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11464__A net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_1141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07661__B _03601_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07776_ net1194 team_03_WB.instance_to_wrap.core.register_file.registers_state\[684\]
+ net897 net1133 vssd1 vssd1 vccd1 vccd1 _03718_ sky130_fd_sc_hd__a211o_1
XFILLER_0_78_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09515_ _05325_ _05327_ _05430_ vssd1 vssd1 vccd1 vccd1 _05457_ sky130_fd_sc_hd__nor3_1
XFILLER_0_149_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_917 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08847__B1 net1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout635_A net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_643 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1377_A net1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09446_ _05346_ _05347_ _05386_ vssd1 vssd1 vccd1 vccd1 _05388_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_82_2070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_149_676 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_490 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09377_ _04445_ _05317_ vssd1 vssd1 vccd1 vccd1 _05319_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout423_X net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout802_A net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11403__S net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1165_X net1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08328_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[693\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[661\]
+ net969 vssd1 vssd1 vccd1 vccd1 _04270_ sky130_fd_sc_hd__mux2_1
XANTENNA__11749__A3 net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15112__1485 vssd1 vssd1 vccd1 vccd1 _15112__1485/HI net1485 sky130_fd_sc_hd__conb_1
XFILLER_0_163_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09272__B1 net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08075__B2 net1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_942 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10957__A1 team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[3\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_771 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08259_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[882\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[850\]
+ net951 vssd1 vssd1 vccd1 vccd1 _04201_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11270_ net504 net634 _06702_ net410 net1974 vssd1 vssd1 vccd1 vccd1 _02160_ sky130_fd_sc_hd__a32o_1
XANTENNA__09024__B1 net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout792_X net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11906__B1 net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09575__A1 net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10221_ _06017_ _06021_ _06062_ vssd1 vssd1 vccd1 vccd1 _06063_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_37_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11382__A1 net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10152_ _03985_ _05993_ vssd1 vssd1 vccd1 vccd1 _05994_ sky130_fd_sc_hd__or2_1
XANTENNA__07050__A2 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_2202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_2213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14960_ clknet_leaf_96_wb_clk_i _02712_ _01325_ vssd1 vssd1 vccd1 vccd1 net212 sky130_fd_sc_hd__dfrtp_1
X_10083_ _02954_ _05107_ _05141_ _05082_ vssd1 vssd1 vccd1 vccd1 _05927_ sky130_fd_sc_hd__a211oi_2
XTAP_TAPCELL_ROW_54_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07338__A0 _03277_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold9 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1014\] vssd1
+ vssd1 vccd1 vccd1 net1502 sky130_fd_sc_hd__dlygate4sd3_1
X_13911_ clknet_leaf_76_wb_clk_i _01675_ _00276_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[265\]
+ sky130_fd_sc_hd__dfrtp_1
X_14891_ clknet_leaf_61_wb_clk_i _02654_ _01256_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.pc.current_pc\[20\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__11685__A2 net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input29_A DAT_I[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13842_ clknet_leaf_164_wb_clk_i _01606_ _00207_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[196\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07063__S net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11093__B net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11437__A2 net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13773_ clknet_leaf_188_wb_clk_i _01537_ _00138_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[127\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_168_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10985_ _06462_ net696 vssd1 vssd1 vccd1 vccd1 _06563_ sky130_fd_sc_hd__nor2_2
XANTENNA__11524__D net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10645__A0 net1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07105__A3 net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12724_ net1304 vssd1 vssd1 vccd1 vccd1 _00488_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_100_2424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_2435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09131__X _05073_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12655_ net1337 vssd1 vssd1 vccd1 vccd1 _00419_ sky130_fd_sc_hd__inv_2
XFILLER_0_154_123 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_152_3502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11313__S net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11606_ _06550_ net2666 net449 vssd1 vssd1 vccd1 vccd1 _01923_ sky130_fd_sc_hd__mux2_1
X_12586_ net1285 vssd1 vssd1 vccd1 vccd1 _00350_ sky130_fd_sc_hd__inv_2
XFILLER_0_81_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_964 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14325_ clknet_leaf_107_wb_clk_i _02089_ _00690_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[679\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_111_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07813__A1 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11537_ net1945 net483 _06786_ net497 vssd1 vssd1 vccd1 vccd1 _01977_ sky130_fd_sc_hd__a22o_1
XFILLER_0_151_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_154 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_463 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold409 net116 vssd1 vssd1 vccd1 vccd1 net1902 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07586__X _03528_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14256_ clknet_leaf_156_wb_clk_i _02020_ _00621_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[610\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_111_716 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08622__S net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11468_ net653 _06593_ vssd1 vssd1 vccd1 vccd1 _06770_ sky130_fd_sc_hd__nor2_1
XFILLER_0_150_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_587 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_1983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09566__A1 net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14921__Q team_03_WB.instance_to_wrap.CPU_DAT_O\[8\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09110__S0 net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13207_ net1391 vssd1 vssd1 vccd1 vccd1 _00971_ sky130_fd_sc_hd__inv_2
XFILLER_0_96_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10419_ _06240_ _06241_ team_03_WB.instance_to_wrap.core.pc.current_pc\[12\] net680
+ vssd1 vssd1 vccd1 vccd1 _02646_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_21_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14187_ clknet_leaf_46_wb_clk_i _01951_ _00552_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[541\]
+ sky130_fd_sc_hd__dfrtp_1
X_11399_ net281 net2565 net396 vssd1 vssd1 vccd1 vccd1 _02081_ sky130_fd_sc_hd__mux2_1
XANTENNA__08774__C1 net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13138_ net1397 vssd1 vssd1 vccd1 vccd1 _00902_ sky130_fd_sc_hd__inv_2
XANTENNA__11983__S net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13069_ net1331 vssd1 vssd1 vccd1 vccd1 _00833_ sky130_fd_sc_hd__inv_2
XANTENNA__09961__B net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_max_cap319_X net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1109 team_03_WB.instance_to_wrap.core.register_file.registers_state\[323\] vssd1
+ vssd1 vccd1 vccd1 net2602 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11125__B2 net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07762__A net1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_119_Right_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10599__S net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_2914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_124_2925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_66 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07630_ net730 _03568_ _03569_ _03570_ _03571_ vssd1 vssd1 vccd1 vccd1 _03572_ sky130_fd_sc_hd__a32o_1
XANTENNA__10884__B1 net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11428__A2 net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07561_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[440\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[408\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[312\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[280\]
+ net772 net1130 vssd1 vssd1 vccd1 vccd1 _03503_ sky130_fd_sc_hd__mux4_1
XFILLER_0_88_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10636__A0 team_03_WB.instance_to_wrap.core.decoder.inst\[25\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09300_ net526 _05144_ net609 vssd1 vssd1 vccd1 vccd1 _05242_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_76_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_158_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07492_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[935\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[903\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[807\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[775\]
+ net785 net1135 vssd1 vssd1 vccd1 vccd1 _03434_ sky130_fd_sc_hd__mux4_1
XANTENNA__07501__B1 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09231_ _03314_ _05161_ vssd1 vssd1 vccd1 vccd1 _05173_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_111_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11223__S net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_wire593_X net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09162_ net547 _04417_ _05103_ net559 vssd1 vssd1 vccd1 vccd1 _05104_ sky130_fd_sc_hd__a211o_1
XFILLER_0_174_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_871 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08113_ net1088 team_03_WB.instance_to_wrap.core.register_file.registers_state\[666\]
+ net892 net1124 vssd1 vssd1 vccd1 vccd1 _04055_ sky130_fd_sc_hd__a211o_1
XFILLER_0_114_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07804__A1 net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09093_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[813\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[781\]
+ net983 vssd1 vssd1 vccd1 vccd1 _05035_ sky130_fd_sc_hd__mux2_1
XANTENNA__12843__A net1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10066__C _02872_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08044_ net613 _03985_ vssd1 vssd1 vccd1 vccd1 _03986_ sky130_fd_sc_hd__nor2_1
XANTENNA__08532__S net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_251 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold910 team_03_WB.instance_to_wrap.core.register_file.registers_state\[521\] vssd1
+ vssd1 vccd1 vccd1 net2403 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06841__A net1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold921 team_03_WB.instance_to_wrap.core.register_file.registers_state\[792\] vssd1
+ vssd1 vccd1 vccd1 net2414 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09557__A1 net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold932 team_03_WB.instance_to_wrap.core.register_file.registers_state\[794\] vssd1
+ vssd1 vccd1 vccd1 net2425 sky130_fd_sc_hd__dlygate4sd3_1
Xhold943 team_03_WB.instance_to_wrap.core.register_file.registers_state\[725\] vssd1
+ vssd1 vccd1 vccd1 net2436 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12054__S net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold954 team_03_WB.instance_to_wrap.core.register_file.registers_state\[333\] vssd1
+ vssd1 vccd1 vccd1 net2447 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1125_A net1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold965 team_03_WB.instance_to_wrap.core.register_file.registers_state\[542\] vssd1
+ vssd1 vccd1 vccd1 net2458 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11364__A1 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07568__B1 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold976 team_03_WB.instance_to_wrap.core.register_file.registers_state\[351\] vssd1
+ vssd1 vccd1 vccd1 net2469 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08765__C1 net1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold987 team_03_WB.instance_to_wrap.core.register_file.registers_state\[881\] vssd1
+ vssd1 vccd1 vccd1 net2480 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11903__A3 net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold998 net209 vssd1 vssd1 vccd1 vccd1 net2491 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11178__B _06517_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09995_ _05880_ net1781 net289 vssd1 vssd1 vccd1 vccd1 _02719_ sky130_fd_sc_hd__mux2_1
XANTENNA__10082__B _05784_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout585_A net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_134_Left_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08946_ net1060 team_03_WB.instance_to_wrap.core.register_file.registers_state\[683\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[651\] net997 net940
+ vssd1 vssd1 vccd1 vccd1 _04888_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_32_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08877_ net556 _04770_ _04817_ net667 vssd1 vssd1 vccd1 vccd1 _04819_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_4_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout373_X net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout752_A net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11194__A net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10875__B1 net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07828_ net1082 team_03_WB.instance_to_wrap.core.register_file.registers_state\[330\]
+ net1149 vssd1 vssd1 vccd1 vccd1 _03770_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_84_2110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_169_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout540_X net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07759_ net819 _03692_ net723 vssd1 vssd1 vccd1 vccd1 _03701_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout1282_X net1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout638_X net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_2018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_80_2029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10770_ team_03_WB.instance_to_wrap.core.decoder.inst\[10\] net1018 vssd1 vssd1 vccd1
+ vccd1 _06380_ sky130_fd_sc_hd__nand2_1
XFILLER_0_17_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12092__A2 net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_143_Left_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09429_ net583 _04830_ vssd1 vssd1 vccd1 vccd1 _05371_ sky130_fd_sc_hd__nor2_4
XFILLER_0_164_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout805_X net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12440_ net1379 vssd1 vssd1 vccd1 vccd1 _00204_ sky130_fd_sc_hd__inv_2
XFILLER_0_81_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08048__B2 _03987_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08008__A net1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_627 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11052__B1 net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12371_ net1255 vssd1 vssd1 vccd1 vccd1 _00135_ sky130_fd_sc_hd__inv_2
X_15066__1452 vssd1 vssd1 vccd1 vccd1 _15066__1452/HI net1452 sky130_fd_sc_hd__conb_1
XANTENNA__10825__X _06429_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12753__A net1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14110_ clknet_leaf_120_wb_clk_i _01874_ _00475_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[464\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07847__A team_03_WB.instance_to_wrap.core.decoder.inst\[30\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11322_ _06628_ net2471 net407 vssd1 vssd1 vccd1 vccd1 _02123_ sky130_fd_sc_hd__mux2_1
X_15090_ net1476 vssd1 vssd1 vccd1 vccd1 la_data_out[26] sky130_fd_sc_hd__buf_2
XFILLER_0_127_1040 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11369__A net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14041_ clknet_leaf_169_wb_clk_i _01805_ _00406_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[395\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_56_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11253_ _06442_ net711 net828 vssd1 vssd1 vccd1 vccd1 _06694_ sky130_fd_sc_hd__and3_1
XFILLER_0_127_1095 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07559__B1 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_152_Left_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08756__C1 net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07058__S net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10204_ net592 _05950_ _06045_ _02994_ vssd1 vssd1 vccd1 vccd1 _06046_ sky130_fd_sc_hd__a211oi_1
XTAP_TAPCELL_ROW_128_3003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08220__A1 net1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_3014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11184_ net659 net705 _06527_ net697 vssd1 vssd1 vccd1 vccd1 _06673_ sky130_fd_sc_hd__and4_1
XFILLER_0_66_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_73_1880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10135_ _05976_ vssd1 vssd1 vccd1 vccd1 _05977_ sky130_fd_sc_hd__inv_2
XANTENNA__08678__A _04619_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_3350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08508__C1 net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_3361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14943_ clknet_leaf_51_wb_clk_i _02698_ _01308_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_O\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_10066_ team_03_WB.instance_to_wrap.core.decoder.inst\[31\] team_03_WB.instance_to_wrap.core.decoder.inst\[30\]
+ _02872_ _05909_ vssd1 vssd1 vccd1 vccd1 _05910_ sky130_fd_sc_hd__or4_1
XANTENNA__11308__S net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10866__B1 net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14874_ clknet_leaf_93_wb_clk_i _02637_ _01239_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.pc.current_pc\[3\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_82_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_141_3269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07731__B1 net1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13825_ clknet_leaf_183_wb_clk_i _01589_ _00190_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[179\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_173_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12928__A net1402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_161_Left_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13756_ clknet_leaf_148_wb_clk_i _01520_ _00121_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[110\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10968_ team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[1\] net308 net688 vssd1
+ vssd1 vccd1 vccd1 _06548_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12083__A2 net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07263__A1_N net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09302__A _04591_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14916__Q team_03_WB.instance_to_wrap.CPU_DAT_O\[3\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_12707_ net1374 vssd1 vssd1 vccd1 vccd1 _00471_ sky130_fd_sc_hd__inv_2
XFILLER_0_167_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07495__C1 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13687_ clknet_leaf_111_wb_clk_i _01451_ _00052_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[41\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10899_ net271 net2039 net520 vssd1 vssd1 vccd1 vccd1 _02320_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12638_ net1387 vssd1 vssd1 vccd1 vccd1 _00402_ sky130_fd_sc_hd__inv_2
XFILLER_0_155_487 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09787__A1 _02954_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11978__S net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12569_ net1355 vssd1 vssd1 vccd1 vccd1 _00333_ sky130_fd_sc_hd__inv_2
XFILLER_0_13_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_117_2773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14308_ clknet_leaf_15_wb_clk_i _02072_ _00673_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[662\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold206 team_03_WB.instance_to_wrap.ADR_I\[29\] vssd1 vssd1 vccd1 vccd1 net1699 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10794__A_N _05799_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08352__S net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_2784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold217 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[12\] vssd1 vssd1 vccd1
+ vccd1 net1710 sky130_fd_sc_hd__dlygate4sd3_1
Xhold228 team_03_WB.instance_to_wrap.CPU_DAT_I\[9\] vssd1 vssd1 vccd1 vccd1 net1721
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_151_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_170_Left_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11279__A net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold239 net197 vssd1 vssd1 vccd1 vccd1 net1732 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_169_3840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14239_ clknet_leaf_171_wb_clk_i _02003_ _00604_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[593\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_169_3851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11346__A1 net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08747__C1 net1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08211__A1 net1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout708 _06461_ vssd1 vssd1 vccd1 vccd1 net708 sky130_fd_sc_hd__buf_4
XFILLER_0_21_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08211__B2 net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout719 net720 vssd1 vssd1 vccd1 vccd1 net719 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_165_3759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13494__A net1328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08800_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[1\] net1008
+ net927 _04741_ vssd1 vssd1 vccd1 vccd1 _04742_ sky130_fd_sc_hd__o211a_1
XFILLER_0_42_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09691__B _05632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09780_ _04649_ _04895_ _04956_ _05071_ net566 net561 vssd1 vssd1 vccd1 vccd1 _05722_
+ sky130_fd_sc_hd__mux4_1
X_06992_ _02829_ _02836_ _02928_ _02933_ vssd1 vssd1 vccd1 vccd1 _02934_ sky130_fd_sc_hd__or4bb_2
XPHY_EDGE_ROW_7_Right_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08731_ net1050 team_03_WB.instance_to_wrap.core.register_file.registers_state\[964\]
+ net1013 team_03_WB.instance_to_wrap.core.register_file.registers_state\[996\] net1067
+ vssd1 vssd1 vccd1 vccd1 _04673_ sky130_fd_sc_hd__a221o_1
XFILLER_0_56_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11218__S net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1290 net1291 vssd1 vssd1 vccd1 vccd1 net1290 sky130_fd_sc_hd__buf_4
XANTENNA_clkbuf_leaf_89_wb_clk_i_A clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09711__B2 _02804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08662_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[423\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[391\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[295\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[263\]
+ net990 net1078 vssd1 vssd1 vccd1 vccd1 _04604_ sky130_fd_sc_hd__mux4_1
XANTENNA__07846__A1_N net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07613_ net1205 team_03_WB.instance_to_wrap.core.register_file.registers_state\[857\]
+ net788 team_03_WB.instance_to_wrap.core.register_file.registers_state\[889\] net1168
+ vssd1 vssd1 vccd1 vccd1 _03555_ sky130_fd_sc_hd__o221a_1
X_08593_ _04478_ _04534_ net553 vssd1 vssd1 vccd1 vccd1 _04535_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_511 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07544_ _03481_ _03485_ _03484_ net1122 vssd1 vssd1 vccd1 vccd1 _03486_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__12074__A2 net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_158_270 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11282__B1 net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07475_ net1184 team_03_WB.instance_to_wrap.core.register_file.registers_state\[853\]
+ net769 team_03_WB.instance_to_wrap.core.register_file.registers_state\[885\] net1129
+ vssd1 vssd1 vccd1 vccd1 _03417_ sky130_fd_sc_hd__o221a_1
XFILLER_0_8_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12049__S net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout333_A _06809_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_808 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1075_A net1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_763 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09214_ _02937_ _05155_ vssd1 vssd1 vccd1 vccd1 _05156_ sky130_fd_sc_hd__and2_1
XFILLER_0_5_1094 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09145_ net432 net425 _04323_ net549 vssd1 vssd1 vccd1 vccd1 _05087_ sky130_fd_sc_hd__o31a_1
XANTENNA_fanout500_A net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06842__Y _02785_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12007__D_N net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1242_A net1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08986__C1 net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_20_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09076_ net1240 team_03_WB.instance_to_wrap.core.register_file.registers_state\[77\]
+ net982 team_03_WB.instance_to_wrap.core.register_file.registers_state\[109\] net926
+ vssd1 vssd1 vccd1 vccd1 _05018_ sky130_fd_sc_hd__o221a_1
XFILLER_0_130_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08027_ net1085 team_03_WB.instance_to_wrap.core.register_file.registers_state\[241\]
+ net890 vssd1 vssd1 vccd1 vccd1 _03969_ sky130_fd_sc_hd__or3_1
XANTENNA__07386__B net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1030_X net1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_855 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold740 team_03_WB.instance_to_wrap.core.register_file.registers_state\[470\] vssd1
+ vssd1 vccd1 vccd1 net2233 sky130_fd_sc_hd__dlygate4sd3_1
Xhold751 team_03_WB.instance_to_wrap.core.register_file.registers_state\[800\] vssd1
+ vssd1 vccd1 vccd1 net2244 sky130_fd_sc_hd__dlygate4sd3_1
Xhold762 team_03_WB.instance_to_wrap.core.register_file.registers_state\[888\] vssd1
+ vssd1 vccd1 vccd1 net2255 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1128_X net1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09882__A _05596_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold773 team_03_WB.instance_to_wrap.core.register_file.registers_state\[905\] vssd1
+ vssd1 vccd1 vccd1 net2266 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout490_X net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold784 team_03_WB.instance_to_wrap.core.register_file.registers_state\[489\] vssd1
+ vssd1 vccd1 vccd1 net2277 sky130_fd_sc_hd__dlygate4sd3_1
Xhold795 team_03_WB.instance_to_wrap.core.register_file.registers_state\[812\] vssd1
+ vssd1 vccd1 vccd1 net2288 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11339__D net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout967_A net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_89_wb_clk_i clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_89_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_09978_ _03023_ net1760 net291 vssd1 vssd1 vccd1 vccd1 _02735_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_51_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10560__A2 net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09093__S net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_18_wb_clk_i clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_18_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_08929_ _04867_ _04870_ net868 vssd1 vssd1 vccd1 vccd1 _04871_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout755_X net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09702__A1 _05073_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09702__B2 _04777_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11940_ _06633_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[192\]
+ net369 vssd1 vssd1 vccd1 vccd1 _01602_ sky130_fd_sc_hd__mux2_1
XANTENNA__11355__C net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11871_ net268 net2139 net377 vssd1 vssd1 vccd1 vccd1 _01669_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout922_X net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_179 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13610_ net1316 vssd1 vssd1 vccd1 vccd1 _01374_ sky130_fd_sc_hd__inv_2
XFILLER_0_157_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10822_ net278 net2610 net519 vssd1 vssd1 vccd1 vccd1 _02332_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14590_ clknet_leaf_115_wb_clk_i _02354_ _00955_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[944\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_39_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_49_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08437__S net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13541_ net1329 vssd1 vssd1 vccd1 vccd1 _01305_ sky130_fd_sc_hd__inv_2
XANTENNA__11371__B net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08364__S1 net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10753_ _05746_ net604 vssd1 vssd1 vccd1 vccd1 _06370_ sky130_fd_sc_hd__nand2_1
XFILLER_0_82_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11812__A2 net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13472_ net1321 vssd1 vssd1 vccd1 vccd1 _01236_ sky130_fd_sc_hd__inv_2
XFILLER_0_138_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input96_A wbs_adr_i[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10684_ _05429_ _06313_ vssd1 vssd1 vccd1 vccd1 _06325_ sky130_fd_sc_hd__or2_1
XFILLER_0_109_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_936 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11798__S net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12423_ net1368 vssd1 vssd1 vccd1 vccd1 _00187_ sky130_fd_sc_hd__inv_2
XFILLER_0_164_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_1124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10555__X _06298_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_97_2367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_97_2378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_608 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12354_ net1360 vssd1 vssd1 vccd1 vccd1 _00118_ sky130_fd_sc_hd__inv_2
XFILLER_0_50_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_991 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10715__B net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11099__A net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11305_ _06615_ net2750 net405 vssd1 vssd1 vccd1 vccd1 _02140_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_75_1920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15073_ net1459 vssd1 vssd1 vccd1 vccd1 la_data_out[9] sky130_fd_sc_hd__buf_2
XFILLER_0_132_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_855 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12285_ net1383 vssd1 vssd1 vccd1 vccd1 _00049_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_147_3401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14024_ clknet_leaf_8_wb_clk_i _01788_ _00389_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[378\]
+ sky130_fd_sc_hd__dfrtp_1
X_11236_ net490 net618 _06685_ net408 net2343 vssd1 vssd1 vccd1 vccd1 _02177_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_112_2670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_123_wb_clk_i_A clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_1839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11167_ _06562_ net713 net297 vssd1 vssd1 vccd1 vccd1 _06662_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_143_3309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10551__A2 _06293_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10118_ _05960_ net2753 _05947_ vssd1 vssd1 vccd1 vccd1 _02666_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11098_ _06625_ net2441 net418 vssd1 vssd1 vccd1 vccd1 _02255_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_1076 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_160_3656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14926_ clknet_leaf_62_wb_clk_i _02681_ _01291_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_O\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_10049_ net7 net1039 net911 net2781 vssd1 vssd1 vccd1 vccd1 _02682_ sky130_fd_sc_hd__a22o_1
XANTENNA__11265__C net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_160_3667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08901__C1 net1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14857_ clknet_leaf_57_wb_clk_i _02621_ _01222_ vssd1 vssd1 vccd1 vccd1 net112 sky130_fd_sc_hd__dfrtp_2
XANTENNA__10877__S net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06927__Y _02869_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_6_wb_clk_i_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_58_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12658__A net1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13808_ clknet_leaf_121_wb_clk_i _01572_ _00173_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[162\]
+ sky130_fd_sc_hd__dfrtp_1
X_14788_ clknet_leaf_102_wb_clk_i _02552_ _01153_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_I\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11264__B1 net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07468__C1 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13739_ clknet_leaf_41_wb_clk_i _01503_ _00104_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[93\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10178__A _03242_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_728 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_2813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09967__A _03788_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_2824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07260_ net1131 _03198_ _03199_ net1119 vssd1 vssd1 vccd1 vccd1 _03202_ sky130_fd_sc_hd__a31o_1
XFILLER_0_144_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11016__B1 net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_324 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13489__A net1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07191_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[883\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[851\]
+ net762 vssd1 vssd1 vccd1 vccd1 _03133_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11501__S net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07487__A _03391_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_162_wb_clk_i_A clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__08968__C1 net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07235__A2 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08432__A1 net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08983__A2 net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09901_ _05834_ _05841_ _05833_ vssd1 vssd1 vccd1 vccd1 _05843_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_10_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_190 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout505 net506 vssd1 vssd1 vccd1 vccd1 net505 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11159__D net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout516 net517 vssd1 vssd1 vccd1 vccd1 net516 sky130_fd_sc_hd__buf_4
XFILLER_0_10_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout527 net528 vssd1 vssd1 vccd1 vccd1 net527 sky130_fd_sc_hd__clkbuf_4
X_09832_ net579 _04711_ net537 _05773_ vssd1 vssd1 vccd1 vccd1 _05774_ sky130_fd_sc_hd__o31a_1
XPHY_EDGE_ROW_171_Right_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout538 net539 vssd1 vssd1 vccd1 vccd1 net538 sky130_fd_sc_hd__buf_2
XFILLER_0_158_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08291__S0 net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout549 _03105_ vssd1 vssd1 vccd1 vccd1 net549 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07943__B1 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09763_ net351 _05463_ _05704_ vssd1 vssd1 vccd1 vccd1 _05705_ sky130_fd_sc_hd__a21oi_1
X_06975_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[517\] net805
+ vssd1 vssd1 vccd1 vccd1 _02917_ sky130_fd_sc_hd__or2_1
XANTENNA__08111__A net1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout283_A net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08714_ net1059 team_03_WB.instance_to_wrap.core.register_file.registers_state\[196\]
+ net1013 team_03_WB.instance_to_wrap.core.register_file.registers_state\[228\] net928
+ vssd1 vssd1 vccd1 vccd1 _04656_ sky130_fd_sc_hd__a221o_1
X_09694_ _05196_ _05203_ _05635_ vssd1 vssd1 vccd1 vccd1 _05636_ sky130_fd_sc_hd__or3_1
XFILLER_0_83_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15065__1451 vssd1 vssd1 vccd1 vccd1 _15065__1451/HI net1451 sky130_fd_sc_hd__conb_1
XFILLER_0_174_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09160__A2 _04476_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07950__A net1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08594__S1 net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08645_ net1053 team_03_WB.instance_to_wrap.core.register_file.registers_state\[582\]
+ net1006 team_03_WB.instance_to_wrap.core.register_file.registers_state\[614\] net941
+ vssd1 vssd1 vccd1 vccd1 _04587_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout450_A _06801_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07171__A1 net1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout548_A net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1192_A net1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08576_ _04512_ _04517_ net872 vssd1 vssd1 vccd1 vccd1 _04518_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_218 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10058__A1 net29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10058__B2 team_03_WB.instance_to_wrap.CPU_DAT_O\[5\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_119_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07527_ _03467_ _03468_ vssd1 vssd1 vccd1 vccd1 _03469_ sky130_fd_sc_hd__and2_1
XFILLER_0_77_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_136_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_136_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_76_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout715_A net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout336_X net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08120__B1 net1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1078_X net1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07458_ net744 _03398_ _03399_ net807 vssd1 vssd1 vccd1 vccd1 _03400_ sky130_fd_sc_hd__a31o_1
XFILLER_0_88_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08671__B2 net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_162_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07389_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[319\] net758
+ net1041 vssd1 vssd1 vccd1 vccd1 _03331_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout503_X net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1245_X net1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11411__S net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_150_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11558__B2 net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09128_ net436 net427 net588 net546 vssd1 vssd1 vccd1 vccd1 _05070_ sky130_fd_sc_hd__o31a_1
XFILLER_0_161_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_40_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09059_ _04999_ _05000_ net1064 vssd1 vssd1 vccd1 vccd1 _05001_ sky130_fd_sc_hd__a21o_1
XFILLER_0_102_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_92_2264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08005__B _03946_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_2275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12070_ net263 net1840 net357 vssd1 vssd1 vccd1 vccd1 _01476_ sky130_fd_sc_hd__mux2_1
Xhold570 team_03_WB.instance_to_wrap.core.register_file.registers_state\[33\] vssd1
+ vssd1 vccd1 vccd1 net2063 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout872_X net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold581 team_03_WB.instance_to_wrap.core.register_file.registers_state\[553\] vssd1
+ vssd1 vccd1 vccd1 net2074 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08187__B1 net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold592 team_03_WB.instance_to_wrap.core.register_file.registers_state\[282\] vssd1
+ vssd1 vccd1 vccd1 net2085 sky130_fd_sc_hd__dlygate4sd3_1
X_11021_ net2480 net420 _06584_ net496 vssd1 vssd1 vccd1 vccd1 _02291_ sky130_fd_sc_hd__a22o_1
XFILLER_0_60_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10533__A2 net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11730__A1 net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09117__A net1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12972_ net1314 vssd1 vssd1 vccd1 vccd1 _00736_ sky130_fd_sc_hd__inv_2
Xhold1270 team_03_WB.instance_to_wrap.core.register_file.registers_state\[476\] vssd1
+ vssd1 vccd1 vccd1 net2763 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_input11_A DAT_I[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1281 team_03_WB.instance_to_wrap.wb.curr_state\[1\] vssd1 vssd1 vccd1 vccd1 net2774
+ sky130_fd_sc_hd__dlygate4sd3_1
X_14711_ clknet_leaf_32_wb_clk_i _02475_ _01076_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.decoder.inst\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_11923_ _06479_ net2395 net367 vssd1 vssd1 vccd1 vccd1 _01619_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14642_ clknet_leaf_121_wb_clk_i _02406_ _01007_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[996\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_157_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12038__A2 net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11854_ net274 net2010 net375 vssd1 vssd1 vccd1 vccd1 _01686_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10049__A1 net7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10805_ _06410_ _06411_ _06412_ vssd1 vssd1 vccd1 vccd1 _06413_ sky130_fd_sc_hd__a21oi_4
XANTENNA__08337__S1 net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11246__B1 net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14573_ clknet_leaf_190_wb_clk_i _02337_ _00938_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[927\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_99_2407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11785_ net2758 _06618_ net327 vssd1 vssd1 vccd1 vccd1 _01753_ sky130_fd_sc_hd__mux2_1
XANTENNA__11532__D net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_2418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11797__A1 _06505_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13524_ net1316 vssd1 vssd1 vccd1 vccd1 _01288_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_64_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10736_ team_03_WB.instance_to_wrap.core.pc.current_pc\[13\] _05659_ net605 vssd1
+ vssd1 vccd1 vccd1 _06360_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_24_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input99_X net99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_878 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_136_3168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_59 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13455_ net1343 vssd1 vssd1 vccd1 vccd1 _01219_ sky130_fd_sc_hd__inv_2
XFILLER_0_82_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10667_ net1142 _06305_ _06306_ _06308_ vssd1 vssd1 vccd1 vccd1 _06309_ sky130_fd_sc_hd__or4_4
XFILLER_0_125_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11549__A1 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11321__S net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12406_ net1280 vssd1 vssd1 vccd1 vccd1 _00170_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_114_2710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13386_ net1427 vssd1 vssd1 vccd1 vccd1 _01150_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10598_ net1708 team_03_WB.instance_to_wrap.CPU_DAT_O\[31\] net841 vssd1 vssd1 vccd1
+ vccd1 _02530_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_114_2721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15125_ net915 vssd1 vssd1 vccd1 vccd1 net256 sky130_fd_sc_hd__clkbuf_1
Xoutput108 net108 vssd1 vssd1 vccd1 vccd1 ADR_O[14] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_11_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12337_ net1265 vssd1 vssd1 vccd1 vccd1 _00101_ sky130_fd_sc_hd__inv_2
XFILLER_0_105_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput119 net119 vssd1 vssd1 vccd1 vccd1 ADR_O[24] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_121_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15056_ net1442 vssd1 vssd1 vccd1 vccd1 gpio_out[2] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_110_2629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12268_ net1331 vssd1 vssd1 vccd1 vccd1 _00032_ sky130_fd_sc_hd__inv_2
X_14007_ clknet_leaf_112_wb_clk_i _01771_ _00372_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[361\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11557__A net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11219_ net297 net2540 net488 vssd1 vssd1 vccd1 vccd1 _02190_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_162_3707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12199_ net1496 vssd1 vssd1 vccd1 vccd1 _02354_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__10524__A2 net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11721__A1 net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07246__S net1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11991__S net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14909_ clknet_leaf_54_wb_clk_i _00003_ _01274_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.ru.state\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_144_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_1022 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07689__C1 net1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07153__A1 net1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08430_ net1049 team_03_WB.instance_to_wrap.core.register_file.registers_state\[666\]
+ net1000 team_03_WB.instance_to_wrap.core.register_file.registers_state\[698\] net920
+ vssd1 vssd1 vccd1 vccd1 _04372_ sky130_fd_sc_hd__a221o_1
XFILLER_0_19_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08361_ net866 _04299_ _04302_ vssd1 vssd1 vccd1 vccd1 _04303_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_59_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11788__A1 _06454_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_160_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07312_ net1152 _03252_ _03253_ net822 vssd1 vssd1 vccd1 vccd1 _03254_ sky130_fd_sc_hd__o31a_1
XFILLER_0_129_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08292_ _04228_ _04233_ net872 vssd1 vssd1 vccd1 vccd1 _04234_ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10460__A1 net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07243_ net1191 team_03_WB.instance_to_wrap.core.register_file.registers_state\[584\]
+ net774 team_03_WB.instance_to_wrap.core.register_file.registers_state\[616\] net730
+ vssd1 vssd1 vccd1 vccd1 _03185_ sky130_fd_sc_hd__o221a_1
XFILLER_0_73_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_147_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11231__S net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_788 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07174_ net811 _03112_ _03115_ vssd1 vssd1 vccd1 vccd1 _03116_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_143_287 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08106__A net1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07010__A net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07613__C1 net1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10923__X _06511_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11960__A1 net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout302 _06422_ vssd1 vssd1 vccd1 vccd1 net302 sky130_fd_sc_hd__buf_2
XANTENNA_fanout498_A net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout313 _05387_ vssd1 vssd1 vccd1 vccd1 net313 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12062__S net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout324 _06811_ vssd1 vssd1 vccd1 vccd1 net324 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10515__A2 net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1205_A net1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11712__A1 _06409_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout335 net337 vssd1 vssd1 vccd1 vccd1 net335 sky130_fd_sc_hd__clkbuf_8
Xfanout346 _06804_ vssd1 vssd1 vccd1 vccd1 net346 sky130_fd_sc_hd__buf_6
XANTENNA__07916__B1 _02870_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09815_ _02954_ _05587_ _05749_ _05756_ vssd1 vssd1 vccd1 vccd1 _05757_ sky130_fd_sc_hd__a211o_4
XANTENNA_input3_A DAT_I[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout357 _06818_ vssd1 vssd1 vccd1 vccd1 net357 sky130_fd_sc_hd__buf_6
XANTENNA__11186__B net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10090__B _05632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout368 _06814_ vssd1 vssd1 vccd1 vccd1 net368 sky130_fd_sc_hd__buf_4
Xfanout379 net387 vssd1 vssd1 vccd1 vccd1 net379 sky130_fd_sc_hd__buf_4
XANTENNA_fanout286_X net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout665_A net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09746_ _05084_ _05086_ _05117_ _05119_ net555 net570 vssd1 vssd1 vccd1 vccd1 _05688_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_94_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09669__B1 _05610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06958_ net808 _02896_ _02899_ vssd1 vssd1 vccd1 vccd1 _02900_ sky130_fd_sc_hd__a21o_1
XFILLER_0_119_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09677_ _03391_ _04119_ net667 _05618_ vssd1 vssd1 vccd1 vccd1 _05619_ sky130_fd_sc_hd__a22o_1
XFILLER_0_119_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06889_ team_03_WB.instance_to_wrap.core.decoder.inst\[12\] _02820_ vssd1 vssd1 vccd1
+ vccd1 _02831_ sky130_fd_sc_hd__and2_2
XFILLER_0_55_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout453_X net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07144__A1 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout832_A _06387_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1195_X net1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11406__S net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08628_ _04568_ _04569_ net857 vssd1 vssd1 vccd1 vccd1 _04570_ sky130_fd_sc_hd__o21a_1
XFILLER_0_68_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11228__A0 _06532_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout620_X net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08559_ net1063 _04497_ _04500_ net870 vssd1 vssd1 vccd1 vccd1 _04501_ sky130_fd_sc_hd__a211o_1
XFILLER_0_76_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout718_X net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11570_ net636 net706 net267 net698 vssd1 vssd1 vccd1 vccd1 _06798_ sky130_fd_sc_hd__and4_1
XANTENNA__08644__A1 net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10521_ net145 net1031 net1023 net1779 vssd1 vssd1 vccd1 vccd1 _02589_ sky130_fd_sc_hd__a22o_1
XFILLER_0_162_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07852__C1 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_2304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_2315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13240_ net1380 vssd1 vssd1 vccd1 vccd1 _01004_ sky130_fd_sc_hd__inv_2
X_10452_ _05925_ net303 _06267_ vssd1 vssd1 vccd1 vccd1 _06268_ sky130_fd_sc_hd__and3_1
XFILLER_0_123_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_162_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08016__A net1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11400__A0 net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_3065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13171_ net1267 vssd1 vssd1 vccd1 vccd1 _00935_ sky130_fd_sc_hd__inv_2
XFILLER_0_62_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10383_ _05994_ _06085_ _05996_ _05992_ vssd1 vssd1 vccd1 vccd1 _06212_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_131_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06958__A1 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11951__A1 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_983 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12122_ net1532 vssd1 vssd1 vccd1 vccd1 _02431_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_33_wb_clk_i clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_33_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_20_447 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07080__B1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input59_A gpio_in[34] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11377__A net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12053_ _06469_ net2654 net355 vssd1 vssd1 vccd1 vccd1 _01493_ sky130_fd_sc_hd__mux2_1
XANTENNA__10506__A2 net1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11004_ net2255 net421 _06574_ net502 vssd1 vssd1 vccd1 vccd1 _02298_ sky130_fd_sc_hd__a22o_1
XANTENNA__07293__C net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09109__C1 net1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07383__A1 net1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08580__B1 net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout880 net887 vssd1 vssd1 vccd1 vccd1 net880 sky130_fd_sc_hd__clkbuf_4
Xfanout891 net904 vssd1 vssd1 vccd1 vccd1 net891 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_172_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09134__X _05076_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07590__A net1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input14_X net14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12955_ net1296 vssd1 vssd1 vccd1 vccd1 _00719_ sky130_fd_sc_hd__inv_2
XANTENNA__09675__A3 net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_2580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11316__S net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11906_ net636 _06715_ net470 net373 net2015 vssd1 vssd1 vccd1 vccd1 _01635_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_66_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12886_ net1258 vssd1 vssd1 vccd1 vccd1 _00650_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_138_3208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11219__A0 net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_3219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_158_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09788__Y _05730_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14625_ clknet_leaf_179_wb_clk_i _02389_ _00990_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[979\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_74_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11837_ net656 _06675_ net473 net325 net1939 vssd1 vssd1 vccd1 vccd1 _01702_ sky130_fd_sc_hd__a32o_1
XFILLER_0_96_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_2488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12936__A net1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_2499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14556_ clknet_leaf_151_wb_clk_i _02320_ _00921_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[910\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08096__C1 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_155_3555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11768_ _06601_ net478 net334 net2542 vssd1 vssd1 vccd1 vccd1 _01769_ sky130_fd_sc_hd__a22o_1
XFILLER_0_138_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_155_3566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10442__A1 _05925_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09310__A net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14924__Q team_03_WB.instance_to_wrap.CPU_DAT_O\[11\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_10719_ _05596_ net602 vssd1 vssd1 vccd1 vccd1 _06351_ sky130_fd_sc_hd__nand2_1
X_13507_ net1322 vssd1 vssd1 vccd1 vccd1 _01271_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14487_ clknet_leaf_79_wb_clk_i _02251_ _00852_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[841\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11699_ _06741_ net385 net341 net1869 vssd1 vssd1 vccd1 vccd1 _01835_ sky130_fd_sc_hd__a22o_1
XANTENNA__10993__A2 net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13438_ net1423 vssd1 vssd1 vccd1 vccd1 _01202_ sky130_fd_sc_hd__inv_2
XFILLER_0_153_596 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08399__B1 net992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11986__S net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15064__1450 vssd1 vssd1 vccd1 vccd1 _15064__1450/HI net1450 sky130_fd_sc_hd__conb_1
XFILLER_0_106_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_658 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13369_ net1322 vssd1 vssd1 vccd1 vccd1 _01133_ sky130_fd_sc_hd__inv_2
XANTENNA__09060__A1 net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06949__A1 net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09060__B2 net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11942__A1 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15108_ net914 vssd1 vssd1 vccd1 vccd1 net243 sky130_fd_sc_hd__clkbuf_1
XANTENNA__07071__B1 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11287__A net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15039_ clknet_leaf_81_wb_clk_i _02759_ _01404_ vssd1 vssd1 vccd1 vccd1 net195 sky130_fd_sc_hd__dfrtp_1
X_07930_ net1181 team_03_WB.instance_to_wrap.core.register_file.registers_state\[87\]
+ net766 team_03_WB.instance_to_wrap.core.register_file.registers_state\[119\] net728
+ vssd1 vssd1 vccd1 vccd1 _03872_ sky130_fd_sc_hd__o221a_1
X_07861_ net1108 team_03_WB.instance_to_wrap.core.register_file.registers_state\[667\]
+ net737 _03791_ vssd1 vssd1 vccd1 vccd1 _03803_ sky130_fd_sc_hd__a211o_1
X_09600_ _05541_ _05500_ _05518_ vssd1 vssd1 vccd1 vccd1 _05542_ sky130_fd_sc_hd__and3b_1
XANTENNA__08571__B1 net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07792_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[683\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[651\]
+ net775 vssd1 vssd1 vccd1 vccd1 _03734_ sky130_fd_sc_hd__mux2_1
XANTENNA__08596__A _02954_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_2978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09531_ _03566_ _04354_ net538 vssd1 vssd1 vccd1 vccd1 _05473_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_127_2989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07931__C net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11226__S net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10130__A0 _04415_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09462_ _05397_ _05403_ net580 vssd1 vssd1 vccd1 vccd1 _05404_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_148_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08413_ net432 net424 _04354_ net547 vssd1 vssd1 vccd1 vccd1 _04355_ sky130_fd_sc_hd__o31a_1
X_09393_ _05318_ _05333_ _05334_ vssd1 vssd1 vccd1 vccd1 _05335_ sky130_fd_sc_hd__or3b_2
XFILLER_0_46_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_171 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08344_ net855 _04284_ _04285_ vssd1 vssd1 vccd1 vccd1 _04286_ sky130_fd_sc_hd__or3_1
XFILLER_0_19_547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07429__A2 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_867 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09858__C _05798_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06844__A net1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10364__A2_N net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1096 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_303 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11630__B1 net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08275_ net855 _04215_ _04216_ _04214_ vssd1 vssd1 vccd1 vccd1 _04217_ sky130_fd_sc_hd__o31a_1
XANTENNA__12057__S net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout413_A _06635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1155_A net1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_574 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07226_ net1146 _03159_ _03167_ vssd1 vssd1 vccd1 vccd1 _03168_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_171_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_71 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09051__A1 net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07157_ net1203 team_03_WB.instance_to_wrap.core.register_file.registers_state\[288\]
+ net885 _02872_ vssd1 vssd1 vccd1 vccd1 _03099_ sky130_fd_sc_hd__a31o_1
XFILLER_0_15_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07088_ net747 _03028_ _03029_ net1165 vssd1 vssd1 vccd1 vccd1 _03030_ sky130_fd_sc_hd__a31o_1
XFILLER_0_140_791 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout782_A net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1108 net1113 vssd1 vssd1 vccd1 vccd1 net1108 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_121_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1208_X net1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1119 net1122 vssd1 vssd1 vccd1 vccd1 net1119 sky130_fd_sc_hd__buf_4
XFILLER_0_10_480 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input6_X net6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11697__B1 net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11161__A2 net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout668_X net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09729_ _04150_ _04269_ _04326_ _04386_ net563 net560 vssd1 vssd1 vccd1 vccd1 _05671_
+ sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_151_wb_clk_i clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_151_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout835_X net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07117__A1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08314__B1 net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12740_ net1382 vssd1 vssd1 vccd1 vccd1 _00504_ sky130_fd_sc_hd__inv_2
XFILLER_0_69_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11363__C net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08865__A1 net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12671_ net1350 vssd1 vssd1 vccd1 vccd1 _00435_ sky130_fd_sc_hd__inv_2
XANTENNA__12756__A net1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14410_ clknet_leaf_1_wb_clk_i _02174_ _00775_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[764\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_93_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11622_ _06696_ net380 net346 net2579 vssd1 vssd1 vccd1 vccd1 _01910_ sky130_fd_sc_hd__a22o_1
XFILLER_0_155_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08617__A1 net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_3105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14341_ clknet_leaf_37_wb_clk_i _02105_ _00706_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[695\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_170_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_133_3116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11553_ net2612 net484 _06791_ net507 vssd1 vssd1 vccd1 vccd1 _01966_ sky130_fd_sc_hd__a22o_1
XANTENNA__11621__B1 net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10504_ net125 net1033 net908 net1761 vssd1 vssd1 vccd1 vccd1 _02605_ sky130_fd_sc_hd__a22o_1
X_14272_ clknet_leaf_191_wb_clk_i _02036_ _00637_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[626\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_150_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11484_ net636 net705 _06550_ net829 vssd1 vssd1 vccd1 vccd1 _06776_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_150_3452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_150_3463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_758 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xwire588 _05068_ vssd1 vssd1 vccd1 vccd1 net588 sky130_fd_sc_hd__buf_4
X_13223_ net1399 vssd1 vssd1 vccd1 vccd1 _00987_ sky130_fd_sc_hd__inv_2
X_10435_ _06253_ _06254_ team_03_WB.instance_to_wrap.core.pc.current_pc\[9\] net682
+ vssd1 vssd1 vccd1 vccd1 _02643_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_150_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_572 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12491__A net1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09042__A1 net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10727__A2 net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_211 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_49 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07585__A team_03_WB.instance_to_wrap.core.decoder.inst\[24\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08180__S net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_628 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13154_ net1289 vssd1 vssd1 vccd1 vccd1 _00918_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_59_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10366_ _05981_ _06089_ _06094_ vssd1 vssd1 vccd1 vccd1 _06198_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_27_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_29_Left_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12105_ _06799_ net477 net442 net2165 vssd1 vssd1 vccd1 vccd1 _01442_ sky130_fd_sc_hd__a22o_1
X_13085_ net1388 vssd1 vssd1 vccd1 vccd1 _00849_ sky130_fd_sc_hd__inv_2
X_10297_ team_03_WB.instance_to_wrap.core.pc.current_pc\[10\] _06138_ vssd1 vssd1
+ vccd1 vccd1 _06139_ sky130_fd_sc_hd__and2_1
X_12036_ _06775_ net471 net361 net2295 vssd1 vssd1 vccd1 vccd1 _01509_ sky130_fd_sc_hd__a22o_1
XANTENNA__11688__B1 net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_2620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07356__A1 net1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_67 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06929__A net1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09728__S0 net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09305__A net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14919__Q team_03_WB.instance_to_wrap.CPU_DAT_O\[6\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__07751__C net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_2528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12101__A1 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13987_ clknet_leaf_36_wb_clk_i _01751_ _00352_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[341\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08305__B1 net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11273__C net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12938_ net1283 vssd1 vssd1 vccd1 vccd1 _00702_ sky130_fd_sc_hd__inv_2
XFILLER_0_34_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_157_3606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_38_Left_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_406 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_122_2875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11860__A0 net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1085 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_122_2886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09959__B net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12869_ net1349 vssd1 vssd1 vccd1 vccd1 _00633_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_174_3942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11570__A net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08608__A1 net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14608_ clknet_leaf_157_wb_clk_i _02372_ _00973_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[962\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_174_3953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08355__S net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_174_3964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_174_3975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09040__A net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_390 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11612__B1 net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14539_ clknet_leaf_46_wb_clk_i _02303_ _00904_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[893\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08084__A2 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10966__A2 net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07292__B1 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08060_ net1186 team_03_WB.instance_to_wrap.core.register_file.registers_state\[470\]
+ vssd1 vssd1 vccd1 vccd1 _04002_ sky130_fd_sc_hd__or2_1
XFILLER_0_114_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_153_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07011_ net526 _02944_ _02948_ _02952_ vssd1 vssd1 vccd1 vccd1 _02953_ sky130_fd_sc_hd__and4_2
XFILLER_0_12_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13497__A net1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09033__A1 net1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10914__A _06503_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12040__D_N net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_47_Left_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07926__C net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08962_ net1245 team_03_WB.instance_to_wrap.core.register_file.registers_state\[457\]
+ net986 team_03_WB.instance_to_wrap.core.register_file.registers_state\[489\] net1216
+ vssd1 vssd1 vccd1 vccd1 _04904_ sky130_fd_sc_hd__o221a_1
XANTENNA__11448__C net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08878__X _04820_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07782__X _03724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07913_ net1085 team_03_WB.instance_to_wrap.core.register_file.registers_state\[975\]
+ vssd1 vssd1 vccd1 vccd1 _03855_ sky130_fd_sc_hd__and2_1
XANTENNA__11679__B1 net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08893_ _02795_ _02796_ net980 vssd1 vssd1 vccd1 vccd1 _04835_ sky130_fd_sc_hd__mux2_1
XANTENNA__10920__Y _06509_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07347__A1 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07844_ _03781_ _03782_ net739 vssd1 vssd1 vccd1 vccd1 _03786_ sky130_fd_sc_hd__mux2_1
XFILLER_0_166_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06839__A team_03_WB.instance_to_wrap.core.decoder.inst\[31\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07898__A2 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07775_ net1194 team_03_WB.instance_to_wrap.core.register_file.registers_state\[556\]
+ net883 vssd1 vssd1 vccd1 vccd1 _03717_ sky130_fd_sc_hd__and3_1
XFILLER_0_155_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout363_A _06815_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09514_ _05327_ _05430_ _05325_ vssd1 vssd1 vccd1 vccd1 _05456_ sky130_fd_sc_hd__o21a_1
XPHY_EDGE_ROW_56_Left_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09445_ _05346_ _05347_ _05386_ vssd1 vssd1 vccd1 vccd1 _05387_ sky130_fd_sc_hd__a21oi_2
XANTENNA__10654__A1 team_03_WB.instance_to_wrap.CPU_DAT_O\[7\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_66_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_2060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11851__A0 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout530_A _06309_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_2071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout628_A net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06845__Y _02788_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1272_A net1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_688 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09376_ _04445_ _05317_ vssd1 vssd1 vccd1 vccd1 _05318_ sky130_fd_sc_hd__and2_1
XANTENNA__08265__S net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11603__A0 _06536_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08327_ net548 _04237_ _04268_ vssd1 vssd1 vccd1 vccd1 _04269_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_152_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07807__C1 net1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10096__A net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1060_X net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout416_X net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_703 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1158_X net1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_954 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08258_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[818\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[786\]
+ net951 vssd1 vssd1 vccd1 vccd1 _04200_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_596 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08480__C1 net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout997_A _04085_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07209_ net1160 _03149_ _03150_ vssd1 vssd1 vccd1 vccd1 _03151_ sky130_fd_sc_hd__o21ai_1
XPHY_EDGE_ROW_65_Left_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09024__A1 net1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_566 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08189_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[435\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[403\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[307\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[275\]
+ net958 net1071 vssd1 vssd1 vccd1 vccd1 _04131_ sky130_fd_sc_hd__mux4_1
XFILLER_0_30_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11906__A1 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09096__S net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10220_ _06057_ _06059_ _06022_ _06024_ vssd1 vssd1 vccd1 vccd1 _06062_ sky130_fd_sc_hd__a211o_1
XFILLER_0_160_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07609__S net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07035__B1 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11198__Y _06680_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout785_X net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11382__A2 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10151_ _04178_ team_03_WB.instance_to_wrap.core.pc.current_pc\[17\] net674 vssd1
+ vssd1 vccd1 vccd1 _05993_ sky130_fd_sc_hd__mux2_1
XANTENNA__09891__Y _05833_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_89_2203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_2214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10082_ _05768_ _05784_ _05798_ vssd1 vssd1 vccd1 vccd1 _05926_ sky130_fd_sc_hd__and3_1
XANTENNA__07338__A1 _03279_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10830__Y _06433_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout952_X net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13910_ clknet_leaf_176_wb_clk_i _01674_ _00275_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[264\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_96_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14890_ clknet_leaf_58_wb_clk_i _02653_ _01255_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.pc.current_pc\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13841_ clknet_leaf_139_wb_clk_i _01605_ _00206_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[195\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_159_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12095__B1 net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13772_ clknet_leaf_19_wb_clk_i _01536_ _00137_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[126\]
+ sky130_fd_sc_hd__dfrtp_1
X_10984_ net1251 net833 vssd1 vssd1 vccd1 vccd1 _06562_ sky130_fd_sc_hd__or2_4
XANTENNA__08964__A net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10645__A1 team_03_WB.instance_to_wrap.CPU_DAT_O\[16\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_12723_ net1255 vssd1 vssd1 vccd1 vccd1 _00487_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_100_2425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06944__S0 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_2436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12654_ net1274 vssd1 vssd1 vccd1 vccd1 _00418_ sky130_fd_sc_hd__inv_2
XFILLER_0_66_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_675 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_152_3503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11605_ _06545_ net2366 net449 vssd1 vssd1 vccd1 vccd1 _01924_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12585_ net1253 vssd1 vssd1 vccd1 vccd1 _00349_ sky130_fd_sc_hd__inv_2
XFILLER_0_92_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09795__A net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14324_ clknet_leaf_133_wb_clk_i _02088_ _00689_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[678\]
+ sky130_fd_sc_hd__dfrtp_1
X_11536_ net627 _06646_ vssd1 vssd1 vccd1 vccd1 _06786_ sky130_fd_sc_hd__and2_1
XFILLER_0_81_976 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14255_ clknet_leaf_136_wb_clk_i _02019_ _00620_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[609\]
+ sky130_fd_sc_hd__dfrtp_1
X_11467_ net2301 net393 _06769_ net507 vssd1 vssd1 vccd1 vccd1 _02030_ sky130_fd_sc_hd__a22o_1
XFILLER_0_80_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_78_1973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13206_ net1257 vssd1 vssd1 vccd1 vccd1 _00970_ sky130_fd_sc_hd__inv_2
X_10418_ net284 _06140_ _06238_ net682 vssd1 vssd1 vccd1 vccd1 _06241_ sky130_fd_sc_hd__o31a_1
XFILLER_0_123_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_78_1984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09110__S1 net1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14186_ clknet_leaf_5_wb_clk_i _01950_ _00551_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[540\]
+ sky130_fd_sc_hd__dfrtp_1
X_11398_ _06449_ _06751_ vssd1 vssd1 vccd1 vccd1 _06752_ sky130_fd_sc_hd__or2_4
XANTENNA__08204__A net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07577__A1 net1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08774__B1 net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13137_ net1268 vssd1 vssd1 vccd1 vccd1 _00901_ sky130_fd_sc_hd__inv_2
X_10349_ _02771_ _06148_ vssd1 vssd1 vccd1 vccd1 _06184_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10581__B1 net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13068_ net1314 vssd1 vssd1 vccd1 vccd1 _00832_ sky130_fd_sc_hd__inv_2
XFILLER_0_40_1051 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11125__A2 net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12019_ net625 _06580_ net455 net359 net2235 vssd1 vssd1 vccd1 vccd1 _01526_ sky130_fd_sc_hd__a32o_1
XFILLER_0_136_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_79_wb_clk_i_A clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_2915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10884__A1 net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12086__B1 net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07560_ net1188 team_03_WB.instance_to_wrap.core.register_file.registers_state\[472\]
+ net772 team_03_WB.instance_to_wrap.core.register_file.registers_state\[504\] net1153
+ vssd1 vssd1 vccd1 vccd1 _03502_ sky130_fd_sc_hd__o221a_1
XFILLER_0_49_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11428__A3 _06756_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06946__X _02888_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11833__B1 net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07491_ _03431_ _03432_ vssd1 vssd1 vccd1 vccd1 _03433_ sky130_fd_sc_hd__and2_1
XFILLER_0_75_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_174_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09230_ _04532_ _05169_ vssd1 vssd1 vccd1 vccd1 _05172_ sky130_fd_sc_hd__and2_2
XANTENNA__11504__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09161_ net438 net424 _04532_ net541 vssd1 vssd1 vccd1 vccd1 _05103_ sky130_fd_sc_hd__o31a_1
XFILLER_0_17_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_161_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_883 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08112_ net1173 team_03_WB.instance_to_wrap.core.register_file.registers_state\[698\]
+ net876 vssd1 vssd1 vccd1 vccd1 _04054_ sky130_fd_sc_hd__and3_1
XFILLER_0_71_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_154_680 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09092_ net1208 _05030_ _05033_ vssd1 vssd1 vccd1 vccd1 _05034_ sky130_fd_sc_hd__or3_1
XFILLER_0_71_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08813__S net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10915__Y _06505_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11299__X _06717_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08043_ net1212 _02821_ _03107_ vssd1 vssd1 vccd1 vccd1 _03985_ sky130_fd_sc_hd__a21o_2
XANTENNA__09006__A1 net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09006__B2 net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold900 team_03_WB.instance_to_wrap.core.register_file.registers_state\[534\] vssd1
+ vssd1 vccd1 vccd1 net2393 sky130_fd_sc_hd__dlygate4sd3_1
Xhold911 team_03_WB.instance_to_wrap.core.register_file.registers_state\[875\] vssd1
+ vssd1 vccd1 vccd1 net2404 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13020__A net1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_263 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold922 team_03_WB.instance_to_wrap.core.register_file.registers_state\[120\] vssd1
+ vssd1 vccd1 vccd1 net2415 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12010__B1 net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08214__C1 net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold933 team_03_WB.instance_to_wrap.core.register_file.registers_state\[382\] vssd1
+ vssd1 vccd1 vccd1 net2426 sky130_fd_sc_hd__dlygate4sd3_1
Xhold944 team_03_WB.instance_to_wrap.core.register_file.registers_state\[625\] vssd1
+ vssd1 vccd1 vccd1 net2437 sky130_fd_sc_hd__dlygate4sd3_1
Xhold955 team_03_WB.instance_to_wrap.core.register_file.registers_state\[138\] vssd1
+ vssd1 vccd1 vccd1 net2448 sky130_fd_sc_hd__dlygate4sd3_1
Xhold966 team_03_WB.instance_to_wrap.core.register_file.registers_state\[479\] vssd1
+ vssd1 vccd1 vccd1 net2459 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08765__B1 net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11364__A2 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold977 team_03_WB.instance_to_wrap.core.register_file.registers_state\[498\] vssd1
+ vssd1 vccd1 vccd1 net2470 sky130_fd_sc_hd__dlygate4sd3_1
X_09994_ _05879_ net1867 net288 vssd1 vssd1 vccd1 vccd1 _02720_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout1020_A net1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold988 team_03_WB.instance_to_wrap.core.register_file.registers_state\[597\] vssd1
+ vssd1 vccd1 vccd1 net2481 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11178__C net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10572__B1 net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold999 team_03_WB.instance_to_wrap.core.register_file.registers_state\[668\] vssd1
+ vssd1 vccd1 vccd1 net2492 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10082__C _05798_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1118_A net1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08945_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[555\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[523\]
+ net977 vssd1 vssd1 vccd1 vccd1 _04887_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout480_A net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout578_A _02993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11475__A net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12070__S net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08876_ _02831_ _02929_ _02935_ vssd1 vssd1 vccd1 vccd1 _04818_ sky130_fd_sc_hd__or3b_2
XTAP_TAPCELL_ROW_32_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09190__B1 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10875__A1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11194__B net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07827_ net1171 team_03_WB.instance_to_wrap.core.register_file.registers_state\[362\]
+ net880 vssd1 vssd1 vccd1 vccd1 _03769_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_84_2100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout745_A net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout366_X net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07758_ net818 _03699_ vssd1 vssd1 vccd1 vccd1 _03700_ sky130_fd_sc_hd__nor2_1
XANTENNA__12077__B1 net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10627__A1 team_03_WB.instance_to_wrap.CPU_DAT_O\[2\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_2019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11824__B1 net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout533_X net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07689_ net1183 team_03_WB.instance_to_wrap.core.register_file.registers_state\[990\]
+ net766 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1022\] net1149
+ vssd1 vssd1 vccd1 vccd1 _03631_ sky130_fd_sc_hd__o221a_1
XFILLER_0_94_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09428_ _04832_ _05368_ _05369_ _05364_ vssd1 vssd1 vccd1 vccd1 _05370_ sky130_fd_sc_hd__o211a_1
XFILLER_0_17_1086 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09359_ _05291_ _05296_ _05300_ vssd1 vssd1 vccd1 vccd1 _05301_ sky130_fd_sc_hd__or3_2
XANTENNA_fanout700_X net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08048__A2 _03946_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_168 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11052__A1 net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12370_ net1395 vssd1 vssd1 vccd1 vccd1 _00134_ sky130_fd_sc_hd__inv_2
XANTENNA__08453__C1 net1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11321_ _06627_ net2627 net404 vssd1 vssd1 vccd1 vccd1 _02124_ sky130_fd_sc_hd__mux2_1
XANTENNA__07847__B net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1052 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12001__A0 net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14040_ clknet_leaf_172_wb_clk_i _01804_ _00405_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[394\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09548__A2 _04267_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11252_ net497 net626 _06693_ net409 net2062 vssd1 vssd1 vccd1 vccd1 _02169_ sky130_fd_sc_hd__a32o_1
XANTENNA__11369__B net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07559__A1 net1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_56_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10203_ team_03_WB.instance_to_wrap.core.pc.current_pc\[2\] net660 vssd1 vssd1 vccd1
+ vccd1 _06045_ sky130_fd_sc_hd__nor2_1
XANTENNA__08756__B1 net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_113_wb_clk_i_A clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__10841__X _06442_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_3004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11183_ net2344 net415 _06672_ net514 vssd1 vssd1 vccd1 vccd1 _02217_ sky130_fd_sc_hd__a22o_1
XANTENNA__10563__B1 net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_761 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08959__A net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10134_ _03565_ _05974_ vssd1 vssd1 vccd1 vccd1 _05976_ sky130_fd_sc_hd__nor2_1
XANTENNA_input41_A gpio_in[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07863__A net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_282 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08508__B1 net995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11385__A net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_3351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14942_ clknet_leaf_61_wb_clk_i _02697_ _01307_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_O\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_145_3362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10065_ team_03_WB.instance_to_wrap.core.decoder.inst\[24\] net1148 net1189 team_03_WB.instance_to_wrap.core.decoder.inst\[19\]
+ vssd1 vssd1 vccd1 vccd1 _05909_ sky130_fd_sc_hd__or4_1
XANTENNA__09126__Y _05068_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10866__A1 net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14873_ clknet_leaf_93_wb_clk_i _02636_ _01238_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.pc.current_pc\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA_output128_A net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12068__A0 net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13824_ clknet_leaf_190_wb_clk_i _01588_ _00189_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[178\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10618__A1 team_03_WB.instance_to_wrap.CPU_DAT_O\[11\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11815__B1 net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10967_ team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[1\] net306 vssd1 vssd1
+ vccd1 vccd1 _06547_ sky130_fd_sc_hd__nand2_2
X_13755_ clknet_leaf_122_wb_clk_i _01519_ _00120_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[109\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11324__S net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12706_ net1351 vssd1 vssd1 vccd1 vccd1 _00470_ sky130_fd_sc_hd__inv_2
XANTENNA__07495__B1 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08692__C1 net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10898_ _06488_ _06489_ _06490_ net586 vssd1 vssd1 vccd1 vccd1 _06491_ sky130_fd_sc_hd__o211a_4
XFILLER_0_127_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13686_ clknet_leaf_153_wb_clk_i _01450_ _00051_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[40\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_66_770 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12637_ net1382 vssd1 vssd1 vccd1 vccd1 _00401_ sky130_fd_sc_hd__inv_2
XANTENNA__08039__A2 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_152_wb_clk_i_A clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_12568_ net1379 vssd1 vssd1 vccd1 vccd1 _00332_ sky130_fd_sc_hd__inv_2
XFILLER_0_81_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_678 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08995__B1 net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_152_Right_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14307_ clknet_leaf_33_wb_clk_i _02071_ _00672_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[661\]
+ sky130_fd_sc_hd__dfrtp_1
X_11519_ _06632_ net2538 net390 vssd1 vssd1 vccd1 vccd1 _01987_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_117_2774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_2785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12499_ net1256 vssd1 vssd1 vccd1 vccd1 _00263_ sky130_fd_sc_hd__inv_2
Xhold207 _02632_ vssd1 vssd1 vccd1 vccd1 net1700 sky130_fd_sc_hd__dlygate4sd3_1
Xhold218 team_03_WB.instance_to_wrap.CPU_DAT_I\[17\] vssd1 vssd1 vccd1 vccd1 net1711
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold229 _02580_ vssd1 vssd1 vccd1 vccd1 net1722 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_169_3841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14238_ clknet_leaf_114_wb_clk_i _02002_ _00603_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[592\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11279__B net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_169_3852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11346__A2 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11994__S net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14169_ clknet_leaf_169_wb_clk_i _01933_ _00534_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[523\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07014__A3 net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10554__B1 net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08869__A _04770_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout709 net711 vssd1 vssd1 vccd1 vccd1 net709 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_0_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11897__A3 net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06991_ net1020 net826 _02825_ team_03_WB.instance_to_wrap.core.decoder.inst\[30\]
+ vssd1 vssd1 vccd1 vccd1 _02933_ sky130_fd_sc_hd__nor4b_1
XFILLER_0_147_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11295__A net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08730_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[804\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[772\]
+ net978 vssd1 vssd1 vccd1 vccd1 _04672_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1280 net1283 vssd1 vssd1 vccd1 vccd1 net1280 sky130_fd_sc_hd__buf_4
XANTENNA__09711__A2 net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1291 net1295 vssd1 vssd1 vccd1 vccd1 net1291 sky130_fd_sc_hd__buf_4
XFILLER_0_56_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08661_ net1056 team_03_WB.instance_to_wrap.core.register_file.registers_state\[455\]
+ net1009 team_03_WB.instance_to_wrap.core.register_file.registers_state\[487\] net1078
+ vssd1 vssd1 vccd1 vccd1 _04603_ sky130_fd_sc_hd__a221o_1
X_07612_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[793\] net802
+ _03548_ net1121 vssd1 vssd1 vccd1 vccd1 _03554_ sky130_fd_sc_hd__o211a_1
X_08592_ _04505_ _04533_ net547 vssd1 vssd1 vccd1 vccd1 _04534_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07543_ net1137 _03483_ net1166 vssd1 vssd1 vccd1 vccd1 _03485_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_89_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07370__A1_N net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_163_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09475__A1 net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_191_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_159_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_400 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07486__A0 _03425_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11282__A1 net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07474_ _03411_ _03415_ net1147 vssd1 vssd1 vccd1 vccd1 _03416_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_5_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_158_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11821__A3 net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09213_ _03429_ _04032_ net431 _05146_ vssd1 vssd1 vccd1 vccd1 _05155_ sky130_fd_sc_hd__or4_1
XANTENNA__07013__A net1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_174_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout326_A _06811_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09144_ net543 _04179_ _05085_ vssd1 vssd1 vccd1 vccd1 _05086_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout1068_A net1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11034__B2 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07948__A net1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08770__C _04711_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14842__Q net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08986__B1 net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09075_ net941 _05015_ _05016_ vssd1 vssd1 vccd1 vccd1 _05017_ sky130_fd_sc_hd__o21a_1
XANTENNA__12065__S net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1235_A net1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08026_ net1177 team_03_WB.instance_to_wrap.core.register_file.registers_state\[81\]
+ net764 team_03_WB.instance_to_wrap.core.register_file.registers_state\[113\] net727
+ vssd1 vssd1 vccd1 vccd1 _03968_ sky130_fd_sc_hd__o221a_1
XFILLER_0_60_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold730 team_03_WB.instance_to_wrap.core.register_file.registers_state\[523\] vssd1
+ vssd1 vccd1 vccd1 net2223 sky130_fd_sc_hd__dlygate4sd3_1
Xhold741 team_03_WB.instance_to_wrap.core.register_file.registers_state\[761\] vssd1
+ vssd1 vccd1 vccd1 net2234 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout695_A net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold752 team_03_WB.instance_to_wrap.core.register_file.registers_state\[742\] vssd1
+ vssd1 vccd1 vccd1 net2245 sky130_fd_sc_hd__dlygate4sd3_1
Xhold763 team_03_WB.instance_to_wrap.core.register_file.registers_state\[235\] vssd1
+ vssd1 vccd1 vccd1 net2256 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold774 team_03_WB.instance_to_wrap.core.register_file.registers_state\[811\] vssd1
+ vssd1 vccd1 vccd1 net2267 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1023_X net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold785 team_03_WB.instance_to_wrap.core.register_file.registers_state\[893\] vssd1
+ vssd1 vccd1 vccd1 net2278 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1402_A net1408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11888__A3 net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold796 team_03_WB.instance_to_wrap.core.register_file.registers_state\[230\] vssd1
+ vssd1 vccd1 vccd1 net2289 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07683__A net1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09977_ net593 net1731 net292 vssd1 vssd1 vccd1 vccd1 _02736_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout483_X net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout862_A net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07961__A1 net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11409__S net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08928_ net862 _04868_ _04869_ vssd1 vssd1 vccd1 vccd1 _04870_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout650_X net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08859_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[928\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[896\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[800\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[768\]
+ net989 net1078 vssd1 vssd1 vccd1 vccd1 _04801_ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout748_X net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_58_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_58_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_11870_ _06536_ net2284 net377 vssd1 vssd1 vccd1 vccd1 _01670_ sky130_fd_sc_hd__mux2_1
X_10821_ _06423_ _06425_ net585 vssd1 vssd1 vccd1 vccd1 _06426_ sky130_fd_sc_hd__o21a_2
XFILLER_0_95_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout915_X net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_400 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10752_ team_03_WB.instance_to_wrap.core.pc.current_pc\[6\] net604 vssd1 vssd1 vccd1
+ vccd1 _06369_ sky130_fd_sc_hd__or2_1
X_13540_ net1320 vssd1 vssd1 vccd1 vccd1 _01304_ sky130_fd_sc_hd__inv_2
XANTENNA__10076__A2 net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07477__B1 net1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11371__C net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08674__C1 net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13471_ net1323 vssd1 vssd1 vccd1 vccd1 _01235_ sky130_fd_sc_hd__inv_2
XFILLER_0_137_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_168_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10683_ _06321_ net522 _06324_ net527 net1587 vssd1 vssd1 vccd1 vccd1 _02465_ sky130_fd_sc_hd__a32o_1
XANTENNA__10836__X _06438_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_239 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12422_ net1336 vssd1 vssd1 vccd1 vccd1 _00186_ sky130_fd_sc_hd__inv_2
XFILLER_0_153_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_1136 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_464 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input89_A wbs_adr_i[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_2368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12353_ net1262 vssd1 vssd1 vccd1 vccd1 _00117_ sky130_fd_sc_hd__inv_2
XFILLER_0_164_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_592 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_1910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11304_ _06614_ net2759 net407 vssd1 vssd1 vccd1 vccd1 _02141_ sky130_fd_sc_hd__mux2_1
X_15072_ net1458 vssd1 vssd1 vccd1 vccd1 la_data_out[8] sky130_fd_sc_hd__buf_2
XFILLER_0_133_694 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12284_ net1411 vssd1 vssd1 vccd1 vccd1 _00048_ sky130_fd_sc_hd__inv_2
XANTENNA__11099__B net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_1921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14023_ clknet_leaf_113_wb_clk_i _01787_ _00388_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[377\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_147_3402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11235_ _06405_ net709 net827 vssd1 vssd1 vccd1 vccd1 _06685_ sky130_fd_sc_hd__and3_1
XFILLER_0_31_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_112_2671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10536__B1 net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11879__A3 net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_2682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_71_1829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11166_ net2440 net414 _06661_ net508 vssd1 vssd1 vccd1 vccd1 _02223_ sky130_fd_sc_hd__a22o_1
XFILLER_0_101_1011 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_1071 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11319__S net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07952__A1 net1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10117_ _05954_ _05955_ _03065_ vssd1 vssd1 vccd1 vccd1 _05960_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_140_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11097_ net835 net298 vssd1 vssd1 vccd1 vccd1 _06625_ sky130_fd_sc_hd__and2_2
XFILLER_0_172_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10048_ net8 net1036 net910 net1849 vssd1 vssd1 vccd1 vccd1 _02683_ sky130_fd_sc_hd__o22a_1
X_14925_ clknet_leaf_44_wb_clk_i _02680_ _01290_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_O\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_160_3657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_3_4_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_160_3668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12939__A net1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07704__A1 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold90 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1017\] vssd1
+ vssd1 vccd1 vccd1 net1583 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08901__B1 net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14856_ clknet_leaf_64_wb_clk_i net1813 _01221_ vssd1 vssd1 vccd1 vccd1 net111 sky130_fd_sc_hd__dfrtp_1
XANTENNA__09313__A net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14927__Q team_03_WB.instance_to_wrap.CPU_DAT_O\[14\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_13807_ clknet_leaf_134_wb_clk_i _01571_ _00172_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[161\]
+ sky130_fd_sc_hd__dfrtp_1
X_14787_ clknet_leaf_102_wb_clk_i _02551_ _01152_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_I\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_147_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11999_ net295 net2390 net444 vssd1 vssd1 vccd1 vccd1 _01545_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_11_Left_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07468__B1 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11264__A1 net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11281__C net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13738_ clknet_leaf_0_wb_clk_i _01502_ _00103_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[92\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09967__B net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_2814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_119_2825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13669_ clknet_leaf_14_wb_clk_i _01433_ _00034_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_143_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11016__A1 net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_848 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07190_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[819\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[787\]
+ net762 vssd1 vssd1 vccd1 vccd1 _03132_ sky130_fd_sc_hd__mux2_1
XANTENNA__08417__C1 net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08968__B1 net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07487__B _03428_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_968 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_151_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09900_ _05834_ _05841_ vssd1 vssd1 vccd1 vccd1 _05842_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_20_Left_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10527__B1 net1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout506 net517 vssd1 vssd1 vccd1 vccd1 net506 sky130_fd_sc_hd__buf_2
XFILLER_0_10_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09831_ net579 _04711_ net667 _05772_ vssd1 vssd1 vccd1 vccd1 _05773_ sky130_fd_sc_hd__a22o_1
Xfanout517 _06448_ vssd1 vssd1 vccd1 vccd1 net517 sky130_fd_sc_hd__clkbuf_8
Xfanout528 _06309_ vssd1 vssd1 vccd1 vccd1 net528 sky130_fd_sc_hd__clkbuf_4
Xfanout539 net540 vssd1 vssd1 vccd1 vccd1 net539 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07943__A1 net1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08291__S1 net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11229__S net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09762_ _04327_ _05073_ _05702_ _05703_ vssd1 vssd1 vccd1 vccd1 _05704_ sky130_fd_sc_hd__a211o_1
X_06974_ net1205 team_03_WB.instance_to_wrap.core.register_file.registers_state\[645\]
+ net787 team_03_WB.instance_to_wrap.core.register_file.registers_state\[677\] net753
+ vssd1 vssd1 vccd1 vccd1 _02916_ sky130_fd_sc_hd__o221a_1
XANTENNA__09145__B1 net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08713_ net1059 team_03_WB.instance_to_wrap.core.register_file.registers_state\[68\]
+ net1013 team_03_WB.instance_to_wrap.core.register_file.registers_state\[100\] net944
+ vssd1 vssd1 vccd1 vccd1 _04655_ sky130_fd_sc_hd__a221o_1
X_09693_ _05276_ _05279_ _05198_ _05207_ vssd1 vssd1 vccd1 vccd1 _05635_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_174_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout276_A _06434_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08644_ net927 _04584_ _04585_ vssd1 vssd1 vccd1 vccd1 _04586_ sky130_fd_sc_hd__a21o_1
XFILLER_0_174_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06847__A net1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09223__A _04503_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08575_ net1220 _04515_ _04516_ vssd1 vssd1 vccd1 vccd1 _04517_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout443_A net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1185_A net1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07526_ net1102 team_03_WB.instance_to_wrap.core.register_file.registers_state\[710\]
+ net799 team_03_WB.instance_to_wrap.core.register_file.registers_state\[742\] net732
+ vssd1 vssd1 vccd1 vccd1 _03468_ sky130_fd_sc_hd__a221o_1
XFILLER_0_49_567 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_824 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_910 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_915 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07457_ net1184 team_03_WB.instance_to_wrap.core.register_file.registers_state\[213\]
+ vssd1 vssd1 vccd1 vccd1 _03399_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout610_A net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_712 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1352_A net1358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout329_X net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_174_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11007__B2 net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_176_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_176_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_07388_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[287\] net791
+ vssd1 vssd1 vccd1 vccd1 _03330_ sky130_fd_sc_hd__or2_1
XFILLER_0_17_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11558__A2 net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09127_ net588 vssd1 vssd1 vccd1 vccd1 _05069_ sky130_fd_sc_hd__inv_2
XANTENNA__09081__C1 net1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1140_X net1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_105_wb_clk_i clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_105_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__10766__B1 net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1238_X net1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09058_ net1047 team_03_WB.instance_to_wrap.core.register_file.registers_state\[591\]
+ net998 team_03_WB.instance_to_wrap.core.register_file.registers_state\[623\] net949
+ vssd1 vssd1 vccd1 vccd1 _05000_ sky130_fd_sc_hd__a221o_1
XFILLER_0_114_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout698_X net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08009_ net1178 team_03_WB.instance_to_wrap.core.register_file.registers_state\[849\]
+ vssd1 vssd1 vccd1 vccd1 _03951_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_92_2265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_2276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold560 team_03_WB.instance_to_wrap.core.register_file.registers_state\[896\] vssd1
+ vssd1 vccd1 vccd1 net2053 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10518__B1 net1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold571 team_03_WB.instance_to_wrap.core.register_file.registers_state\[462\] vssd1
+ vssd1 vccd1 vccd1 net2064 sky130_fd_sc_hd__dlygate4sd3_1
Xhold582 team_03_WB.instance_to_wrap.core.register_file.registers_state\[275\] vssd1
+ vssd1 vccd1 vccd1 net2075 sky130_fd_sc_hd__dlygate4sd3_1
X_11020_ net624 _06583_ vssd1 vssd1 vccd1 vccd1 _06584_ sky130_fd_sc_hd__nor2_1
Xhold593 team_03_WB.instance_to_wrap.core.register_file.registers_state\[628\] vssd1
+ vssd1 vccd1 vccd1 net2086 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08302__A net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout865_X net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_10__f_wb_clk_i_A clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07934__A1 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12971_ net1283 vssd1 vssd1 vccd1 vccd1 _00735_ sky130_fd_sc_hd__inv_2
XANTENNA__07147__C1 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1260 team_03_WB.instance_to_wrap.core.pc.current_pc\[0\] vssd1 vssd1 vccd1 vccd1
+ net2753 sky130_fd_sc_hd__dlygate4sd3_1
X_14710_ clknet_leaf_31_wb_clk_i _02474_ _01075_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.decoder.inst\[7\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1271 team_03_WB.instance_to_wrap.core.register_file.registers_state\[348\] vssd1
+ vssd1 vccd1 vccd1 net2764 sky130_fd_sc_hd__dlygate4sd3_1
X_11922_ _06621_ net2558 net367 vssd1 vssd1 vccd1 vccd1 _01620_ sky130_fd_sc_hd__mux2_1
Xhold1282 team_03_WB.instance_to_wrap.core.register_file.registers_state\[193\] vssd1
+ vssd1 vccd1 vccd1 net2775 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08895__C1 net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09133__A _02804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14641_ clknet_leaf_140_wb_clk_i _02405_ _01006_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[995\]
+ sky130_fd_sc_hd__dfstp_1
X_11853_ net275 net2070 net376 vssd1 vssd1 vccd1 vccd1 _01687_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_68_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10804_ net687 _05563_ _06401_ vssd1 vssd1 vccd1 vccd1 _06412_ sky130_fd_sc_hd__a21o_1
XFILLER_0_32_1112 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11246__A1 net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11784_ net2412 _06617_ net328 vssd1 vssd1 vccd1 vccd1 _01754_ sky130_fd_sc_hd__mux2_1
X_14572_ clknet_leaf_14_wb_clk_i _02336_ _00937_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[926\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_99_2408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_2419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13523_ net1306 vssd1 vssd1 vccd1 vccd1 _01287_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_64_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10735_ net1658 net529 net524 _06359_ vssd1 vssd1 vccd1 vccd1 _02448_ sky130_fd_sc_hd__a22o_1
XFILLER_0_153_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12494__A net1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11602__S net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_153_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_136_3158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_3169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07588__A net1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13454_ net1345 vssd1 vssd1 vccd1 vccd1 _01218_ sky130_fd_sc_hd__inv_2
X_10666_ net1145 _06307_ _06302_ team_03_WB.instance_to_wrap.core.ru.state\[3\] vssd1
+ vssd1 vccd1 vccd1 _06308_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__07870__B1 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_153_767 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10206__C1 _02994_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11549__A2 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06923__C net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12405_ net1271 vssd1 vssd1 vccd1 vccd1 _00169_ sky130_fd_sc_hd__inv_2
XANTENNA__10757__A0 team_03_WB.instance_to_wrap.core.pc.current_pc\[4\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13385_ net1415 vssd1 vssd1 vccd1 vccd1 _01149_ sky130_fd_sc_hd__inv_2
X_10597_ net1142 team_03_WB.instance_to_wrap.core.d_hit team_03_WB.instance_to_wrap.core.ru.state\[5\]
+ _06281_ net840 vssd1 vssd1 vccd1 vccd1 _02531_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_114_2711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_220 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_114_2722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_11_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15124_ net1489 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[29] sky130_fd_sc_hd__buf_2
Xoutput109 net109 vssd1 vssd1 vccd1 vccd1 ADR_O[15] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_50_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12336_ net1410 vssd1 vssd1 vccd1 vccd1 _00100_ sky130_fd_sc_hd__inv_2
XFILLER_0_121_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06976__A2 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11397__X _06751_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15055_ net1441 vssd1 vssd1 vccd1 vccd1 gpio_out[1] sky130_fd_sc_hd__buf_2
XFILLER_0_10_128 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12267_ net1291 vssd1 vssd1 vccd1 vccd1 _00031_ sky130_fd_sc_hd__inv_2
XANTENNA__10509__B1 net1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14006_ clknet_leaf_178_wb_clk_i _01770_ _00371_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[360\]
+ sky130_fd_sc_hd__dfrtp_1
X_11218_ _06495_ net2655 net488 vssd1 vssd1 vccd1 vccd1 _02191_ sky130_fd_sc_hd__mux2_1
XANTENNA__09308__A _04565_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12198_ net1497 vssd1 vssd1 vccd1 vccd1 _02355_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_162_3708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07925__A1 net1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11149_ net493 net647 _06651_ net412 net1930 vssd1 vssd1 vccd1 vccd1 _02230_ sky130_fd_sc_hd__a32o_1
XANTENNA__08866__B _04807_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14908_ clknet_leaf_54_wb_clk_i _00002_ _01273_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.ru.state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07689__B1 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11485__B2 net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08350__A1 net1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14839_ clknet_leaf_83_wb_clk_i _02603_ _01204_ vssd1 vssd1 vccd1 vccd1 net103 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10189__A _03460_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1078 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12029__A3 net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_651 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08360_ net855 _04300_ _04301_ vssd1 vssd1 vccd1 vccd1 _04302_ sky130_fd_sc_hd__or3_1
XANTENNA__08638__C1 net1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08882__A _04080_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07311_ net1185 team_03_WB.instance_to_wrap.core.register_file.registers_state\[861\]
+ net768 team_03_WB.instance_to_wrap.core.register_file.registers_state\[893\] net1162
+ vssd1 vssd1 vccd1 vccd1 _03253_ sky130_fd_sc_hd__o221a_1
Xclkbuf_leaf_3_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_3_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__09697__B net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08291_ _04229_ _04230_ _04231_ _04232_ net861 net937 vssd1 vssd1 vccd1 vccd1 _04233_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__07310__C1 net1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11512__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07242_ net1191 team_03_WB.instance_to_wrap.core.register_file.registers_state\[712\]
+ vssd1 vssd1 vccd1 vccd1 _03184_ sky130_fd_sc_hd__or2_1
XANTENNA__10460__A2 _05945_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07861__B1 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07173_ net806 _03113_ _03114_ vssd1 vssd1 vccd1 vccd1 _03115_ sky130_fd_sc_hd__or3_1
XANTENNA__10748__B1 net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_6__f_wb_clk_i_A clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_143_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07010__B net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07613__B1 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout303 _05945_ vssd1 vssd1 vccd1 vccd1 net303 sky130_fd_sc_hd__buf_4
Xfanout314 _05387_ vssd1 vssd1 vccd1 vccd1 net314 sky130_fd_sc_hd__buf_2
XANTENNA__07664__C net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout325 _06811_ vssd1 vssd1 vccd1 vccd1 net325 sky130_fd_sc_hd__clkbuf_8
XANTENNA__07916__A1 net1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout393_A net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout336 net337 vssd1 vssd1 vccd1 vccd1 net336 sky130_fd_sc_hd__buf_6
X_09814_ _05754_ _05755_ _05752_ vssd1 vssd1 vccd1 vccd1 _05756_ sky130_fd_sc_hd__or3b_1
Xfanout347 _06804_ vssd1 vssd1 vccd1 vccd1 net347 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11186__C net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout358 _06818_ vssd1 vssd1 vccd1 vccd1 net358 sky130_fd_sc_hd__buf_4
XANTENNA_fanout1100_A net1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout369 _06814_ vssd1 vssd1 vccd1 vccd1 net369 sky130_fd_sc_hd__buf_6
XANTENNA__10090__C _05659_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09745_ _05213_ _05235_ _05275_ vssd1 vssd1 vccd1 vccd1 _05687_ sky130_fd_sc_hd__nand3_1
XANTENNA_fanout560_A _03063_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09669__A1 net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06957_ net814 _02897_ _02898_ vssd1 vssd1 vccd1 vccd1 _02899_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout658_A net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout279_X net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09676_ _03391_ _04119_ net539 vssd1 vssd1 vccd1 vccd1 _05618_ sky130_fd_sc_hd__o21ai_1
X_06888_ _02822_ _02823_ _02827_ _02829_ vssd1 vssd1 vccd1 vccd1 _02830_ sky130_fd_sc_hd__or4_2
XANTENNA__11476__B2 net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08341__A1 net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08627_ net1240 team_03_WB.instance_to_wrap.core.register_file.registers_state\[134\]
+ net983 team_03_WB.instance_to_wrap.core.register_file.registers_state\[166\] net941
+ vssd1 vssd1 vccd1 vccd1 _04569_ sky130_fd_sc_hd__o221a_1
XFILLER_0_96_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_139_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1090_X net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout446_X net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1188_X net1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08629__C1 net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08558_ _04498_ _04499_ net1219 vssd1 vssd1 vccd1 vccd1 _04500_ sky130_fd_sc_hd__o21a_1
XFILLER_0_65_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07509_ net1110 team_03_WB.instance_to_wrap.core.register_file.registers_state\[327\]
+ net803 team_03_WB.instance_to_wrap.core.register_file.registers_state\[359\] net1158
+ vssd1 vssd1 vccd1 vccd1 _03451_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_147_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout613_X net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08489_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[59\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[27\]
+ net987 vssd1 vssd1 vccd1 vccd1 _04431_ sky130_fd_sc_hd__mux2_1
XANTENNA__09841__A1 _02992_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11422__S net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13203__A net1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10520_ net146 net1034 net1026 net1656 vssd1 vssd1 vccd1 vccd1 _02590_ sky130_fd_sc_hd__a22o_1
XFILLER_0_174_380 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09400__B _04475_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07852__B1 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_570 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_2305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10451_ _06135_ _06266_ vssd1 vssd1 vccd1 vccd1 _06267_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_94_2316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10739__B1 net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13170_ net1397 vssd1 vssd1 vccd1 vccd1 _00934_ sky130_fd_sc_hd__inv_2
XANTENNA__07604__B1 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10382_ team_03_WB.instance_to_wrap.core.pc.current_pc\[18\] _06144_ vssd1 vssd1
+ vccd1 vccd1 _06211_ sky130_fd_sc_hd__xor2_1
XFILLER_0_150_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_131_3066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08801__C1 net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout982_X net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12121_ net1563 vssd1 vssd1 vccd1 vccd1 _02432_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__07080__A1 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_995 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12052_ _06454_ net2559 net355 vssd1 vssd1 vccd1 vccd1 _01494_ sky130_fd_sc_hd__mux2_1
Xhold390 net196 vssd1 vssd1 vccd1 vccd1 net1883 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11377__B net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07368__C1 net1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11003_ net276 net650 net704 net828 vssd1 vssd1 vccd1 vccd1 _06574_ sky130_fd_sc_hd__and4_1
XANTENNA__11703__A2 net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_73_wb_clk_i clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_73_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08580__A1 net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout870 _04082_ vssd1 vssd1 vccd1 vccd1 net870 sky130_fd_sc_hd__buf_4
XANTENNA__09109__B1 net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout881 net882 vssd1 vssd1 vccd1 vccd1 net881 sky130_fd_sc_hd__clkbuf_4
Xfanout892 net893 vssd1 vssd1 vccd1 vccd1 net892 sky130_fd_sc_hd__buf_2
XFILLER_0_99_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11393__A net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12954_ net1378 vssd1 vssd1 vccd1 vccd1 _00718_ sky130_fd_sc_hd__inv_2
XANTENNA__11467__B2 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_2570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1090 team_03_WB.instance_to_wrap.core.register_file.registers_state\[95\] vssd1
+ vssd1 vccd1 vccd1 net2583 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_158_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_107_2581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11905_ net633 _06714_ net467 net373 net2097 vssd1 vssd1 vccd1 vccd1 _01636_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_66_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_139 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_303 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12885_ net1273 vssd1 vssd1 vccd1 vccd1 _00649_ sky130_fd_sc_hd__inv_2
XFILLER_0_68_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_3209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14624_ clknet_leaf_192_wb_clk_i _02388_ _00989_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[978\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_114_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11836_ net657 _06674_ net478 net326 net1882 vssd1 vssd1 vccd1 vccd1 _01703_ sky130_fd_sc_hd__a32o_1
XFILLER_0_56_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_2489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08096__B1 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14555_ clknet_leaf_121_wb_clk_i _02319_ _00920_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[909\]
+ sky130_fd_sc_hd__dfrtp_1
X_11767_ _06599_ net464 net331 net2336 vssd1 vssd1 vccd1 vccd1 _01770_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_155_3556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_155_3567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13506_ net1321 vssd1 vssd1 vccd1 vccd1 _01270_ sky130_fd_sc_hd__inv_2
XANTENNA__10442__A2 _05945_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10718_ team_03_WB.instance_to_wrap.core.pc.current_pc\[21\] net602 vssd1 vssd1 vccd1
+ vccd1 _06350_ sky130_fd_sc_hd__or2_1
X_14486_ clknet_leaf_152_wb_clk_i _02250_ _00851_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[840\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08207__A net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11698_ _06740_ net379 net338 net2069 vssd1 vssd1 vccd1 vccd1 _01836_ sky130_fd_sc_hd__a22o_1
XANTENNA__07111__A net1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13437_ net1424 vssd1 vssd1 vccd1 vccd1 _01201_ sky130_fd_sc_hd__inv_2
X_10649_ team_03_WB.instance_to_wrap.core.decoder.inst\[12\] team_03_WB.instance_to_wrap.CPU_DAT_O\[12\]
+ net846 vssd1 vssd1 vccd1 vccd1 _02479_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12952__A net1380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08399__A1 net1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_299 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13368_ net1319 vssd1 vssd1 vccd1 vccd1 _01132_ sky130_fd_sc_hd__inv_2
XFILLER_0_51_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_415 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06949__A2 _02888_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15107_ net912 vssd1 vssd1 vccd1 vccd1 net242 sky130_fd_sc_hd__clkbuf_1
XANTENNA__07071__A1 net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12319_ net1285 vssd1 vssd1 vccd1 vccd1 _00083_ sky130_fd_sc_hd__inv_2
XFILLER_0_107_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13299_ net1327 vssd1 vssd1 vccd1 vccd1 _01063_ sky130_fd_sc_hd__inv_2
X_15038_ clknet_leaf_91_wb_clk_i _02758_ _01403_ vssd1 vssd1 vccd1 vccd1 net194 sky130_fd_sc_hd__dfrtp_1
XANTENNA__11287__B net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10191__B net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09899__A1 net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07359__C1 net1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07860_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[539\] net783
+ net751 _03801_ vssd1 vssd1 vccd1 vccd1 _03802_ sky130_fd_sc_hd__a211o_1
XANTENNA__08571__A1 net1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07791_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[555\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[523\]
+ net775 vssd1 vssd1 vccd1 vccd1 _03733_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_127_2979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11507__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09530_ net580 _05471_ net351 vssd1 vssd1 vccd1 vccd1 _05472_ sky130_fd_sc_hd__o21a_1
XFILLER_0_64_64 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07126__A2 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08323__A1 net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09461_ _05399_ _05402_ net570 vssd1 vssd1 vccd1 vccd1 _05403_ sky130_fd_sc_hd__mux2_1
XANTENNA__09204__C _05144_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08412_ net853 _04340_ _04353_ vssd1 vssd1 vccd1 vccd1 _04354_ sky130_fd_sc_hd__o21ba_4
X_09392_ _04382_ _05312_ _05319_ vssd1 vssd1 vccd1 vccd1 _05334_ sky130_fd_sc_hd__or3_1
XFILLER_0_4_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08343_ net1238 team_03_WB.instance_to_wrap.core.register_file.registers_state\[213\]
+ net968 team_03_WB.instance_to_wrap.core.register_file.registers_state\[245\] net938
+ vssd1 vssd1 vccd1 vccd1 _04285_ sky130_fd_sc_hd__o221a_1
XFILLER_0_4_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_183 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_15_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07834__B1 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08274_ net1234 team_03_WB.instance_to_wrap.core.register_file.registers_state\[215\]
+ net963 team_03_WB.instance_to_wrap.core.register_file.registers_state\[247\] net937
+ vssd1 vssd1 vccd1 vccd1 _04216_ sky130_fd_sc_hd__o221a_1
XFILLER_0_104_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_156_391 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07225_ net1138 _03162_ _03164_ _03166_ net721 vssd1 vssd1 vccd1 vccd1 _03167_ sky130_fd_sc_hd__o41a_1
XFILLER_0_61_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15011__Q team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[30\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout406_A _06717_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1050_A net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10085__C net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1148_A team_03_WB.instance_to_wrap.core.decoder.inst\[23\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07156_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[384\] net785
+ _03097_ vssd1 vssd1 vccd1 vccd1 _03098_ sky130_fd_sc_hd__a21o_1
XFILLER_0_89_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10197__A1 team_03_WB.instance_to_wrap.core.pc.current_pc\[4\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_258 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11394__B1 net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07062__A1 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07087_ net1102 team_03_WB.instance_to_wrap.core.register_file.registers_state\[673\]
+ net899 vssd1 vssd1 vccd1 vccd1 _03029_ sky130_fd_sc_hd__or3_1
XFILLER_0_112_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1315_A net1330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_160_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout775_A net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout396_X net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1109 net1111 vssd1 vssd1 vccd1 vccd1 net1109 sky130_fd_sc_hd__buf_2
XFILLER_0_10_492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07365__A2 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout942_A net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_29_Right_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07989_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[816\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[784\]
+ net782 vssd1 vssd1 vccd1 vccd1 _03931_ sky130_fd_sc_hd__mux2_1
XANTENNA__07770__C1 net1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11417__S net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09728_ _04210_ _05014_ _05071_ _04895_ net558 net571 vssd1 vssd1 vccd1 vccd1 _05670_
+ sky130_fd_sc_hd__mux4_2
XTAP_TAPCELL_ROW_87_2164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11449__B2 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08314__A1 net1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09659_ _05084_ _05089_ _05091_ _05098_ net563 net560 vssd1 vssd1 vccd1 vccd1 _05601_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_26_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout730_X net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout828_X net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11941__A net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_166_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_191_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_191_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_38_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12670_ net1387 vssd1 vssd1 vccd1 vccd1 _00434_ sky130_fd_sc_hd__inv_2
XFILLER_0_166_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_139_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11621_ _06695_ net381 net347 net2489 vssd1 vssd1 vccd1 vccd1 _01911_ sky130_fd_sc_hd__a22o_1
XFILLER_0_166_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_61_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_120_wb_clk_i clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_120_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_61_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_120 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14340_ clknet_leaf_36_wb_clk_i _02104_ _00705_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[694\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_147_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_133_3106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11552_ net655 _06662_ vssd1 vssd1 vccd1 vccd1 _06791_ sky130_fd_sc_hd__nor2_1
XFILLER_0_107_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08027__A net1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_38_Right_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10503_ net128 net1033 net907 net1679 vssd1 vssd1 vccd1 vccd1 _02606_ sky130_fd_sc_hd__a22o_1
XFILLER_0_150_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11483_ net505 net633 _06606_ net393 net2152 vssd1 vssd1 vccd1 vccd1 _02020_ sky130_fd_sc_hd__a32o_1
XFILLER_0_52_348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14271_ clknet_leaf_171_wb_clk_i _02035_ _00636_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[625\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_163_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_150_3453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10434_ net285 _06138_ _06250_ net682 vssd1 vssd1 vccd1 vccd1 _06254_ sky130_fd_sc_hd__o31a_1
XANTENNA_input71_A wbs_adr_i[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07866__A net1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13222_ net1301 vssd1 vssd1 vccd1 vccd1 _00986_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_150_3464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire589 _05012_ vssd1 vssd1 vccd1 vccd1 net589 sky130_fd_sc_hd__buf_4
XFILLER_0_33_584 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_223 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10365_ team_03_WB.instance_to_wrap.core.pc.current_pc\[20\] _06145_ team_03_WB.instance_to_wrap.core.pc.current_pc\[21\]
+ vssd1 vssd1 vccd1 vccd1 _06197_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07585__B net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13153_ net1261 vssd1 vssd1 vccd1 vccd1 _00917_ sky130_fd_sc_hd__inv_2
XFILLER_0_104_984 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_59_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_5__f_wb_clk_i_X clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_12104_ _06798_ net470 net441 net2063 vssd1 vssd1 vccd1 vccd1 _01443_ sky130_fd_sc_hd__a22o_1
X_13084_ net1419 vssd1 vssd1 vccd1 vccd1 _00848_ sky130_fd_sc_hd__inv_2
X_10296_ team_03_WB.instance_to_wrap.core.pc.current_pc\[9\] team_03_WB.instance_to_wrap.core.pc.current_pc\[8\]
+ _06136_ vssd1 vssd1 vccd1 vccd1 _06138_ sky130_fd_sc_hd__and3_1
X_12035_ net639 _06604_ net473 net362 net2291 vssd1 vssd1 vccd1 vccd1 _01510_ sky130_fd_sc_hd__a32o_1
XFILLER_0_100_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_69_wb_clk_i_A clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_2610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_47_Right_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_109_2621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06929__B net1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11327__S net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09305__B _05144_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_2529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13986_ clknet_leaf_175_wb_clk_i _01750_ _00351_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[340\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08305__A1 net1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12101__A2 _06675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07106__A net1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10112__A1 _04807_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12937_ net1259 vssd1 vssd1 vccd1 vccd1 _00701_ sky130_fd_sc_hd__inv_2
XFILLER_0_73_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_157_3607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_2876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_122_2887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12868_ net1382 vssd1 vssd1 vccd1 vccd1 _00632_ sky130_fd_sc_hd__inv_2
XFILLER_0_69_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_312 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14607_ clknet_leaf_135_wb_clk_i _02371_ _00972_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[961\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11570__B net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08069__B1 net1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_174_3943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11819_ _06649_ net459 net324 net1904 vssd1 vssd1 vccd1 vccd1 _01720_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_174_3954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_174_3965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12799_ net1349 vssd1 vssd1 vccd1 vccd1 _00563_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_56_Right_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_174_3976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_520 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_840 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14538_ clknet_leaf_7_wb_clk_i _02302_ _00903_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[892\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_996 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11997__S net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10966__A3 net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10820__C1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07292__A1 net1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09018__C1 net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14469_ clknet_leaf_37_wb_clk_i _02233_ _00834_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[823\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06951__Y _02893_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07010_ net1020 net582 vssd1 vssd1 vccd1 vccd1 _02952_ sky130_fd_sc_hd__nor2_1
XANTENNA__09569__B1 net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_759 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08371__S net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11376__B1 net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08792__A1 net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08961_ net1245 team_03_WB.instance_to_wrap.core.register_file.registers_state\[329\]
+ net986 team_03_WB.instance_to_wrap.core.register_file.registers_state\[361\] net1079
+ vssd1 vssd1 vccd1 vccd1 _04903_ sky130_fd_sc_hd__o221a_1
XFILLER_0_80_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_65_Right_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11448__D _06558_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07912_ net1178 team_03_WB.instance_to_wrap.core.register_file.registers_state\[879\]
+ net878 _03853_ vssd1 vssd1 vccd1 vccd1 _03854_ sky130_fd_sc_hd__a31o_1
X_08892_ net578 net351 vssd1 vssd1 vccd1 vccd1 _04834_ sky130_fd_sc_hd__nand2_1
X_07843_ _03783_ _03784_ vssd1 vssd1 vccd1 vccd1 _03785_ sky130_fd_sc_hd__and2_1
XFILLER_0_75_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07774_ net1098 net897 team_03_WB.instance_to_wrap.core.register_file.registers_state\[524\]
+ vssd1 vssd1 vccd1 vccd1 _03716_ sky130_fd_sc_hd__o21a_1
XANTENNA__09930__S net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_3_Left_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09513_ _05435_ _05453_ vssd1 vssd1 vccd1 vccd1 _05455_ sky130_fd_sc_hd__or2_1
XFILLER_0_79_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15006__Q team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[25\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout356_A _06818_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1098_A net1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09444_ _05371_ _05385_ _05370_ vssd1 vssd1 vccd1 vccd1 _05386_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_82_2061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_166_Right_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_74_Right_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09231__A _03314_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09375_ _05160_ _05316_ vssd1 vssd1 vccd1 vccd1 _05317_ sky130_fd_sc_hd__nand2b_1
XANTENNA__12068__S net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout523_A _06322_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1265_A net1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_451 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08326_ net432 net424 _04267_ net541 vssd1 vssd1 vccd1 vccd1 _04268_ sky130_fd_sc_hd__o31a_1
XANTENNA__07807__B1 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10096__B _05429_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_151_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08257_ net934 _04197_ _04198_ net854 vssd1 vssd1 vccd1 vccd1 _04199_ sky130_fd_sc_hd__o211a_1
XFILLER_0_46_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout311_X net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09885__B _04148_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_966 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08480__B1 net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1053_X net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout409_X net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07208_ net1114 _03147_ _03148_ vssd1 vssd1 vccd1 vccd1 _03150_ sky130_fd_sc_hd__or3_1
XFILLER_0_171_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08188_ net1231 team_03_WB.instance_to_wrap.core.register_file.registers_state\[467\]
+ net957 team_03_WB.instance_to_wrap.core.register_file.registers_state\[499\] net1211
+ vssd1 vssd1 vccd1 vccd1 _04130_ sky130_fd_sc_hd__o221a_1
XANTENNA__08281__S net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout892_A net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_595 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07139_ _03077_ _03080_ net819 vssd1 vssd1 vccd1 vccd1 _03081_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout1220_X net1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_103_wb_clk_i_A clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09980__A0 _03103_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11001__A net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_83_Right_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10150_ _03139_ _05990_ vssd1 vssd1 vccd1 vccd1 _05992_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_37_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout680_X net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout778_X net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_2204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10081_ _05918_ _05923_ _05924_ _02831_ vssd1 vssd1 vccd1 vccd1 _05925_ sky130_fd_sc_hd__a211o_4
XTAP_TAPCELL_ROW_54_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09732__B1 net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout945_X net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13840_ clknet_leaf_158_wb_clk_i _01604_ _00205_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[194\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12095__A1 net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13771_ clknet_leaf_41_wb_clk_i _01535_ _00136_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[125\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_234 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08299__B1 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10983_ net1251 net833 vssd1 vssd1 vccd1 vccd1 _06561_ sky130_fd_sc_hd__nor2_2
XPHY_EDGE_ROW_92_Right_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_139_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12722_ net1396 vssd1 vssd1 vccd1 vccd1 _00486_ sky130_fd_sc_hd__inv_2
XFILLER_0_69_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09141__A net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_2426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_133_Right_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06944__S1 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_2437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12653_ net1311 vssd1 vssd1 vccd1 vccd1 _00417_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_152_3504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11604_ net268 net2681 net449 vssd1 vssd1 vccd1 vccd1 _01925_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_1081 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_142_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_38_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12584_ net1297 vssd1 vssd1 vccd1 vccd1 _00348_ sky130_fd_sc_hd__inv_2
XFILLER_0_52_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_1111 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07274__A1 _02872_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14323_ clknet_leaf_99_wb_clk_i _02087_ _00688_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[677\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09795__B _05736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07274__B2 _02870_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11535_ net2438 net485 _06785_ net511 vssd1 vssd1 vccd1 vccd1 _01978_ sky130_fd_sc_hd__a22o_1
XFILLER_0_151_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14254_ clknet_leaf_131_wb_clk_i _02018_ _00619_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[608\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_123_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11466_ net655 _06591_ vssd1 vssd1 vccd1 vccd1 _06769_ sky130_fd_sc_hd__nor2_1
XANTENNA__11358__B1 net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07026__A1 net1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_1974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13205_ net1276 vssd1 vssd1 vccd1 vccd1 _00969_ sky130_fd_sc_hd__inv_2
X_10417_ net304 net303 _06067_ _06239_ vssd1 vssd1 vccd1 vccd1 _06240_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_78_1985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09566__A3 _05125_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14185_ clknet_leaf_77_wb_clk_i _01949_ _00550_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[539\]
+ sky130_fd_sc_hd__dfrtp_1
X_11397_ net650 _06459_ vssd1 vssd1 vccd1 vccd1 _06751_ sky130_fd_sc_hd__or2_4
XANTENNA__12007__A net1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08774__A1 net1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13136_ net1403 vssd1 vssd1 vccd1 vccd1 _00900_ sky130_fd_sc_hd__inv_2
X_10348_ _06107_ _06109_ vssd1 vssd1 vccd1 vccd1 _06183_ sky130_fd_sc_hd__xor2_1
XFILLER_0_21_598 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10581__B2 _03458_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10750__A _05730_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10279_ _03822_ _06117_ _06114_ vssd1 vssd1 vccd1 vccd1 _06121_ sky130_fd_sc_hd__a21bo_1
X_13067_ net1288 vssd1 vssd1 vccd1 vccd1 _00831_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08526__A1 net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09316__A net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12018_ net628 _06579_ net459 net360 net2401 vssd1 vssd1 vccd1 vccd1 _01527_ sky130_fd_sc_hd__a32o_1
XFILLER_0_174_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07762__C net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_124_2916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10884__A2 net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_2927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09603__X _05545_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12086__A1 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13969_ clknet_leaf_138_wb_clk_i _01733_ _00334_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[323\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_99 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_932 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_181_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__08385__S0 net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07490_ net1110 team_03_WB.instance_to_wrap.core.register_file.registers_state\[967\]
+ net802 team_03_WB.instance_to_wrap.core.register_file.registers_state\[999\] net1135
+ vssd1 vssd1 vccd1 vccd1 _03432_ sky130_fd_sc_hd__a221o_1
XFILLER_0_0_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07501__A2 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_100_Right_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09160_ net541 _04476_ _05101_ net553 vssd1 vssd1 vccd1 vccd1 _05102_ sky130_fd_sc_hd__a211o_1
XFILLER_0_174_968 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08890__A net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08111_ net1172 team_03_WB.instance_to_wrap.core.register_file.registers_state\[570\]
+ net876 vssd1 vssd1 vccd1 vccd1 _04053_ sky130_fd_sc_hd__and3_1
XFILLER_0_43_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09091_ net941 _05032_ _05031_ net1066 vssd1 vssd1 vccd1 vccd1 _05033_ sky130_fd_sc_hd__o211a_1
XFILLER_0_127_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11520__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08042_ net717 _03962_ _03983_ vssd1 vssd1 vccd1 vccd1 _03984_ sky130_fd_sc_hd__o21a_2
XFILLER_0_25_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold901 team_03_WB.instance_to_wrap.core.register_file.registers_state\[856\] vssd1
+ vssd1 vccd1 vccd1 net2394 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07017__A1 net1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold912 team_03_WB.instance_to_wrap.core.register_file.registers_state\[619\] vssd1
+ vssd1 vccd1 vccd1 net2405 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold923 team_03_WB.instance_to_wrap.core.register_file.registers_state\[380\] vssd1
+ vssd1 vccd1 vccd1 net2416 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08214__B1 net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold934 net135 vssd1 vssd1 vccd1 vccd1 net2427 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10136__S net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold945 team_03_WB.instance_to_wrap.core.register_file.registers_state\[568\] vssd1
+ vssd1 vccd1 vccd1 net2438 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08765__A1 net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold956 team_03_WB.instance_to_wrap.core.register_file.registers_state\[639\] vssd1
+ vssd1 vccd1 vccd1 net2449 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07568__A2 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09962__A0 _05885_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold967 team_03_WB.instance_to_wrap.core.register_file.registers_state\[464\] vssd1
+ vssd1 vccd1 vccd1 net2460 sky130_fd_sc_hd__dlygate4sd3_1
Xhold978 team_03_WB.instance_to_wrap.core.register_file.registers_state\[713\] vssd1
+ vssd1 vccd1 vccd1 net2471 sky130_fd_sc_hd__dlygate4sd3_1
X_09993_ _05878_ net1763 net288 vssd1 vssd1 vccd1 vccd1 _02721_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold989 team_03_WB.instance_to_wrap.core.register_file.registers_state\[525\] vssd1
+ vssd1 vccd1 vccd1 net2482 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10572__B2 _05882_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08944_ net1050 team_03_WB.instance_to_wrap.core.register_file.registers_state\[715\]
+ net1002 team_03_WB.instance_to_wrap.core.register_file.registers_state\[747\] net924
+ vssd1 vssd1 vccd1 vccd1 _04886_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout1013_A _04085_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_32_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08875_ net556 _04770_ net540 vssd1 vssd1 vccd1 vccd1 _04817_ sky130_fd_sc_hd__o21ai_1
XANTENNA__11875__D_N net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout473_A net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07826_ _03764_ _03767_ net817 vssd1 vssd1 vccd1 vccd1 _03768_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_98_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10875__A2 net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11194__C net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12077__A1 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09478__C1 net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout640_A net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07757_ net1165 _03697_ _03698_ vssd1 vssd1 vccd1 vccd1 _03699_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout359_X net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07688_ net1183 team_03_WB.instance_to_wrap.core.register_file.registers_state\[862\]
+ net766 team_03_WB.instance_to_wrap.core.register_file.registers_state\[894\] net1129
+ vssd1 vssd1 vccd1 vccd1 _03630_ sky130_fd_sc_hd__o221a_1
XANTENNA__07180__S net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08150__C1 net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_149_475 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09427_ _04476_ _05081_ _05126_ vssd1 vssd1 vccd1 vccd1 _05369_ sky130_fd_sc_hd__or3b_1
XFILLER_0_137_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout905_A net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout526_X net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_131 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1170_X net1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09358_ _05298_ _05299_ vssd1 vssd1 vccd1 vccd1 _05300_ sky130_fd_sc_hd__nand2_1
XFILLER_0_118_840 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11588__A0 _06468_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08008__C net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08309_ net870 _04250_ _04245_ net849 vssd1 vssd1 vccd1 vccd1 _04251_ sky130_fd_sc_hd__o211a_1
XANTENNA__11052__A2 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09289_ _05230_ vssd1 vssd1 vccd1 vccd1 _05231_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout1435_X net1435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13211__A net1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07351__S1 net1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11320_ _06505_ net2566 net406 vssd1 vssd1 vccd1 vccd1 _02125_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout895_X net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11251_ net1250 net837 net301 net670 vssd1 vssd1 vccd1 vccd1 _06693_ sky130_fd_sc_hd__and4_1
XFILLER_0_63_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11369__C net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10012__A0 _03059_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_56_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08756__A1 net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10202_ team_03_WB.instance_to_wrap.core.pc.current_pc\[2\] net676 vssd1 vssd1 vccd1
+ vccd1 _06044_ sky130_fd_sc_hd__nand2_1
XFILLER_0_63_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11182_ net642 _06671_ vssd1 vssd1 vccd1 vccd1 _06672_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_128_3005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11760__B1 net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10133_ _03565_ _05974_ vssd1 vssd1 vccd1 vccd1 _05975_ sky130_fd_sc_hd__nand2_1
XFILLER_0_101_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_73_1871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_1882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08508__A1 net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_294 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input34_A gpio_in[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09136__A net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_3352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14941_ clknet_leaf_52_wb_clk_i _02696_ _01306_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_O\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_10064_ team_03_WB.instance_to_wrap.core.decoder.inst\[11\] team_03_WB.instance_to_wrap.core.decoder.inst\[10\]
+ net1248 net1251 vssd1 vssd1 vccd1 vccd1 _05908_ sky130_fd_sc_hd__or4_1
XANTENNA__11385__B net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11512__A0 _06519_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14872_ clknet_leaf_52_wb_clk_i net1901 _01237_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.wb.prev_BUSY_O
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10866__A2 _06454_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07731__A2 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13823_ clknet_leaf_20_wb_clk_i _01587_ _00188_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[177\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_106_16 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12497__A net1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_874 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10079__B1 net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11605__S net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13754_ clknet_leaf_142_wb_clk_i _01518_ _00119_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[108\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11815__A1 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10966_ net506 net597 net263 net520 net1788 vssd1 vssd1 vccd1 vccd1 _02308_ sky130_fd_sc_hd__a32o_1
XFILLER_0_168_773 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12705_ net1281 vssd1 vssd1 vccd1 vccd1 _00469_ sky130_fd_sc_hd__inv_2
XFILLER_0_57_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_167_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_248 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13685_ clknet_leaf_126_wb_clk_i _01449_ _00050_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[39\]
+ sky130_fd_sc_hd__dfrtp_1
X_10897_ net686 _05821_ vssd1 vssd1 vccd1 vccd1 _06490_ sky130_fd_sc_hd__nand2_1
XFILLER_0_127_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12636_ net1409 vssd1 vssd1 vccd1 vccd1 _00400_ sky130_fd_sc_hd__inv_2
XANTENNA__08914__S net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_35 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11579__A0 net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10745__A _05706_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12567_ net1390 vssd1 vssd1 vccd1 vccd1 _00331_ sky130_fd_sc_hd__inv_2
XFILLER_0_81_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14306_ clknet_leaf_185_wb_clk_i _02070_ _00671_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[660\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11518_ net263 net2483 net390 vssd1 vssd1 vccd1 vccd1 _01988_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_117_2775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12498_ net1394 vssd1 vssd1 vccd1 vccd1 _00262_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_117_2786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold208 net215 vssd1 vssd1 vccd1 vccd1 net1701 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold219 _02588_ vssd1 vssd1 vccd1 vccd1 net1712 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14237_ clknet_leaf_25_wb_clk_i _02001_ _00602_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[591\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_151_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11449_ net2733 net393 _06763_ net511 vssd1 vssd1 vccd1 vccd1 _02042_ sky130_fd_sc_hd__a22o_1
XANTENNA__10003__A0 _05888_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_169_3842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11279__C net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09944__A0 _05876_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_169_3853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08747__A1 net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14168_ clknet_leaf_5_wb_clk_i _01932_ _00533_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[522\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08502__X _04444_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11751__B1 net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07955__C1 net1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13119_ net1347 vssd1 vssd1 vccd1 vccd1 _00883_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_84_Left_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06990_ _02929_ _02930_ vssd1 vssd1 vccd1 vccd1 _02932_ sky130_fd_sc_hd__or2_2
X_14099_ clknet_leaf_103_wb_clk_i _01863_ _00464_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[453\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11295__B _06550_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11503__A0 _06479_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1270 net1278 vssd1 vssd1 vccd1 vccd1 net1270 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_1_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1281 net1282 vssd1 vssd1 vccd1 vccd1 net1281 sky130_fd_sc_hd__buf_4
X_08660_ net1057 team_03_WB.instance_to_wrap.core.register_file.registers_state\[327\]
+ net1010 team_03_WB.instance_to_wrap.core.register_file.registers_state\[359\] team_03_WB.instance_to_wrap.core.decoder.inst\[17\]
+ vssd1 vssd1 vccd1 vccd1 _04602_ sky130_fd_sc_hd__a221o_1
XANTENNA__09711__A3 _05041_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1292 net1294 vssd1 vssd1 vccd1 vccd1 net1292 sky130_fd_sc_hd__buf_4
X_07611_ net1121 _03551_ _03552_ net1137 vssd1 vssd1 vccd1 vccd1 _03553_ sky130_fd_sc_hd__a211o_1
X_08591_ net438 net424 _04532_ vssd1 vssd1 vccd1 vccd1 _04533_ sky130_fd_sc_hd__nor3_1
XFILLER_0_163_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11515__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_66 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11806__A1 net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07542_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[422\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[390\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[294\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[262\]
+ net779 net1137 vssd1 vssd1 vccd1 vccd1 _03484_ sky130_fd_sc_hd__mux4_1
XFILLER_0_88_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_226 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07473_ _03413_ _03414_ net1162 vssd1 vssd1 vccd1 vccd1 _03415_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_93_Left_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_626 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11282__A2 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09212_ _03391_ _03428_ _05152_ net607 vssd1 vssd1 vccd1 vccd1 _05154_ sky130_fd_sc_hd__a31o_1
XFILLER_0_174_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10490__B1 net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_147 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07238__A1 net1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09143_ net433 net427 net590 net550 vssd1 vssd1 vccd1 vccd1 _05085_ sky130_fd_sc_hd__o31a_1
XFILLER_0_17_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11034__A2 net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08986__A1 net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13031__A net1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07300__Y _03242_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_854 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09074_ net1240 team_03_WB.instance_to_wrap.core.register_file.registers_state\[173\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[141\] net982 net927
+ vssd1 vssd1 vccd1 vccd1 _05016_ sky130_fd_sc_hd__a221o_1
XANTENNA__11990__A0 net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08025_ net745 _03963_ _03964_ _03965_ _03966_ vssd1 vssd1 vccd1 vccd1 _03967_ sky130_fd_sc_hd__o32a_1
XANTENNA__10942__X _06527_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold720 team_03_WB.instance_to_wrap.core.register_file.registers_state\[125\] vssd1
+ vssd1 vccd1 vccd1 net2213 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1130_A _02785_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold731 team_03_WB.instance_to_wrap.core.register_file.registers_state\[177\] vssd1
+ vssd1 vccd1 vccd1 net2224 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold742 team_03_WB.instance_to_wrap.core.register_file.registers_state\[116\] vssd1
+ vssd1 vccd1 vccd1 net2235 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_660 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1228_A net1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold753 team_03_WB.instance_to_wrap.core.register_file.registers_state\[596\] vssd1
+ vssd1 vccd1 vccd1 net2246 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07964__A net1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold764 team_03_WB.instance_to_wrap.core.register_file.registers_state\[264\] vssd1
+ vssd1 vccd1 vccd1 net2257 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08412__X _04354_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold775 team_03_WB.instance_to_wrap.core.register_file.registers_state\[785\] vssd1
+ vssd1 vccd1 vccd1 net2268 sky130_fd_sc_hd__dlygate4sd3_1
Xhold786 team_03_WB.instance_to_wrap.core.register_file.registers_state\[519\] vssd1
+ vssd1 vccd1 vccd1 net2279 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07410__A1 _03351_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold797 team_03_WB.instance_to_wrap.core.register_file.registers_state\[492\] vssd1
+ vssd1 vccd1 vccd1 net2290 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11486__A net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09976_ _02888_ net1846 net291 vssd1 vssd1 vccd1 vccd1 _02737_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_51_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07961__A2 _03900_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08927_ net1050 team_03_WB.instance_to_wrap.core.register_file.registers_state\[203\]
+ net1002 team_03_WB.instance_to_wrap.core.register_file.registers_state\[235\] net924
+ vssd1 vssd1 vccd1 vccd1 _04869_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_51_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout855_A net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout476_X net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08858_ net864 _04799_ _04796_ net868 vssd1 vssd1 vccd1 vccd1 _04800_ sky130_fd_sc_hd__o211a_1
X_07809_ net1191 team_03_WB.instance_to_wrap.core.register_file.registers_state\[491\]
+ net881 _03750_ vssd1 vssd1 vccd1 vccd1 _03751_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout643_X net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08789_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[930\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[898\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[802\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[770\]
+ net978 net1075 vssd1 vssd1 vccd1 vccd1 _04731_ sky130_fd_sc_hd__mux4_1
XFILLER_0_79_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_140_3260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10820_ team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[26\] net305 _06424_ net691
+ vssd1 vssd1 vccd1 vccd1 _06425_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_49_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10751_ net524 _06367_ _06368_ net529 net1562 vssd1 vssd1 vccd1 vccd1 _02441_ sky130_fd_sc_hd__a32o_1
XFILLER_0_149_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_98_wb_clk_i clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_98_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout810_X net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08674__B1 net1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_412 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout908_X net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10481__B1 net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07698__X _03640_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13470_ net1323 vssd1 vssd1 vccd1 vccd1 _01234_ sky130_fd_sc_hd__inv_2
XFILLER_0_138_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_27_wb_clk_i clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_27_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_10682_ net602 _06323_ vssd1 vssd1 vccd1 vccd1 _06324_ sky130_fd_sc_hd__nand2_1
XFILLER_0_164_264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12421_ net1353 vssd1 vssd1 vccd1 vccd1 _00185_ sky130_fd_sc_hd__inv_2
XFILLER_0_36_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_97_2369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12352_ net1399 vssd1 vssd1 vccd1 vccd1 _00116_ sky130_fd_sc_hd__inv_2
XANTENNA__11981__A0 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11303_ _06613_ net2651 net404 vssd1 vssd1 vccd1 vccd1 _02142_ sky130_fd_sc_hd__mux2_1
X_15071_ net1457 vssd1 vssd1 vccd1 vccd1 la_data_out[7] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_75_1911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_75_1922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12283_ net1362 vssd1 vssd1 vccd1 vccd1 _00047_ sky130_fd_sc_hd__inv_2
X_14022_ clknet_leaf_72_wb_clk_i _01786_ _00387_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[376\]
+ sky130_fd_sc_hd__dfrtp_1
X_11234_ net1042 _06449_ net650 net701 vssd1 vssd1 vccd1 vccd1 _06684_ sky130_fd_sc_hd__or4_4
XTAP_TAPCELL_ROW_147_3403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_3_1_0_wb_clk_i_X clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_378 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_2672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11165_ net637 _06660_ vssd1 vssd1 vccd1 vccd1 _06661_ sky130_fd_sc_hd__nor2_1
XFILLER_0_101_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_164_3750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10116_ _05947_ _05957_ _05958_ _05959_ vssd1 vssd1 vccd1 vccd1 _02667_ sky130_fd_sc_hd__o31ai_1
X_11096_ _06624_ net2697 net418 vssd1 vssd1 vccd1 vccd1 _02256_ sky130_fd_sc_hd__mux2_1
XANTENNA__08588__S0 net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10047_ net9 net1036 net909 net2778 vssd1 vssd1 vccd1 vccd1 _02684_ sky130_fd_sc_hd__o22a_1
X_14924_ clknet_leaf_42_wb_clk_i _02679_ _01289_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_O\[11\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__07165__B1 team_03_WB.instance_to_wrap.core.decoder.inst\[31\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_160_3658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold80 team_03_WB.instance_to_wrap.core.register_file.registers_state\[994\] vssd1
+ vssd1 vccd1 vccd1 net1573 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_160_3669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold91 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1004\] vssd1
+ vssd1 vccd1 vccd1 net1584 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08901__A1 net1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08362__C1 net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14855_ clknet_leaf_65_wb_clk_i net1744 _01220_ vssd1 vssd1 vccd1 vccd1 net110 sky130_fd_sc_hd__dfrtp_1
X_13806_ clknet_leaf_124_wb_clk_i _01570_ _00171_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[160\]
+ sky130_fd_sc_hd__dfrtp_1
X_14786_ clknet_leaf_100_wb_clk_i _02550_ _01151_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_I\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_11998_ _06755_ net464 net445 net2708 vssd1 vssd1 vccd1 vccd1 _01546_ sky130_fd_sc_hd__a22o_1
XFILLER_0_97_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07468__A1 net1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13737_ clknet_leaf_117_wb_clk_i _01501_ _00102_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[91\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10949_ _06532_ net2430 net521 vssd1 vssd1 vccd1 vccd1 _02311_ sky130_fd_sc_hd__mux2_1
XANTENNA__11264__A2 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_168_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12955__A net1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_2815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13668_ clknet_leaf_30_wb_clk_i _01432_ _00033_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_156_776 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_2826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11016__A2 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12619_ net1288 vssd1 vssd1 vccd1 vccd1 _00383_ sky130_fd_sc_hd__inv_2
XFILLER_0_137_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13599_ net1342 vssd1 vssd1 vccd1 vccd1 _01363_ sky130_fd_sc_hd__inv_2
XFILLER_0_143_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_171_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07120__Y _03062_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08968__A1 net1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11972__B1 net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12690__A net1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_158_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07928__C1 net1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09830_ net578 _04711_ net540 vssd1 vssd1 vccd1 vccd1 _05772_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_6_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout507 net510 vssd1 vssd1 vccd1 vccd1 net507 sky130_fd_sc_hd__clkbuf_4
Xfanout518 _06395_ vssd1 vssd1 vccd1 vccd1 net518 sky130_fd_sc_hd__buf_8
Xfanout529 _06309_ vssd1 vssd1 vccd1 vccd1 net529 sky130_fd_sc_hd__clkbuf_4
X_09761_ _05654_ _04536_ vssd1 vssd1 vccd1 vccd1 _05703_ sky130_fd_sc_hd__and2b_1
X_06973_ net1112 team_03_WB.instance_to_wrap.core.register_file.registers_state\[709\]
+ net802 team_03_WB.instance_to_wrap.core.register_file.registers_state\[741\] net736
+ vssd1 vssd1 vccd1 vccd1 _02915_ sky130_fd_sc_hd__a221o_1
XANTENNA__08111__C net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1029 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08712_ _04652_ _04653_ net856 vssd1 vssd1 vccd1 vccd1 _04654_ sky130_fd_sc_hd__o21a_1
X_09692_ _05276_ _05279_ _05207_ vssd1 vssd1 vccd1 vccd1 _05634_ sky130_fd_sc_hd__a21o_1
X_08643_ net1054 team_03_WB.instance_to_wrap.core.register_file.registers_state\[678\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[646\] net1007 net941
+ vssd1 vssd1 vccd1 vccd1 _04585_ sky130_fd_sc_hd__o221a_1
XANTENNA__07950__C net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout269_A _06532_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_822 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08574_ net1063 _04513_ _04514_ vssd1 vssd1 vccd1 vccd1 _04516_ sky130_fd_sc_hd__or3_1
XFILLER_0_89_693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1096 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07459__A1 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07525_ net1102 team_03_WB.instance_to_wrap.core.register_file.registers_state\[582\]
+ net799 team_03_WB.instance_to_wrap.core.register_file.registers_state\[614\] net747
+ vssd1 vssd1 vccd1 vccd1 _03467_ sky130_fd_sc_hd__a221o_1
XANTENNA__08656__B1 net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10937__X _06523_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1080_A _02789_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout436_A net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1178_A net1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07456_ net1089 team_03_WB.instance_to_wrap.core.register_file.registers_state\[245\]
+ net893 vssd1 vssd1 vccd1 vccd1 _03398_ sky130_fd_sc_hd__or3_1
XFILLER_0_135_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_79_2000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_162_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11007__A2 net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_44_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout603_A _06295_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07387_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[447\] net758
+ net1014 vssd1 vssd1 vccd1 vccd1 _03329_ sky130_fd_sc_hd__o21a_1
XFILLER_0_33_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_44_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1345_A net1346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09126_ net852 _05055_ _05067_ vssd1 vssd1 vccd1 vccd1 _05068_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_44_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09081__B1 net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11963__B1 net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09057_ net1047 team_03_WB.instance_to_wrap.core.register_file.registers_state\[719\]
+ net998 team_03_WB.instance_to_wrap.core.register_file.registers_state\[751\] net921
+ vssd1 vssd1 vccd1 vccd1 _04999_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout1133_X net1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08008_ net1085 team_03_WB.instance_to_wrap.core.register_file.registers_state\[881\]
+ net890 vssd1 vssd1 vccd1 vccd1 _03950_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_92_2266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold550 team_03_WB.instance_to_wrap.core.register_file.registers_state\[283\] vssd1
+ vssd1 vccd1 vccd1 net2043 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_145_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_145_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout972_A net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold561 team_03_WB.instance_to_wrap.core.register_file.registers_state\[463\] vssd1
+ vssd1 vccd1 vccd1 net2054 sky130_fd_sc_hd__dlygate4sd3_1
Xhold572 team_03_WB.instance_to_wrap.core.register_file.registers_state\[233\] vssd1
+ vssd1 vccd1 vccd1 net2065 sky130_fd_sc_hd__dlygate4sd3_1
Xhold583 team_03_WB.instance_to_wrap.core.register_file.registers_state\[529\] vssd1
+ vssd1 vccd1 vccd1 net2076 sky130_fd_sc_hd__dlygate4sd3_1
Xhold594 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[27\] vssd1 vssd1 vccd1
+ vccd1 net2087 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1300_X net1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11191__B2 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09959_ _03600_ net661 vssd1 vssd1 vccd1 vccd1 _05884_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout760_X net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_142_3300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout858_X net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12970_ net1283 vssd1 vssd1 vccd1 vccd1 _00734_ sky130_fd_sc_hd__inv_2
XANTENNA__08729__S net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07147__B1 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1250 team_03_WB.instance_to_wrap.core.register_file.registers_state\[200\] vssd1
+ vssd1 vccd1 vccd1 net2743 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1261 team_03_WB.instance_to_wrap.core.register_file.registers_state\[70\] vssd1
+ vssd1 vccd1 vccd1 net2754 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09414__A net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11921_ _06469_ net2732 net367 vssd1 vssd1 vccd1 vccd1 _01621_ sky130_fd_sc_hd__mux2_1
Xhold1272 team_03_WB.instance_to_wrap.CPU_DAT_O\[26\] vssd1 vssd1 vccd1 vccd1 net2765
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1283 team_03_WB.instance_to_wrap.CPU_DAT_O\[19\] vssd1 vssd1 vccd1 vccd1 net2776
+ sky130_fd_sc_hd__dlygate4sd3_1
X_14640_ clknet_leaf_156_wb_clk_i _02404_ _01005_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[994\]
+ sky130_fd_sc_hd__dfstp_1
X_11852_ net300 net2455 net376 vssd1 vssd1 vccd1 vccd1 _01688_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_68_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10803_ _02798_ _05866_ net316 _06404_ net693 vssd1 vssd1 vccd1 vccd1 _06411_ sky130_fd_sc_hd__o41a_2
XFILLER_0_68_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14571_ clknet_leaf_45_wb_clk_i _02335_ _00936_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[925\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11246__A2 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12775__A net1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11783_ net2129 _06616_ net330 vssd1 vssd1 vccd1 vccd1 _01755_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_1124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_2409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13522_ net1307 vssd1 vssd1 vccd1 vccd1 _01286_ sky130_fd_sc_hd__inv_2
XANTENNA__07869__A net1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10734_ team_03_WB.instance_to_wrap.core.pc.current_pc\[14\] _05822_ _06295_ vssd1
+ vssd1 vccd1 vccd1 _06359_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_3159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13453_ net1343 vssd1 vssd1 vccd1 vccd1 _01217_ sky130_fd_sc_hd__inv_2
X_10665_ team_03_WB.instance_to_wrap.core.ru.state\[3\] team_03_WB.instance_to_wrap.core.ru.state\[4\]
+ team_03_WB.instance_to_wrap.core.ru.state\[5\] vssd1 vssd1 vccd1 vccd1 _06307_ sky130_fd_sc_hd__or3_1
XPHY_EDGE_ROW_149_Left_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12404_ net1305 vssd1 vssd1 vccd1 vccd1 _00168_ sky130_fd_sc_hd__inv_2
XFILLER_0_153_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13384_ net1427 vssd1 vssd1 vccd1 vccd1 _01148_ sky130_fd_sc_hd__inv_2
X_10596_ team_03_WB.instance_to_wrap.core.ru.state\[4\] _06281_ vssd1 vssd1 vccd1
+ vccd1 _06304_ sky130_fd_sc_hd__and2_1
XFILLER_0_2_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_2712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11954__B1 net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15123_ net914 vssd1 vssd1 vccd1 vccd1 net254 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_140_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_114_2723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_232 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12335_ net1336 vssd1 vssd1 vccd1 vccd1 _00099_ sky130_fd_sc_hd__inv_2
X_15054_ net1440 vssd1 vssd1 vccd1 vccd1 gpio_oeb[37] sky130_fd_sc_hd__buf_2
XFILLER_0_50_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12266_ net1279 vssd1 vssd1 vccd1 vccd1 _00030_ sky130_fd_sc_hd__inv_2
XANTENNA__11706__B1 net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14005_ clknet_leaf_106_wb_clk_i _01769_ _00370_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[359\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_120_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11217_ net271 net2056 net488 vssd1 vssd1 vccd1 vccd1 _02192_ sky130_fd_sc_hd__mux2_1
X_12197_ net1571 vssd1 vssd1 vccd1 vccd1 _02356_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_162_3709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07925__A2 net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11148_ net274 net703 net695 vssd1 vssd1 vccd1 vccd1 _06651_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_158_Left_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11079_ _06617_ net2394 net416 vssd1 vssd1 vccd1 vccd1 _02266_ sky130_fd_sc_hd__mux2_1
XANTENNA__06948__A net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09324__A _04679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14907_ clknet_leaf_54_wb_clk_i _00001_ _01272_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.ru.state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07689__A1 net1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11485__A2 net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11065__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07153__A3 net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10693__B1 net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14838_ clknet_leaf_92_wb_clk_i net1759 _01203_ vssd1 vssd1 vccd1 vccd1 net160 sky130_fd_sc_hd__dfrtp_1
X_14769_ clknet_leaf_55_wb_clk_i _02533_ _01134_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.READ_I
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08882__B _04807_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07310_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[797\] net794
+ _03246_ net1116 vssd1 vssd1 vccd1 vccd1 _03252_ sky130_fd_sc_hd__o211a_1
XFILLER_0_156_540 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08290_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[1015\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[983\]
+ net966 vssd1 vssd1 vccd1 vccd1 _04232_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_167_Left_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07241_ net1096 team_03_WB.instance_to_wrap.core.register_file.registers_state\[744\]
+ net896 vssd1 vssd1 vccd1 vccd1 _03183_ sky130_fd_sc_hd__or3_1
XFILLER_0_143_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07861__A1 net1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_144_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_448 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07172_ net1176 team_03_WB.instance_to_wrap.core.register_file.registers_state\[211\]
+ net762 team_03_WB.instance_to_wrap.core.register_file.registers_state\[243\] net741
+ vssd1 vssd1 vccd1 vccd1 _03114_ sky130_fd_sc_hd__o221a_1
XANTENNA__09063__B1 net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_171_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11945__B1 net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08106__C net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07613__A1 net1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07074__C1 net1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11960__A3 net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_996 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout304 _05925_ vssd1 vssd1 vccd1 vccd1 net304 sky130_fd_sc_hd__buf_4
Xfanout326 _06811_ vssd1 vssd1 vccd1 vccd1 net326 sky130_fd_sc_hd__clkbuf_4
X_09813_ net322 _05545_ _05650_ _05073_ vssd1 vssd1 vccd1 vccd1 _05755_ sky130_fd_sc_hd__a22o_1
Xfanout337 _06807_ vssd1 vssd1 vccd1 vccd1 net337 sky130_fd_sc_hd__buf_4
Xfanout348 _06804_ vssd1 vssd1 vccd1 vccd1 net348 sky130_fd_sc_hd__clkbuf_8
Xfanout359 _06817_ vssd1 vssd1 vccd1 vccd1 net359 sky130_fd_sc_hd__clkbuf_8
XANTENNA__09118__A1 net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout386_A net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09744_ net351 _05523_ _05678_ _05685_ vssd1 vssd1 vccd1 vccd1 _05686_ sky130_fd_sc_hd__a211o_4
X_06956_ net1112 team_03_WB.instance_to_wrap.core.register_file.registers_state\[197\]
+ net802 team_03_WB.instance_to_wrap.core.register_file.registers_state\[229\] net736
+ vssd1 vssd1 vccd1 vccd1 _02898_ sky130_fd_sc_hd__a221o_1
XANTENNA__09234__A _04235_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09675_ _03391_ _04119_ net536 _02804_ net1108 vssd1 vssd1 vccd1 vccd1 _05617_ sky130_fd_sc_hd__o32a_1
XANTENNA__11476__A2 net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout553_A net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06887_ _02792_ net1015 vssd1 vssd1 vccd1 vccd1 _02829_ sky130_fd_sc_hd__nor2_4
XANTENNA_fanout1295_A net1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08626_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[6\] net1007
+ net927 _04567_ vssd1 vssd1 vccd1 vccd1 _04568_ sky130_fd_sc_hd__o211a_1
XFILLER_0_55_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10099__B net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08557_ net1232 team_03_WB.instance_to_wrap.core.register_file.registers_state\[478\]
+ net970 team_03_WB.instance_to_wrap.core.register_file.registers_state\[510\] net1210
+ vssd1 vssd1 vccd1 vccd1 _04499_ sky130_fd_sc_hd__o221a_1
XFILLER_0_166_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10667__X _06309_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout341_X net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout439_X net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout818_A net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1083_X net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07508_ _03446_ _03449_ net819 vssd1 vssd1 vccd1 vccd1 _03450_ sky130_fd_sc_hd__o21a_1
XANTENNA__07301__A0 _03241_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08284__S net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08488_ net869 _04429_ _04424_ vssd1 vssd1 vccd1 vccd1 _04430_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_9_451 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07439_ net806 _03379_ _03380_ vssd1 vssd1 vccd1 vccd1 _03381_ sky130_fd_sc_hd__or3_1
XANTENNA__07852__A1 net1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1250_X net1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_763 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout606_X net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_2306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10450_ team_03_WB.instance_to_wrap.core.pc.current_pc\[4\] team_03_WB.instance_to_wrap.core.pc.current_pc\[3\]
+ team_03_WB.instance_to_wrap.core.pc.current_pc\[2\] team_03_WB.instance_to_wrap.core.pc.current_pc\[5\]
+ vssd1 vssd1 vccd1 vccd1 _06266_ sky130_fd_sc_hd__a31o_1
XFILLER_0_45_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_94_2317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_960 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11936__A0 net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09109_ net1051 team_03_WB.instance_to_wrap.core.register_file.registers_state\[462\]
+ net1001 team_03_WB.instance_to_wrap.core.register_file.registers_state\[494\] net1075
+ vssd1 vssd1 vccd1 vccd1 _05051_ sky130_fd_sc_hd__a221o_1
XFILLER_0_60_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08016__C net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07604__A1 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10381_ _06209_ _06210_ team_03_WB.instance_to_wrap.core.pc.current_pc\[19\] net677
+ vssd1 vssd1 vccd1 vccd1 _02653_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_131_3056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08801__B1 net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_3067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12120_ net1546 vssd1 vssd1 vccd1 vccd1 _02433_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__11951__A3 net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12051_ _06620_ net2597 net356 vssd1 vssd1 vccd1 vccd1 _01495_ sky130_fd_sc_hd__mux2_1
Xhold380 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[26\] vssd1 vssd1 vccd1
+ vccd1 net1873 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11377__C net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold391 team_03_WB.instance_to_wrap.core.register_file.registers_state\[41\] vssd1
+ vssd1 vccd1 vccd1 net1884 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11002_ net2389 net423 _06573_ net515 vssd1 vssd1 vccd1 vccd1 _02299_ sky130_fd_sc_hd__a22o_1
XANTENNA__08565__C1 net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_59_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_99_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10911__A1 net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09109__A1 net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout860 net866 vssd1 vssd1 vccd1 vccd1 net860 sky130_fd_sc_hd__buf_4
Xfanout871 net872 vssd1 vssd1 vccd1 vccd1 net871 sky130_fd_sc_hd__buf_4
Xfanout882 net887 vssd1 vssd1 vccd1 vccd1 net882 sky130_fd_sc_hd__clkbuf_2
Xfanout893 net904 vssd1 vssd1 vccd1 vccd1 net893 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08317__C1 net1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11393__B net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11467__A2 net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12953_ net1351 vssd1 vssd1 vccd1 vccd1 _00717_ sky130_fd_sc_hd__inv_2
Xhold1080 team_03_WB.instance_to_wrap.core.register_file.registers_state\[358\] vssd1
+ vssd1 vccd1 vccd1 net2573 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1091 team_03_WB.instance_to_wrap.core.register_file.registers_state\[858\] vssd1
+ vssd1 vccd1 vccd1 net2584 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08963__S0 net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_2571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11904_ net635 _06713_ net468 net373 net2030 vssd1 vssd1 vccd1 vccd1 _01637_ sky130_fd_sc_hd__a32o_1
Xclkbuf_leaf_42_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_42_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_107_2582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12884_ net1306 vssd1 vssd1 vccd1 vccd1 _00648_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_29_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_315 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14623_ clknet_leaf_168_wb_clk_i _02387_ _00988_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[977\]
+ sky130_fd_sc_hd__dfstp_1
X_11835_ _06673_ net469 net325 net2207 vssd1 vssd1 vccd1 vccd1 _01704_ sky130_fd_sc_hd__a22o_1
XANTENNA_output103_A net103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07599__A net1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14554_ clknet_leaf_148_wb_clk_i _02318_ _00919_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[908\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08096__A1 net1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11766_ _06597_ net475 net334 net2196 vssd1 vssd1 vccd1 vccd1 _01771_ sky130_fd_sc_hd__a22o_1
XFILLER_0_67_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09832__A2 _04711_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13505_ net1425 vssd1 vssd1 vccd1 vccd1 _01269_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_155_3557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10717_ net522 _06348_ _06349_ net527 net1676 vssd1 vssd1 vccd1 vccd1 _02456_ sky130_fd_sc_hd__a32o_1
XFILLER_0_125_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14485_ clknet_leaf_105_wb_clk_i _02249_ _00850_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[839\]
+ sky130_fd_sc_hd__dfrtp_1
X_11697_ _06739_ net383 net338 net2003 vssd1 vssd1 vccd1 vccd1 _01837_ sky130_fd_sc_hd__a22o_1
XANTENNA__08207__B net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13436_ net1424 vssd1 vssd1 vccd1 vccd1 _01200_ sky130_fd_sc_hd__inv_2
X_10648_ team_03_WB.instance_to_wrap.core.decoder.inst\[13\] net1715 net847 vssd1
+ vssd1 vccd1 vccd1 _02480_ sky130_fd_sc_hd__mux2_1
XANTENNA__09045__B1 net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_141_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09596__A1 _04778_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13367_ net1309 vssd1 vssd1 vccd1 vccd1 _01131_ sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_98_wb_clk_i_A clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_24_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10579_ net1721 net531 net598 _05889_ vssd1 vssd1 vccd1 vccd1 _02544_ sky130_fd_sc_hd__a22o_1
XFILLER_0_23_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15106_ net912 vssd1 vssd1 vccd1 vccd1 net241 sky130_fd_sc_hd__clkbuf_1
XANTENNA__09319__A net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12318_ net1390 vssd1 vssd1 vccd1 vccd1 _00082_ sky130_fd_sc_hd__inv_2
XANTENNA__11942__A3 net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13298_ net1340 vssd1 vssd1 vccd1 vccd1 _01062_ sky130_fd_sc_hd__inv_2
XFILLER_0_121_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15037_ clknet_leaf_93_wb_clk_i _02757_ _01402_ vssd1 vssd1 vccd1 vccd1 net193 sky130_fd_sc_hd__dfrtp_1
X_12249_ net1366 vssd1 vssd1 vccd1 vccd1 _00013_ sky130_fd_sc_hd__inv_2
XANTENNA__11287__C net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07359__B1 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09899__A2 _05735_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08556__C1 net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08020__A1 net1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10899__S net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07790_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[939\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[907\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[811\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[779\]
+ net775 net1126 vssd1 vssd1 vccd1 vccd1 _03732_ sky130_fd_sc_hd__mux4_1
XANTENNA__12104__B1 net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_147_Right_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07273__S net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09054__A net1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09460_ _05400_ _05401_ net561 vssd1 vssd1 vccd1 vccd1 _05402_ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07531__B1 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08411_ net869 _04352_ _04347_ net853 vssd1 vssd1 vccd1 vccd1 _04353_ sky130_fd_sc_hd__o211a_1
XFILLER_0_59_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09391_ _05321_ _05324_ _05332_ vssd1 vssd1 vccd1 vccd1 _05333_ sky130_fd_sc_hd__and3_1
XFILLER_0_4_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10418__B1 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08342_ net1235 team_03_WB.instance_to_wrap.core.register_file.registers_state\[85\]
+ net968 team_03_WB.instance_to_wrap.core.register_file.registers_state\[117\] net920
+ vssd1 vssd1 vccd1 vccd1 _04284_ sky130_fd_sc_hd__o221a_1
XANTENNA__08087__A1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09501__B _04444_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10969__A1 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07834__A1 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08273_ net1234 team_03_WB.instance_to_wrap.core.register_file.registers_state\[87\]
+ net964 team_03_WB.instance_to_wrap.core.register_file.registers_state\[119\] net920
+ vssd1 vssd1 vccd1 vccd1 _04215_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_15_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11630__A2 net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09928__S net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07224_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[818\] net757
+ net1041 _03165_ vssd1 vssd1 vccd1 vccd1 _03166_ sky130_fd_sc_hd__o211a_1
XANTENNA__11918__A0 _06619_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_850 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07155_ net1204 team_03_WB.instance_to_wrap.core.register_file.registers_state\[416\]
+ net885 _02870_ vssd1 vssd1 vccd1 vccd1 _03097_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout301_A _06438_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10197__A2 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11394__A1 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1043_A net1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07086_ net1196 net884 team_03_WB.instance_to_wrap.core.register_file.registers_state\[641\]
+ vssd1 vssd1 vccd1 vccd1 _03028_ sky130_fd_sc_hd__a21o_1
XFILLER_0_160_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10382__B _06144_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10950__X _06533_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1210_A net1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1308_A net1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08547__C1 net1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11697__A2 net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout291_X net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout670_A _06563_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout389_X net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout768_A net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10602__S net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07988_ net1136 _03926_ _03927_ _03929_ net1120 vssd1 vssd1 vccd1 vccd1 _03930_ sky130_fd_sc_hd__a311o_1
XANTENNA__07770__B1 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_114_Right_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09727_ _04150_ _04269_ _04326_ _04386_ net563 net560 vssd1 vssd1 vccd1 vccd1 _05669_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_87_2154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06939_ _02877_ _02878_ _02880_ _02879_ net750 net813 vssd1 vssd1 vccd1 vccd1 _02881_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_87_2165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11449__A2 net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout935_A net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11143__C_N net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09658_ _05089_ _05098_ net559 vssd1 vssd1 vccd1 vccd1 _05600_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_26_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_235 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08609_ net874 _04549_ _04550_ vssd1 vssd1 vccd1 vccd1 _04551_ sky130_fd_sc_hd__a21o_1
XFILLER_0_167_646 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09589_ _02783_ _02804_ net535 _05528_ _05530_ vssd1 vssd1 vccd1 vccd1 _05531_ sky130_fd_sc_hd__o221a_1
XFILLER_0_139_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout723_X net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11433__S net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11620_ _06694_ net382 net347 net2371 vssd1 vssd1 vccd1 vccd1 _01912_ sky130_fd_sc_hd__a22o_1
XANTENNA__13214__A net1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_318 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_132_wb_clk_i_A clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_13_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11551_ net2335 net484 _06790_ net508 vssd1 vssd1 vccd1 vccd1 _01967_ sky130_fd_sc_hd__a22o_1
XFILLER_0_9_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11621__A2 net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_3107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10502_ net129 net1030 net907 net1638 vssd1 vssd1 vccd1 vccd1 _02607_ sky130_fd_sc_hd__a22o_1
XFILLER_0_162_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14270_ clknet_leaf_114_wb_clk_i _02034_ _00635_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[624\]
+ sky130_fd_sc_hd__dfrtp_1
X_11482_ net2508 net393 _06775_ net510 vssd1 vssd1 vccd1 vccd1 _02021_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_160_wb_clk_i clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_160_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_45_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07038__C1 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13221_ net1353 vssd1 vssd1 vccd1 vccd1 _00985_ sky130_fd_sc_hd__inv_2
X_10433_ net285 _06251_ _06252_ vssd1 vssd1 vccd1 vccd1 _06253_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_150_3454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_150_3465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07589__B1 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08786__C1 net1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input64_A gpio_in[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09139__A net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13152_ net1403 vssd1 vssd1 vccd1 vccd1 _00916_ sky130_fd_sc_hd__inv_2
XFILLER_0_33_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10364_ team_03_WB.instance_to_wrap.core.pc.current_pc\[22\] net679 _06194_ _06196_
+ vssd1 vssd1 vccd1 vccd1 _02656_ sky130_fd_sc_hd__a2bb2oi_1
XANTENNA__08250__A1 net1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_59_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12103_ net634 _06677_ net466 net441 net1941 vssd1 vssd1 vccd1 vccd1 _01444_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_59_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13083_ net1364 vssd1 vssd1 vccd1 vccd1 _00847_ sky130_fd_sc_hd__inv_2
X_10295_ team_03_WB.instance_to_wrap.core.pc.current_pc\[8\] _06136_ vssd1 vssd1 vccd1
+ vccd1 _06137_ sky130_fd_sc_hd__and2_1
XANTENNA__11137__B2 net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08538__C1 net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07882__A net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12034_ net643 _06603_ net479 net362 net2068 vssd1 vssd1 vccd1 vccd1 _01511_ sky130_fd_sc_hd__a32o_1
XFILLER_0_109_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11688__A2 net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_2611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_2622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout690 _02840_ vssd1 vssd1 vccd1 vccd1 net690 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07093__S net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13985_ clknet_leaf_177_wb_clk_i _01749_ _00350_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[339\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10648__A0 team_03_WB.instance_to_wrap.core.decoder.inst\[13\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_171_wb_clk_i_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12101__A3 net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12936_ net1295 vssd1 vssd1 vccd1 vccd1 _00700_ sky130_fd_sc_hd__inv_2
XANTENNA__10112__A2 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07513__B1 net1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_157_3608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_122_2877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12867_ net1371 vssd1 vssd1 vccd1 vccd1 _00631_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_122_2888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_668 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14606_ clknet_leaf_130_wb_clk_i _02370_ _00971_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[960\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__08069__A1 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11818_ _06647_ net458 net324 net1940 vssd1 vssd1 vccd1 vccd1 _01721_ sky130_fd_sc_hd__a22o_1
XFILLER_0_28_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11570__C net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_174_3944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12798_ net1409 vssd1 vssd1 vccd1 vccd1 _00562_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_174_3955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_174_3966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_174_3977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07816__A1 net1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14537_ clknet_leaf_76_wb_clk_i _02301_ _00902_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[891\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07277__C1 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11749_ net649 _06572_ net460 net332 net2348 vssd1 vssd1 vccd1 vccd1 _01788_ sky130_fd_sc_hd__a32o_1
XANTENNA__11612__A2 net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14468_ clknet_leaf_23_wb_clk_i _02232_ _00833_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[822\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09569__B2 net1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13419_ net1427 vssd1 vssd1 vccd1 vccd1 _01183_ sky130_fd_sc_hd__inv_2
XFILLER_0_10_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14399_ clknet_leaf_172_wb_clk_i _02163_ _00764_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[753\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_10 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11376__A1 net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_144_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08777__C1 net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08241__A1 net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07675__S0 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08960_ net864 _04898_ _04901_ vssd1 vssd1 vccd1 vccd1 _04902_ sky130_fd_sc_hd__o21ai_1
XANTENNA__11128__B2 net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09336__X _05278_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07911_ net1091 team_03_WB.instance_to_wrap.core.register_file.registers_state\[847\]
+ net1150 vssd1 vssd1 vccd1 vccd1 _03853_ sky130_fd_sc_hd__a21o_1
XFILLER_0_166_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08891_ net580 _04832_ vssd1 vssd1 vccd1 vccd1 _04833_ sky130_fd_sc_hd__nor2_1
XANTENNA__11679__A2 net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07201__C1 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11518__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07842_ net1082 team_03_WB.instance_to_wrap.core.register_file.registers_state\[714\]
+ net791 team_03_WB.instance_to_wrap.core.register_file.registers_state\[746\] net725
+ vssd1 vssd1 vccd1 vccd1 _03784_ sky130_fd_sc_hd__a221o_1
X_07773_ net1133 _03711_ _03712_ _03714_ net824 vssd1 vssd1 vccd1 vccd1 _03715_ sky130_fd_sc_hd__o311ai_2
XANTENNA__10639__A0 net1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09512_ _05435_ _05453_ vssd1 vssd1 vccd1 vccd1 _05454_ sky130_fd_sc_hd__nor2_1
XFILLER_0_116_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_235 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_1019 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07504__B1 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09443_ _05378_ _05384_ net580 vssd1 vssd1 vccd1 vccd1 _05385_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_82_2051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_2062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout349_A _06804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09374_ _05143_ _05159_ _03823_ vssd1 vssd1 vccd1 vccd1 _05316_ sky130_fd_sc_hd__a21o_1
XFILLER_0_136_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_90 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07032__A net1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08325_ net850 _04266_ _04251_ vssd1 vssd1 vccd1 vccd1 _04267_ sky130_fd_sc_hd__a21oi_4
XANTENNA__07807__A1 net1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12873__A net1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout516_A net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1160_A net1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08256_ net1045 team_03_WB.instance_to_wrap.core.register_file.registers_state\[658\]
+ net995 team_03_WB.instance_to_wrap.core.register_file.registers_state\[690\] net916
+ vssd1 vssd1 vccd1 vccd1 _04198_ sky130_fd_sc_hd__a221o_1
XFILLER_0_160_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08480__A1 net1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07207_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[434\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[402\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[306\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[274\]
+ net757 net1123 vssd1 vssd1 vccd1 vccd1 _03149_ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout304_X net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08187_ net1231 team_03_WB.instance_to_wrap.core.register_file.registers_state\[339\]
+ net957 team_03_WB.instance_to_wrap.core.register_file.registers_state\[371\] net1071
+ vssd1 vssd1 vccd1 vccd1 _04129_ sky130_fd_sc_hd__o221a_1
XFILLER_0_30_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1046_X net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_104_Left_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07035__A2 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11906__A3 net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07138_ net1167 _03078_ _03079_ vssd1 vssd1 vccd1 vccd1 _03080_ sky130_fd_sc_hd__nand3_1
XFILLER_0_30_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout885_A net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11776__X _06810_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11001__B net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07069_ _03008_ _03010_ net809 vssd1 vssd1 vccd1 vccd1 _03011_ sky130_fd_sc_hd__o21a_1
Xoutput260 net260 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[6] sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout1213_X net1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10080_ _02925_ _02927_ _05918_ vssd1 vssd1 vccd1 vccd1 _05924_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_89_2205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout673_X net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_6_0_wb_clk_i_X clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10878__B1 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08310__B net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08940__C1 net1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout938_X net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_113_Left_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09496__A0 _05436_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13770_ clknet_leaf_1_wb_clk_i _01534_ _00135_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[124\]
+ sky130_fd_sc_hd__dfrtp_1
X_10982_ net1248 _06449_ net629 net701 vssd1 vssd1 vccd1 vccd1 _06560_ sky130_fd_sc_hd__or4_4
XFILLER_0_69_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12721_ net1266 vssd1 vssd1 vccd1 vccd1 _00485_ sky130_fd_sc_hd__inv_2
XFILLER_0_84_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_100_2427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_2438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12652_ net1331 vssd1 vssd1 vccd1 vccd1 _00416_ sky130_fd_sc_hd__inv_2
XFILLER_0_127_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_750 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11603_ _06536_ net2500 net449 vssd1 vssd1 vccd1 vccd1 _01926_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_152_3505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10855__X _06454_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12583_ net1387 vssd1 vssd1 vccd1 vccd1 _00347_ sky130_fd_sc_hd__inv_2
XFILLER_0_33_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_154_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1123 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14322_ clknet_leaf_164_wb_clk_i _02086_ _00687_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[676\]
+ sky130_fd_sc_hd__dfrtp_1
X_11534_ net276 net639 net704 net699 vssd1 vssd1 vccd1 vccd1 _06785_ sky130_fd_sc_hd__and4_1
XFILLER_0_20_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08471__A1 net1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08472__S net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xwire354 _04149_ vssd1 vssd1 vccd1 vccd1 net354 sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_122_Left_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_850 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14253_ clknet_leaf_189_wb_clk_i _02017_ _00618_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[607\]
+ sky130_fd_sc_hd__dfrtp_1
X_11465_ net2675 net393 _06768_ net508 vssd1 vssd1 vccd1 vccd1 _02031_ sky130_fd_sc_hd__a22o_1
XFILLER_0_80_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11358__A1 net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13204_ net1318 vssd1 vssd1 vccd1 vccd1 _00968_ sky130_fd_sc_hd__inv_2
X_10416_ _06008_ _06066_ vssd1 vssd1 vccd1 vccd1 _06239_ sky130_fd_sc_hd__and2_1
XFILLER_0_150_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input67_X net67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14184_ clknet_leaf_13_wb_clk_i _01948_ _00549_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[538\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_78_1975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09420__B1 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11396_ net516 net642 _06750_ net402 net2347 vssd1 vssd1 vccd1 vccd1 _02082_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_78_1986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13135_ net1338 vssd1 vssd1 vccd1 vccd1 _00899_ sky130_fd_sc_hd__inv_2
X_10347_ team_03_WB.instance_to_wrap.core.pc.current_pc\[25\] _06182_ net680 vssd1
+ vssd1 vccd1 vccd1 _02659_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10581__A2 net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07982__B1 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13066_ net1279 vssd1 vssd1 vccd1 vccd1 _00830_ sky130_fd_sc_hd__inv_2
X_10278_ _06119_ vssd1 vssd1 vccd1 vccd1 _06120_ sky130_fd_sc_hd__inv_2
XANTENNA__10750__B net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_1106 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1430 net1435 vssd1 vssd1 vccd1 vccd1 net1430 sky130_fd_sc_hd__buf_4
XANTENNA__13119__A net1347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12017_ _06765_ net461 net360 net2611 vssd1 vssd1 vccd1 vccd1 _01528_ sky130_fd_sc_hd__a22o_1
XANTENNA__11530__B2 net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08931__C1 net1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_2917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10884__A3 _06479_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09487__B1 _05428_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13968_ clknet_leaf_157_wb_clk_i _01732_ _00333_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[322\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_159_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_17_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11294__B1 net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12919_ net1386 vssd1 vssd1 vccd1 vccd1 _00683_ sky130_fd_sc_hd__inv_2
XANTENNA__11833__A2 net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13899_ clknet_leaf_41_wb_clk_i _01663_ _00264_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[253\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11073__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07123__Y _03065_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_150_1074 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_290 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_145_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_411 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08110_ net1087 net893 team_03_WB.instance_to_wrap.core.register_file.registers_state\[538\]
+ vssd1 vssd1 vccd1 vccd1 _04052_ sky130_fd_sc_hd__o21a_1
XANTENNA__11801__S net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08998__C1 net1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08462__A1 net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09090_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[557\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[525\]
+ net982 vssd1 vssd1 vccd1 vccd1 _05032_ sky130_fd_sc_hd__mux2_1
XFILLER_0_142_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08041_ net817 _03972_ _03982_ vssd1 vssd1 vccd1 vccd1 _03983_ sky130_fd_sc_hd__a21o_1
XANTENNA__11102__A net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold902 team_03_WB.instance_to_wrap.core.register_file.registers_state\[209\] vssd1
+ vssd1 vccd1 vccd1 net2395 sky130_fd_sc_hd__dlygate4sd3_1
Xhold913 team_03_WB.instance_to_wrap.core.register_file.registers_state\[609\] vssd1
+ vssd1 vccd1 vccd1 net2406 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08214__A1 net1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12010__A2 net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold924 team_03_WB.instance_to_wrap.core.register_file.registers_state\[540\] vssd1
+ vssd1 vccd1 vccd1 net2417 sky130_fd_sc_hd__dlygate4sd3_1
Xhold935 team_03_WB.instance_to_wrap.core.register_file.registers_state\[96\] vssd1
+ vssd1 vccd1 vccd1 net2428 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold946 team_03_WB.instance_to_wrap.core.register_file.registers_state\[592\] vssd1
+ vssd1 vccd1 vccd1 net2439 sky130_fd_sc_hd__dlygate4sd3_1
Xhold957 team_03_WB.instance_to_wrap.core.register_file.registers_state\[217\] vssd1
+ vssd1 vccd1 vccd1 net2450 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07422__C1 net1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold968 team_03_WB.instance_to_wrap.core.register_file.registers_state\[538\] vssd1
+ vssd1 vccd1 vccd1 net2461 sky130_fd_sc_hd__dlygate4sd3_1
X_09992_ _05877_ net1826 net288 vssd1 vssd1 vccd1 vccd1 _02722_ sky130_fd_sc_hd__mux2_1
Xhold979 team_03_WB.instance_to_wrap.core.register_file.registers_state\[532\] vssd1
+ vssd1 vccd1 vccd1 net2472 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10572__A2 net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08943_ net1046 team_03_WB.instance_to_wrap.core.register_file.registers_state\[587\]
+ net997 team_03_WB.instance_to_wrap.core.register_file.registers_state\[619\] net940
+ vssd1 vssd1 vccd1 vccd1 _04885_ sky130_fd_sc_hd__a221o_1
XFILLER_0_86_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09714__A1 _05073_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout299_A _06487_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08874_ _02944_ _02947_ vssd1 vssd1 vccd1 vccd1 _04816_ sky130_fd_sc_hd__or2_4
XTAP_TAPCELL_ROW_32_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07725__B1 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1006_A net1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07027__A net1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07825_ net811 _03765_ _03766_ vssd1 vssd1 vccd1 vccd1 _03767_ sky130_fd_sc_hd__and3_1
XANTENNA__11194__D net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout466_A net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07756_ net1133 _03693_ _03694_ _03696_ net1118 vssd1 vssd1 vccd1 vccd1 _03698_ sky130_fd_sc_hd__a311o_1
XANTENNA__10088__A1 net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09242__A _03391_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07489__C1 net1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11824__A2 net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07687_ _03624_ _03628_ net1146 vssd1 vssd1 vccd1 vccd1 _03629_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_17_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08150__B1 net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout633_A net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_903 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1375_A net1376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09426_ net574 _05354_ _05367_ vssd1 vssd1 vccd1 vccd1 _05368_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_149_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09357_ net590 _05297_ vssd1 vssd1 vccd1 vccd1 _05299_ sky130_fd_sc_hd__nand2_1
XFILLER_0_87_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout421_X net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout800_A net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1163_X net1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11711__S net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout519_X net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07697__A team_03_WB.instance_to_wrap.core.decoder.inst\[30\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08308_ net1225 _04248_ _04249_ vssd1 vssd1 vccd1 vccd1 _04250_ sky130_fd_sc_hd__o21a_1
XANTENNA__08453__A1 net1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08292__S net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09288_ _04646_ _05229_ vssd1 vssd1 vccd1 vccd1 _05230_ sky130_fd_sc_hd__nand2_1
XFILLER_0_133_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08239_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[50\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[18\]
+ net950 vssd1 vssd1 vccd1 vccd1 _04181_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1330_X net1330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08205__A1 net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11250_ net502 net631 _06692_ net408 net2369 vssd1 vssd1 vccd1 vccd1 _02170_ sky130_fd_sc_hd__a32o_1
XANTENNA__09402__B1 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout790_X net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout888_X net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10201_ _02990_ _06041_ vssd1 vssd1 vccd1 vccd1 _06043_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_56_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07413__C1 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11181_ net694 net715 net295 vssd1 vssd1 vccd1 vccd1 _06671_ sky130_fd_sc_hd__or3b_1
XANTENNA__10563__A2 net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_3006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10132_ _04354_ _02770_ net673 vssd1 vssd1 vccd1 vccd1 _05974_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_1872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08321__A net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09136__B _05076_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14940_ clknet_leaf_61_wb_clk_i _02695_ _01305_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_O\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_10063_ net2 net1036 net909 net2766 vssd1 vssd1 vccd1 vccd1 _02668_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_145_3353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11385__C net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07716__B1 _02871_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09704__X _05646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input27_A DAT_I[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14871_ clknet_leaf_55_wb_clk_i _02635_ _01236_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.ru.prev_busy
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10866__A3 net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13822_ clknet_leaf_118_wb_clk_i _01586_ _00187_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[176\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_173_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11276__B1 net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13753_ clknet_leaf_162_wb_clk_i _01517_ _00118_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[107\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_98_886 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10965_ net834 _06545_ vssd1 vssd1 vccd1 vccd1 _06546_ sky130_fd_sc_hd__and2_1
X_12704_ net1399 vssd1 vssd1 vccd1 vccd1 _00468_ sky130_fd_sc_hd__inv_2
XFILLER_0_168_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08692__A1 net1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13684_ clknet_leaf_124_wb_clk_i _01448_ _00049_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[38\]
+ sky130_fd_sc_hd__dfrtp_1
X_10896_ team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[14\] net307 net686 vssd1
+ vssd1 vccd1 vccd1 _06489_ sky130_fd_sc_hd__a21o_1
XANTENNA__08692__B2 net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11028__B1 net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12635_ net1361 vssd1 vssd1 vccd1 vccd1 _00399_ sky130_fd_sc_hd__inv_2
XFILLER_0_127_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_130_Left_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12566_ net1262 vssd1 vssd1 vccd1 vccd1 _00330_ sky130_fd_sc_hd__inv_2
XANTENNA__09641__B1 _05582_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10745__B net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07400__A net1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14305_ clknet_leaf_183_wb_clk_i _02069_ _00670_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[659\]
+ sky130_fd_sc_hd__dfrtp_1
X_11517_ _06631_ net2362 net390 vssd1 vssd1 vccd1 vccd1 _01989_ sky130_fd_sc_hd__mux2_1
XANTENNA__07652__C1 net1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12497_ net1267 vssd1 vssd1 vccd1 vccd1 _00261_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_117_2776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_117_2787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold209 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[24\] vssd1 vssd1 vccd1
+ vccd1 net1702 sky130_fd_sc_hd__dlygate4sd3_1
X_14236_ clknet_leaf_150_wb_clk_i _02000_ _00601_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[590\]
+ sky130_fd_sc_hd__dfrtp_1
X_11448_ net276 net629 net708 _06558_ vssd1 vssd1 vccd1 vccd1 _06763_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_169_3843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11200__A0 _06409_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_169_3854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07404__C1 net1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14167_ clknet_leaf_79_wb_clk_i _01931_ _00532_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[521\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_106_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11379_ net713 _06518_ net698 vssd1 vssd1 vccd1 vccd1 _06742_ sky130_fd_sc_hd__and3_1
XFILLER_0_42_1126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13118_ net1414 vssd1 vssd1 vccd1 vccd1 _00882_ sky130_fd_sc_hd__inv_2
XANTENNA__08231__A net1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14098_ clknet_leaf_165_wb_clk_i _01862_ _00463_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[452\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07118__Y _03060_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13049_ net1359 vssd1 vssd1 vccd1 vccd1 _00813_ sky130_fd_sc_hd__inv_2
XANTENNA__11295__C net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1260 net1263 vssd1 vssd1 vccd1 vccd1 net1260 sky130_fd_sc_hd__buf_4
XFILLER_0_79_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1271 net1273 vssd1 vssd1 vccd1 vccd1 net1271 sky130_fd_sc_hd__buf_4
XFILLER_0_56_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1282 net1283 vssd1 vssd1 vccd1 vccd1 net1282 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_1_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1293 net1294 vssd1 vssd1 vccd1 vccd1 net1293 sky130_fd_sc_hd__buf_4
XFILLER_0_79_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07610_ net1205 team_03_WB.instance_to_wrap.core.register_file.registers_state\[985\]
+ net789 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1017\] net1168
+ vssd1 vssd1 vccd1 vccd1 _03552_ sky130_fd_sc_hd__o221a_1
X_08590_ net851 _04518_ _04531_ vssd1 vssd1 vccd1 vccd1 _04532_ sky130_fd_sc_hd__o21ba_4
XANTENNA__08377__S net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12040__X _06818_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07541_ net1198 team_03_WB.instance_to_wrap.core.register_file.registers_state\[486\]
+ net884 _03482_ vssd1 vssd1 vccd1 vccd1 _03483_ sky130_fd_sc_hd__a31o_1
XFILLER_0_152_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07472_ net1184 team_03_WB.instance_to_wrap.core.register_file.registers_state\[693\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[661\] net769 net728
+ vssd1 vssd1 vccd1 vccd1 _03414_ sky130_fd_sc_hd__a221o_1
XFILLER_0_159_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09211_ net607 _05152_ vssd1 vssd1 vccd1 vccd1 _05153_ sky130_fd_sc_hd__or2_1
XFILLER_0_119_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10936__A team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[7\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_wire591_X net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09142_ net354 _04208_ net549 vssd1 vssd1 vccd1 vccd1 _05084_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_591 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_161_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09073_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[45\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[13\]
+ net982 vssd1 vssd1 vccd1 vccd1 _05015_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_866 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09181__A1_N net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09936__S net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08024_ net1177 team_03_WB.instance_to_wrap.core.register_file.registers_state\[177\]
+ net890 net1126 vssd1 vssd1 vccd1 vccd1 _03966_ sky130_fd_sc_hd__a211o_1
XFILLER_0_170_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold710 team_03_WB.instance_to_wrap.core.register_file.registers_state\[629\] vssd1
+ vssd1 vccd1 vccd1 net2203 sky130_fd_sc_hd__dlygate4sd3_1
Xhold721 team_03_WB.instance_to_wrap.core.register_file.registers_state\[531\] vssd1
+ vssd1 vccd1 vccd1 net2214 sky130_fd_sc_hd__dlygate4sd3_1
Xhold732 team_03_WB.instance_to_wrap.core.register_file.registers_state\[357\] vssd1
+ vssd1 vccd1 vccd1 net2225 sky130_fd_sc_hd__dlygate4sd3_1
Xhold743 team_03_WB.instance_to_wrap.core.register_file.registers_state\[573\] vssd1
+ vssd1 vccd1 vccd1 net2236 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold754 team_03_WB.instance_to_wrap.core.register_file.registers_state\[352\] vssd1
+ vssd1 vccd1 vccd1 net2247 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1123_A net1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold765 team_03_WB.instance_to_wrap.core.register_file.registers_state\[303\] vssd1
+ vssd1 vccd1 vccd1 net2258 sky130_fd_sc_hd__dlygate4sd3_1
Xhold776 team_03_WB.instance_to_wrap.core.register_file.registers_state\[459\] vssd1
+ vssd1 vccd1 vccd1 net2269 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11742__A1 net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold787 team_03_WB.instance_to_wrap.core.register_file.registers_state\[175\] vssd1
+ vssd1 vccd1 vccd1 net2280 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11486__B net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09975_ _02921_ net2577 net292 vssd1 vssd1 vccd1 vccd1 _02738_ sky130_fd_sc_hd__mux2_1
XANTENNA__07683__C net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold798 team_03_WB.instance_to_wrap.core.register_file.registers_state\[100\] vssd1
+ vssd1 vccd1 vccd1 net2291 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08141__A net1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08926_ net1046 team_03_WB.instance_to_wrap.core.register_file.registers_state\[75\]
+ net997 team_03_WB.instance_to_wrap.core.register_file.registers_state\[107\] net940
+ vssd1 vssd1 vccd1 vccd1 _04868_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_51_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09699__B1 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07980__A net1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1009_X net1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09794__S0 net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08857_ _04797_ _04798_ net946 vssd1 vssd1 vccd1 vccd1 _04799_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07174__A1 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout371_X net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout750_A net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout848_A net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout469_X net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07808_ net1096 team_03_WB.instance_to_wrap.core.register_file.registers_state\[459\]
+ vssd1 vssd1 vccd1 vccd1 _03750_ sky130_fd_sc_hd__and2_1
XANTENNA__10610__S net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08788_ _04728_ _04729_ vssd1 vssd1 vccd1 vccd1 _04730_ sky130_fd_sc_hd__and2_1
XFILLER_0_93_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08287__S net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_140_3250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11258__B1 net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07739_ _03669_ _03677_ net617 _03660_ vssd1 vssd1 vccd1 vccd1 _03681_ sky130_fd_sc_hd__o211a_2
XFILLER_0_79_363 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1280_X net1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout636_X net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10549__C _02837_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_240 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10750_ _05730_ net605 vssd1 vssd1 vccd1 vccd1 _06368_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_49_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09871__B1 net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09409_ net550 _04985_ _04180_ vssd1 vssd1 vccd1 vccd1 _05351_ sky130_fd_sc_hd__o21a_1
X_10681_ net313 _06314_ vssd1 vssd1 vccd1 vccd1 _06323_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_109_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout803_X net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12420_ net1357 vssd1 vssd1 vccd1 vccd1 _00184_ sky130_fd_sc_hd__inv_2
XANTENNA__13222__A net1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_165_799 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_146_991 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_2359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12351_ net1285 vssd1 vssd1 vccd1 vccd1 _00115_ sky130_fd_sc_hd__inv_2
XANTENNA__11430__B1 net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_67_wb_clk_i clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_67_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_7_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_161_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11302_ _06612_ net2637 net404 vssd1 vssd1 vccd1 vccd1 _02143_ sky130_fd_sc_hd__mux2_1
X_15070_ net1456 vssd1 vssd1 vccd1 vccd1 la_data_out[6] sky130_fd_sc_hd__buf_2
X_12282_ net1372 vssd1 vssd1 vccd1 vccd1 _00046_ sky130_fd_sc_hd__inv_2
XFILLER_0_132_162 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_1912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14021_ clknet_leaf_39_wb_clk_i _01785_ _00386_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[375\]
+ sky130_fd_sc_hd__dfrtp_1
X_11233_ net266 net2146 net488 vssd1 vssd1 vccd1 vccd1 _02178_ sky130_fd_sc_hd__mux2_1
XANTENNA__11733__A1 net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10536__A2 net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07366__S net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_2673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11164_ net694 net713 net298 vssd1 vssd1 vccd1 vccd1 _06660_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_8_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08051__A net1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_164_3740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10115_ net683 net285 team_03_WB.instance_to_wrap.core.pc.current_pc\[1\] vssd1 vssd1
+ vccd1 vccd1 _05959_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_164_3751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11095_ net834 net271 vssd1 vssd1 vccd1 vccd1 _06624_ sky130_fd_sc_hd__and2_2
XANTENNA__09154__A2 net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10046_ net10 net1040 _05906_ team_03_WB.instance_to_wrap.CPU_DAT_O\[17\] vssd1 vssd1
+ vccd1 vccd1 _02685_ sky130_fd_sc_hd__a22o_1
X_14923_ clknet_leaf_51_wb_clk_i _02678_ _01288_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_O\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08588__S1 net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10839__A3 net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_160_3659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold70 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1022\] vssd1
+ vssd1 vccd1 vccd1 net1563 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08362__B1 net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold81 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[2\] vssd1 vssd1 vccd1
+ vccd1 net1574 sky130_fd_sc_hd__dlygate4sd3_1
Xhold92 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1000\] vssd1
+ vssd1 vccd1 vccd1 net1585 sky130_fd_sc_hd__dlygate4sd3_1
X_14854_ clknet_leaf_65_wb_clk_i net1804 _01219_ vssd1 vssd1 vccd1 vccd1 net109 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_158_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13805_ clknet_leaf_182_wb_clk_i _01569_ _00170_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[159\]
+ sky130_fd_sc_hd__dfrtp_1
X_14785_ clknet_leaf_95_wb_clk_i _02549_ _01150_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_I\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_11997_ net296 net2468 net444 vssd1 vssd1 vccd1 vccd1 _01547_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10948_ _06529_ _06530_ _06531_ vssd1 vssd1 vccd1 vccd1 _06532_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_58_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13736_ clknet_leaf_7_wb_clk_i _01500_ _00101_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[90\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09610__A _05551_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_68 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10879_ net311 net310 net317 _02779_ vssd1 vssd1 vccd1 vccd1 _06475_ sky130_fd_sc_hd__a31o_2
X_13667_ clknet_leaf_30_wb_clk_i _01431_ _00032_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_2816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_119_2827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12618_ net1286 vssd1 vssd1 vccd1 vccd1 _00382_ sky130_fd_sc_hd__inv_2
XANTENNA__08417__A1 net1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13598_ net1344 vssd1 vssd1 vccd1 vccd1 _01362_ sky130_fd_sc_hd__inv_2
XFILLER_0_109_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12549_ net1355 vssd1 vssd1 vccd1 vccd1 _00313_ sky130_fd_sc_hd__inv_2
XFILLER_0_152_950 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12971__A net1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06979__A1 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11972__A1 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_1 _05870_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14219_ clknet_leaf_46_wb_clk_i _01983_ _00584_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[573\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_50_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10527__A2 net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_171 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07928__B1 net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout508 net510 vssd1 vssd1 vccd1 vccd1 net508 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_67_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout519 _06395_ vssd1 vssd1 vccd1 vccd1 net519 sky130_fd_sc_hd__clkbuf_4
X_09760_ _04777_ _05072_ _05701_ vssd1 vssd1 vccd1 vccd1 _05702_ sky130_fd_sc_hd__a21bo_1
X_06972_ net1112 team_03_WB.instance_to_wrap.core.register_file.registers_state\[581\]
+ net802 team_03_WB.instance_to_wrap.core.register_file.registers_state\[613\] net753
+ vssd1 vssd1 vccd1 vccd1 _02914_ sky130_fd_sc_hd__a221o_1
X_08711_ net1242 team_03_WB.instance_to_wrap.core.register_file.registers_state\[132\]
+ net984 team_03_WB.instance_to_wrap.core.register_file.registers_state\[164\] net944
+ vssd1 vssd1 vccd1 vccd1 _04653_ sky130_fd_sc_hd__o221a_1
X_09691_ _05623_ _05632_ vssd1 vssd1 vccd1 vccd1 _05633_ sky130_fd_sc_hd__nand2_1
Xfanout1090 net1092 vssd1 vssd1 vccd1 vccd1 net1090 sky130_fd_sc_hd__buf_2
X_08642_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[550\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[518\]
+ net983 vssd1 vssd1 vccd1 vccd1 _04584_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08573_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[445\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[413\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[317\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[285\]
+ net966 net1073 vssd1 vssd1 vccd1 vccd1 _04515_ sky130_fd_sc_hd__mux4_1
XFILLER_0_49_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08105__B1 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_166_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07524_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[678\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[646\]
+ net779 vssd1 vssd1 vccd1 vccd1 _03466_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07455_ net1184 team_03_WB.instance_to_wrap.core.register_file.registers_state\[85\]
+ net769 team_03_WB.instance_to_wrap.core.register_file.registers_state\[117\] net728
+ vssd1 vssd1 vccd1 vccd1 _03397_ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout331_A _06809_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1073_A net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_2001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_479 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07386_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[415\] net791
+ vssd1 vssd1 vccd1 vccd1 _03328_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_44_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_438 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09125_ net1081 _05060_ _05066_ vssd1 vssd1 vccd1 vccd1 _05067_ sky130_fd_sc_hd__o21ai_1
XANTENNA__10953__X _06536_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold1279_A team_03_WB.instance_to_wrap.CPU_DAT_O\[4\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09081__A1 net1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1240_A net1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10766__A2 net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11963__A1 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1338_A net1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_600 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07975__A net1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09056_ _04992_ _04997_ net875 vssd1 vssd1 vccd1 vccd1 _04998_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout798_A net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08007_ net1086 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1009\]
+ net900 _03948_ net1150 vssd1 vssd1 vccd1 vccd1 _03949_ sky130_fd_sc_hd__o311a_1
XTAP_TAPCELL_ROW_92_2256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10605__S _06304_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold540 team_03_WB.instance_to_wrap.core.register_file.registers_state\[444\] vssd1
+ vssd1 vccd1 vccd1 net2033 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_2267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold551 team_03_WB.instance_to_wrap.core.register_file.registers_state\[878\] vssd1
+ vssd1 vccd1 vccd1 net2044 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10518__A2 net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11715__A1 net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1126_X net1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold562 team_03_WB.instance_to_wrap.core.register_file.registers_state\[266\] vssd1
+ vssd1 vccd1 vccd1 net2055 sky130_fd_sc_hd__dlygate4sd3_1
Xhold573 team_03_WB.instance_to_wrap.core.register_file.registers_state\[441\] vssd1
+ vssd1 vccd1 vccd1 net2066 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_49_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold584 team_03_WB.instance_to_wrap.core.register_file.registers_state\[301\] vssd1
+ vssd1 vccd1 vccd1 net2077 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold595 team_03_WB.instance_to_wrap.core.register_file.registers_state\[691\] vssd1
+ vssd1 vccd1 vccd1 net2088 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout586_X net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout965_A net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11191__A2 net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09958_ net587 net1790 net294 vssd1 vssd1 vccd1 vccd1 _02748_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_185_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_185_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_142_3301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11479__B1 net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08909_ net1051 team_03_WB.instance_to_wrap.core.register_file.registers_state\[652\]
+ net1003 team_03_WB.instance_to_wrap.core.register_file.registers_state\[684\] net926
+ vssd1 vssd1 vccd1 vccd1 _04851_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout753_X net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09889_ net321 _05449_ _05513_ _05436_ _05830_ vssd1 vssd1 vccd1 vccd1 _05831_ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_114_wb_clk_i clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_114_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xhold1240 team_03_WB.instance_to_wrap.core.register_file.registers_state\[632\] vssd1
+ vssd1 vccd1 vccd1 net2733 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1251 team_03_WB.instance_to_wrap.core.register_file.registers_state\[218\] vssd1
+ vssd1 vccd1 vccd1 net2744 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10340__S net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10151__A0 _04178_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1262 team_03_WB.instance_to_wrap.core.register_file.registers_state\[645\] vssd1
+ vssd1 vccd1 vccd1 net2755 sky130_fd_sc_hd__dlygate4sd3_1
X_11920_ _06454_ net2582 net367 vssd1 vssd1 vccd1 vccd1 _01622_ sky130_fd_sc_hd__mux2_1
Xhold1273 team_03_WB.instance_to_wrap.CPU_DAT_O\[0\] vssd1 vssd1 vccd1 vccd1 net2766
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08895__A1 net1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1284 team_03_WB.instance_to_wrap.CPU_DAT_O\[9\] vssd1 vssd1 vccd1 vccd1 net2777
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08895__B2 net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11851_ net301 net1971 net376 vssd1 vssd1 vccd1 vccd1 _01689_ sky130_fd_sc_hd__mux2_1
XFILLER_0_170_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_169_346 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09133__C net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout920_X net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10802_ net311 net310 net317 _02778_ vssd1 vssd1 vccd1 vccd1 _06410_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_68_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_631 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14570_ clknet_leaf_6_wb_clk_i _02334_ _00935_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[924\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_71_1141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11782_ net2747 _06615_ net327 vssd1 vssd1 vccd1 vccd1 _01756_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10454__A1 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10733_ net1803 net528 net523 _06358_ vssd1 vssd1 vccd1 vccd1 _02449_ sky130_fd_sc_hd__a22o_1
X_13521_ net1306 vssd1 vssd1 vccd1 vccd1 _01285_ sky130_fd_sc_hd__inv_2
XFILLER_0_32_1136 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07855__C1 net1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13452_ net1345 vssd1 vssd1 vccd1 vccd1 _01216_ sky130_fd_sc_hd__inv_2
X_10664_ team_03_WB.instance_to_wrap.core.ru.state\[4\] team_03_WB.instance_to_wrap.core.ru.state\[5\]
+ team_03_WB.instance_to_wrap.BUSY_O vssd1 vssd1 vccd1 vccd1 _06306_ sky130_fd_sc_hd__o21a_1
XANTENNA_input94_A wbs_adr_i[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07588__C net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10295__B _06136_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_904 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10206__A1 net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11403__A0 net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12403_ net1256 vssd1 vssd1 vccd1 vccd1 _00167_ sky130_fd_sc_hd__inv_2
XFILLER_0_63_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_712 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07607__C1 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13383_ net1430 vssd1 vssd1 vccd1 vccd1 _01147_ sky130_fd_sc_hd__inv_2
XFILLER_0_134_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_88_wb_clk_i_A clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_10595_ net1142 net2004 net844 vssd1 vssd1 vccd1 vccd1 _02532_ sky130_fd_sc_hd__a21o_1
XFILLER_0_50_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_114_2713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11954__A1 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15122_ net913 vssd1 vssd1 vccd1 vccd1 net253 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_114_2724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12334_ net1268 vssd1 vssd1 vccd1 vccd1 _00098_ sky130_fd_sc_hd__inv_2
XFILLER_0_50_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15053_ net1439 vssd1 vssd1 vccd1 vccd1 gpio_oeb[36] sky130_fd_sc_hd__buf_2
XFILLER_0_120_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12265_ net1253 vssd1 vssd1 vccd1 vccd1 _00029_ sky130_fd_sc_hd__inv_2
XANTENNA__10509__A2 net1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_128_Right_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14004_ clknet_leaf_132_wb_clk_i _01768_ _00369_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[358\]
+ sky130_fd_sc_hd__dfrtp_1
X_11216_ net299 net2505 net486 vssd1 vssd1 vccd1 vccd1 _02193_ sky130_fd_sc_hd__mux2_1
XANTENNA__08032__C1 net1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12196_ net1528 vssd1 vssd1 vccd1 vccd1 _02357_ sky130_fd_sc_hd__clkbuf_1
X_11147_ net499 net649 _06650_ net413 net1953 vssd1 vssd1 vccd1 vccd1 _02231_ sky130_fd_sc_hd__a32o_1
XFILLER_0_101_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11078_ net833 _06434_ vssd1 vssd1 vccd1 vccd1 _06617_ sky130_fd_sc_hd__and2_2
XANTENNA__06948__B _02889_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14906_ clknet_leaf_54_wb_clk_i _00000_ _01271_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.ru.state\[0\]
+ sky130_fd_sc_hd__dfstp_1
X_10029_ team_03_WB.instance_to_wrap.wb.curr_state\[1\] net1 vssd1 vssd1 vccd1 vccd1
+ _05905_ sky130_fd_sc_hd__nand2_1
XFILLER_0_76_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07125__A net1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14837_ clknet_leaf_85_wb_clk_i net1730 _01202_ vssd1 vssd1 vccd1 vccd1 net159 sky130_fd_sc_hd__dfrtp_1
XANTENNA__11890__B1 net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09043__C net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_508 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08638__A1 net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14768_ clknet_leaf_54_wb_clk_i _02532_ _01133_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.i_hit
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_169_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_878 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11642__B1 net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13719_ clknet_leaf_115_wb_clk_i _01483_ _00084_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[73\]
+ sky130_fd_sc_hd__dfrtp_1
X_14699_ clknet_leaf_58_wb_clk_i _02463_ _01064_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.ADR_I\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_156_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11081__S net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_603 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07240_ net1191 team_03_WB.instance_to_wrap.core.register_file.registers_state\[968\]
+ net774 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1000\] net1154
+ vssd1 vssd1 vccd1 vccd1 _03182_ sky130_fd_sc_hd__o221a_1
XFILLER_0_116_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_246 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07171_ net1176 team_03_WB.instance_to_wrap.core.register_file.registers_state\[83\]
+ net762 team_03_WB.instance_to_wrap.core.register_file.registers_state\[115\] net726
+ vssd1 vssd1 vccd1 vccd1 _03113_ sky130_fd_sc_hd__o221a_1
XFILLER_0_82_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09063__A1 net1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10748__A2 net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11945__A1 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09339__X _05281_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07074__B1 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08271__C1 net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11110__A net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout305 net306 vssd1 vssd1 vccd1 vccd1 net305 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07377__A1 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout316 _05928_ vssd1 vssd1 vccd1 vccd1 net316 sky130_fd_sc_hd__buf_2
X_09812_ _03024_ _04957_ _05753_ _04777_ vssd1 vssd1 vccd1 vccd1 _05754_ sky130_fd_sc_hd__o211a_1
XANTENNA__07916__A3 net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout327 _06810_ vssd1 vssd1 vccd1 vccd1 net327 sky130_fd_sc_hd__buf_6
Xfanout338 _06806_ vssd1 vssd1 vccd1 vccd1 net338 sky130_fd_sc_hd__clkbuf_8
Xfanout349 _06804_ vssd1 vssd1 vccd1 vccd1 net349 sky130_fd_sc_hd__clkbuf_4
X_09743_ _05073_ _05601_ _05682_ _05684_ vssd1 vssd1 vccd1 vccd1 _05685_ sky130_fd_sc_hd__a211o_1
X_06955_ net1112 team_03_WB.instance_to_wrap.core.register_file.registers_state\[69\]
+ net802 team_03_WB.instance_to_wrap.core.register_file.registers_state\[101\] net753
+ vssd1 vssd1 vccd1 vccd1 _02897_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout281_A _06405_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout379_A net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09674_ _05614_ _05615_ net353 vssd1 vssd1 vccd1 vccd1 _05616_ sky130_fd_sc_hd__o21a_1
XFILLER_0_118_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_154_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06886_ _02823_ _02827_ vssd1 vssd1 vccd1 vccd1 _02828_ sky130_fd_sc_hd__or2_1
XANTENNA__08877__B2 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08625_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[38\] net983
+ vssd1 vssd1 vccd1 vccd1 _04567_ sky130_fd_sc_hd__or2_1
XANTENNA__11881__B1 net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1190_A net1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout546_A _03106_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1288_A net1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08629__A1 net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08556_ net1232 team_03_WB.instance_to_wrap.core.register_file.registers_state\[350\]
+ net970 team_03_WB.instance_to_wrap.core.register_file.registers_state\[382\] net1072
+ vssd1 vssd1 vccd1 vccd1 _04498_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_46_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10436__A1 _05925_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07507_ net813 _03447_ _03448_ vssd1 vssd1 vccd1 vccd1 _03449_ sky130_fd_sc_hd__and3_1
XFILLER_0_159_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_122_wb_clk_i_A clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11633__B1 net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08487_ _04425_ _04426_ _04428_ _04427_ net929 net864 vssd1 vssd1 vccd1 vccd1 _04429_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__07301__A1 _03242_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout713_A net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout334_X net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08137__Y _04079_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1076_X net1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07438_ net1179 team_03_WB.instance_to_wrap.core.register_file.registers_state\[212\]
+ net764 team_03_WB.instance_to_wrap.core.register_file.registers_state\[244\] net742
+ vssd1 vssd1 vccd1 vccd1 _03380_ sky130_fd_sc_hd__o221a_1
XFILLER_0_9_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_174_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_162_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07369_ net1114 _03309_ _03310_ _03304_ _03305_ vssd1 vssd1 vccd1 vccd1 _03311_ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout501_X net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_2307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1243_X net1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10739__A2 net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13500__A net1328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09108_ net1051 team_03_WB.instance_to_wrap.core.register_file.registers_state\[334\]
+ net1001 team_03_WB.instance_to_wrap.core.register_file.registers_state\[366\] net1214
+ vssd1 vssd1 vccd1 vccd1 _05050_ sky130_fd_sc_hd__a221o_1
XFILLER_0_60_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10380_ net282 _06145_ _06206_ net677 vssd1 vssd1 vccd1 vccd1 _06210_ sky130_fd_sc_hd__o31a_1
XFILLER_0_131_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08801__A1 net1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_3057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_131_3068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_255 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_5_wb_clk_i_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09039_ _04977_ _04978_ _04979_ _04980_ net864 net944 vssd1 vssd1 vccd1 vccd1 _04981_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_60_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11020__A net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12050_ _06619_ net2625 net356 vssd1 vssd1 vccd1 vccd1 _01496_ sky130_fd_sc_hd__mux2_1
Xhold370 team_03_WB.instance_to_wrap.ADR_I\[5\] vssd1 vssd1 vccd1 vccd1 net1863 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout870_X net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold381 team_03_WB.instance_to_wrap.core.register_file.registers_state\[393\] vssd1
+ vssd1 vccd1 vccd1 net1874 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07698__A_N net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07368__A1 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold392 net229 vssd1 vssd1 vccd1 vccd1 net1885 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout968_X net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11001_ net277 net657 net707 net830 vssd1 vssd1 vccd1 vccd1 _06573_ sky130_fd_sc_hd__and4_1
XFILLER_0_102_1130 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10911__A2 _05845_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout850 _04096_ vssd1 vssd1 vccd1 vccd1 net850 sky130_fd_sc_hd__buf_8
Xfanout861 net866 vssd1 vssd1 vccd1 vccd1 net861 sky130_fd_sc_hd__buf_4
Xfanout872 net875 vssd1 vssd1 vccd1 vccd1 net872 sky130_fd_sc_hd__clkbuf_8
Xfanout883 net884 vssd1 vssd1 vccd1 vccd1 net883 sky130_fd_sc_hd__buf_4
Xfanout894 net904 vssd1 vssd1 vccd1 vccd1 net894 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08317__B1 net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08868__A1 _02937_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11393__C net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12952_ net1380 vssd1 vssd1 vccd1 vccd1 _00716_ sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_161_wb_clk_i_A clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold1070 team_03_WB.instance_to_wrap.core.register_file.registers_state\[706\] vssd1
+ vssd1 vccd1 vccd1 net2563 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1081 team_03_WB.instance_to_wrap.core.register_file.registers_state\[74\] vssd1
+ vssd1 vccd1 vccd1 net2574 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_107_2572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11872__A0 _06545_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11903_ net639 _06712_ net473 net374 net2398 vssd1 vssd1 vccd1 vccd1 _01638_ sky130_fd_sc_hd__a32o_1
Xhold1092 team_03_WB.instance_to_wrap.core.register_file.registers_state\[871\] vssd1
+ vssd1 vccd1 vccd1 net2585 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08963__S1 net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_107_2583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12883_ net1265 vssd1 vssd1 vccd1 vccd1 _00647_ sky130_fd_sc_hd__inv_2
X_14622_ clknet_leaf_115_wb_clk_i _02386_ _00987_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[976\]
+ sky130_fd_sc_hd__dfstp_1
X_11834_ _06672_ net477 net326 net2179 vssd1 vssd1 vccd1 vccd1 _01705_ sky130_fd_sc_hd__a22o_1
XFILLER_0_157_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09817__B1 net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10427__A1 net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11624__B1 net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11765_ net646 _06595_ net451 net331 net1917 vssd1 vssd1 vccd1 vccd1 _01772_ sky130_fd_sc_hd__a32o_1
X_14553_ clknet_leaf_175_wb_clk_i _02317_ _00918_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[907\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_82_wb_clk_i clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_82_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_138_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_172_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_166_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09832__A3 net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10716_ _05842_ net603 vssd1 vssd1 vccd1 vccd1 _06349_ sky130_fd_sc_hd__nand2_1
X_13504_ net1425 vssd1 vssd1 vccd1 vccd1 _01268_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_155_3558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11696_ _06738_ net384 net340 net1996 vssd1 vssd1 vccd1 vccd1 _01838_ sky130_fd_sc_hd__a22o_1
X_14484_ clknet_leaf_132_wb_clk_i _02248_ _00849_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[838\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_11_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_11_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_130_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08207__C _04148_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13435_ net1431 vssd1 vssd1 vccd1 vccd1 _01199_ sky130_fd_sc_hd__inv_2
X_10647_ team_03_WB.instance_to_wrap.core.decoder.inst\[14\] team_03_WB.instance_to_wrap.CPU_DAT_O\[14\]
+ net846 vssd1 vssd1 vccd1 vccd1 _02481_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07111__C net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_408 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13366_ net1325 vssd1 vssd1 vccd1 vccd1 _01130_ sky130_fd_sc_hd__inv_2
XANTENNA__08253__C1 net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10578_ net1782 net531 net598 _05888_ vssd1 vssd1 vccd1 vccd1 _02545_ sky130_fd_sc_hd__a22o_1
XANTENNA__10753__B net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08504__A _04080_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15105_ net915 vssd1 vssd1 vccd1 vccd1 net240 sky130_fd_sc_hd__clkbuf_1
X_12317_ net1388 vssd1 vssd1 vccd1 vccd1 _00081_ sky130_fd_sc_hd__inv_2
X_13297_ net1340 vssd1 vssd1 vccd1 vccd1 _01061_ sky130_fd_sc_hd__inv_2
XFILLER_0_146_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15036_ clknet_leaf_87_wb_clk_i _02756_ _01401_ vssd1 vssd1 vccd1 vccd1 net192 sky130_fd_sc_hd__dfrtp_1
X_12248_ net1374 vssd1 vssd1 vccd1 vccd1 _00012_ sky130_fd_sc_hd__inv_2
XFILLER_0_107_1085 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07359__A1 net1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08556__B1 net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12179_ net1572 vssd1 vssd1 vccd1 vccd1 _02374_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__10363__B1 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11863__B1 net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08410_ _04348_ _04349_ _04351_ _04350_ net947 net865 vssd1 vssd1 vccd1 vccd1 _04352_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__11804__S net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09390_ _05323_ _05327_ vssd1 vssd1 vccd1 vccd1 _05332_ sky130_fd_sc_hd__or2_1
XFILLER_0_80_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09808__B1 net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10418__A1 net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08341_ net938 _04281_ _04282_ vssd1 vssd1 vccd1 vccd1 _04283_ sky130_fd_sc_hd__o21a_1
XFILLER_0_47_826 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_686 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1022 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11615__B1 net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10969__A2 _05082_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_61 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08272_ _04212_ _04213_ net861 vssd1 vssd1 vccd1 vccd1 _04214_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_15_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08492__C1 net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07223_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[786\] net791
+ vssd1 vssd1 vccd1 vccd1 _03165_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_17_Left_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_171_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07154_ _03093_ _03095_ net1122 vssd1 vssd1 vccd1 vccd1 _03096_ sky130_fd_sc_hd__a21o_1
XFILLER_0_6_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10663__B net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11394__A2 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07085_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[513\] net799
+ net732 _03026_ vssd1 vssd1 vccd1 vccd1 _03027_ sky130_fd_sc_hd__o211a_1
XFILLER_0_140_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1036_A net1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09944__S net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout496_A net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1203_A net1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input1_A ACK_I vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07987_ net1107 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1008\]
+ net901 _03928_ net1158 vssd1 vssd1 vccd1 vccd1 _03929_ sky130_fd_sc_hd__o311a_1
XANTENNA_fanout284_X net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09726_ net351 _05438_ _05665_ _04820_ _05667_ vssd1 vssd1 vccd1 vccd1 _05668_ sky130_fd_sc_hd__a221o_1
X_06938_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[612\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[580\]
+ net775 vssd1 vssd1 vccd1 vccd1 _02880_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_87_2155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10657__A1 team_03_WB.instance_to_wrap.CPU_DAT_O\[4\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11854__A0 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09657_ _05293_ _05298_ _05597_ _05294_ _05285_ vssd1 vssd1 vccd1 vccd1 _05599_ sky130_fd_sc_hd__a311oi_4
X_06869_ team_03_WB.instance_to_wrap.core.control_logic.instruction\[4\] team_03_WB.instance_to_wrap.core.control_logic.instruction\[5\]
+ team_03_WB.instance_to_wrap.core.control_logic.instruction\[6\] vssd1 vssd1 vccd1
+ vccd1 _02811_ sky130_fd_sc_hd__nand3b_4
XANTENNA_fanout451_X net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout830_A net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout549_X net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1193_X net1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout928_A net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_26_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11714__S net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08608_ net869 _04541_ _04544_ _04097_ vssd1 vssd1 vccd1 vccd1 _04550_ sky130_fd_sc_hd__a31o_1
XFILLER_0_96_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09588_ _04071_ _04382_ net664 _05529_ vssd1 vssd1 vccd1 vccd1 _05530_ sky130_fd_sc_hd__a22o_1
XFILLER_0_132_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11941__C net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07052__X _02994_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_658 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11606__A0 _06550_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08539_ net1063 _04479_ _04480_ vssd1 vssd1 vccd1 vccd1 _04481_ sky130_fd_sc_hd__or3_1
XFILLER_0_166_146 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_850 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout716_X net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_2480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11015__A net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07286__B1 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11550_ net655 _06660_ vssd1 vssd1 vccd1 vccd1 _06790_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_61_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_807 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_133_3108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10501_ net130 net1033 net908 net1863 vssd1 vssd1 vccd1 vccd1 _02608_ sky130_fd_sc_hd__a22o_1
XFILLER_0_163_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08027__C net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11481_ net635 net705 _06541_ net829 vssd1 vssd1 vccd1 vccd1 _06775_ sky130_fd_sc_hd__and4_1
XANTENNA__09027__A1 net1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_199 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13220_ net1370 vssd1 vssd1 vccd1 vccd1 _00984_ sky130_fd_sc_hd__inv_2
X_10432_ _06020_ _06022_ _06061_ vssd1 vssd1 vccd1 vccd1 _06252_ sky130_fd_sc_hd__or3_1
XANTENNA__07038__B1 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12031__B1 net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_150_3455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08786__B1 net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13151_ net1347 vssd1 vssd1 vccd1 vccd1 _00915_ sky130_fd_sc_hd__inv_2
XFILLER_0_104_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10363_ net283 _06147_ _06195_ net679 vssd1 vssd1 vccd1 vccd1 _06196_ sky130_fd_sc_hd__o31a_1
XFILLER_0_131_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12102_ _06797_ net468 net441 net1858 vssd1 vssd1 vccd1 vccd1 _01445_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_59_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13082_ net1378 vssd1 vssd1 vccd1 vccd1 _00846_ sky130_fd_sc_hd__inv_2
X_10294_ team_03_WB.instance_to_wrap.core.pc.current_pc\[7\] team_03_WB.instance_to_wrap.core.pc.current_pc\[6\]
+ _06135_ vssd1 vssd1 vccd1 vccd1 _06136_ sky130_fd_sc_hd__and3_1
XANTENNA_input57_A gpio_in[32] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11137__A2 net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08538__B1 net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12033_ _06774_ net470 net361 net2423 vssd1 vssd1 vccd1 vccd1 _01512_ sky130_fd_sc_hd__a22o_1
XFILLER_0_18_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07227__X _03169_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10896__A1 team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[14\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_2612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_2623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout680 net681 vssd1 vssd1 vccd1 vccd1 net680 sky130_fd_sc_hd__buf_2
Xfanout691 net693 vssd1 vssd1 vccd1 vccd1 net691 sky130_fd_sc_hd__buf_4
XANTENNA__12098__B1 net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13984_ clknet_leaf_192_wb_clk_i _01748_ _00349_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[338\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08994__A net1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09442__X _05384_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input12_X net12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_16 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11845__A0 _06413_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12935_ net1363 vssd1 vssd1 vccd1 vccd1 _00699_ sky130_fd_sc_hd__inv_2
XANTENNA__07513__A1 net1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08710__B1 net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12866_ net1350 vssd1 vssd1 vccd1 vccd1 _00630_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_122_2878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_2889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14605_ clknet_leaf_190_wb_clk_i _02369_ _00970_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[959\]
+ sky130_fd_sc_hd__dfstp_1
X_11817_ _06645_ net461 net324 net2032 vssd1 vssd1 vccd1 vccd1 _01722_ sky130_fd_sc_hd__a22o_1
XANTENNA__11570__D net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_174_3945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12797_ net1384 vssd1 vssd1 vccd1 vccd1 _00561_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_174_3956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_13 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07277__B1 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_174_3967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14536_ clknet_leaf_10_wb_clk_i _02300_ _00901_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[890\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_83_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11748_ _06571_ net475 net334 net2351 vssd1 vssd1 vccd1 vccd1 _01789_ sky130_fd_sc_hd__a22o_1
XFILLER_0_126_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09018__A1 net1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14467_ clknet_leaf_33_wb_clk_i _02231_ _00832_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[821\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09018__B2 net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11679_ _06721_ net381 net339 net1934 vssd1 vssd1 vccd1 vccd1 _01855_ sky130_fd_sc_hd__a22o_1
XFILLER_0_24_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13418_ net1431 vssd1 vssd1 vccd1 vccd1 _01182_ sky130_fd_sc_hd__inv_2
XANTENNA__09569__A2 _04235_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12022__B1 net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08226__C1 net1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08234__A net1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14398_ clknet_leaf_119_wb_clk_i _02162_ _00763_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[752\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11376__A2 net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08777__B1 net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_22 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13349_ net1329 vssd1 vssd1 vccd1 vccd1 _01113_ sky130_fd_sc_hd__inv_2
XANTENNA__10584__B1 net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07675__S1 net1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11128__A2 net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15019_ clknet_leaf_88_wb_clk_i _02739_ _01384_ vssd1 vssd1 vccd1 vccd1 net175 sky130_fd_sc_hd__dfrtp_1
X_07910_ net1163 _03845_ _03846_ _03848_ _03851_ vssd1 vssd1 vccd1 vccd1 _03852_ sky130_fd_sc_hd__a32o_1
X_08890_ net584 _04830_ vssd1 vssd1 vccd1 vccd1 _04832_ sky130_fd_sc_hd__or2_2
XFILLER_0_110_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07841_ net1082 team_03_WB.instance_to_wrap.core.register_file.registers_state\[586\]
+ net791 team_03_WB.instance_to_wrap.core.register_file.registers_state\[618\] net739
+ vssd1 vssd1 vccd1 vccd1 _03783_ sky130_fd_sc_hd__a221o_1
XFILLER_0_120_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07772_ net1118 _03704_ _03705_ _03713_ net1155 vssd1 vssd1 vccd1 vccd1 _03714_ sky130_fd_sc_hd__a311o_1
XANTENNA__12089__B1 net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06960__C1 net1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09511_ _05371_ _05438_ _05450_ _05452_ _05448_ vssd1 vssd1 vccd1 vccd1 _05453_ sky130_fd_sc_hd__a221o_2
XANTENNA__11836__B1 net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09442_ _05381_ _05383_ net566 vssd1 vssd1 vccd1 vccd1 _05384_ sky130_fd_sc_hd__mux2_2
XANTENNA__13315__A net1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09512__B _05453_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_2052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07313__A net1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09373_ _05313_ _05314_ vssd1 vssd1 vccd1 vccd1 _05315_ sky130_fd_sc_hd__nor2_1
XFILLER_0_75_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_25_Left_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08324_ _04257_ _04260_ _04265_ net867 vssd1 vssd1 vccd1 vccd1 _04266_ sky130_fd_sc_hd__a22o_1
XFILLER_0_117_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_818 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08255_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[562\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[530\]
+ net950 vssd1 vssd1 vccd1 vccd1 _04197_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout411_A _06684_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1153_A net1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout509_A net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_136 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07206_ net1170 team_03_WB.instance_to_wrap.core.register_file.registers_state\[466\]
+ net756 team_03_WB.instance_to_wrap.core.register_file.registers_state\[498\] net1149
+ vssd1 vssd1 vccd1 vccd1 _03148_ sky130_fd_sc_hd__o221a_1
XFILLER_0_7_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08217__C1 net1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12013__B1 net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08186_ net860 _04124_ _04127_ vssd1 vssd1 vccd1 vccd1 _04128_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_61_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08768__B1 net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07137_ net1109 team_03_WB.instance_to_wrap.core.register_file.registers_state\[832\]
+ net803 team_03_WB.instance_to_wrap.core.register_file.registers_state\[864\] net1156
+ vssd1 vssd1 vccd1 vccd1 _03079_ sky130_fd_sc_hd__a221o_1
XFILLER_0_162_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10961__X _06542_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1320_A net1330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10575__B1 net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1418_A net1436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11001__C net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07440__B1 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07068_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[2\] net797
+ net733 _03009_ vssd1 vssd1 vccd1 vccd1 _03010_ sky130_fd_sc_hd__o211a_1
XANTENNA__10680__Y _06322_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout780_A _02851_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput250 net250 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[23] sky130_fd_sc_hd__buf_2
XFILLER_0_30_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput261 net261 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[7] sky130_fd_sc_hd__buf_2
XANTENNA_fanout499_X net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout878_A net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07991__A1 _02872_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07991__B2 _02870_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10613__S net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1206_X net1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_2206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07194__S net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout666_X net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07743__A1 net1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08940__B1 net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09709_ _03682_ _05041_ net539 vssd1 vssd1 vccd1 vccd1 _05651_ sky130_fd_sc_hd__o21ai_1
XANTENNA__11827__B1 net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10981_ net1251 net839 vssd1 vssd1 vccd1 vccd1 _06559_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout833_X net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12095__A3 net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_2520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12720_ net1401 vssd1 vssd1 vccd1 vccd1 _00484_ sky130_fd_sc_hd__inv_2
XFILLER_0_128_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12651_ net1297 vssd1 vssd1 vccd1 vccd1 _00415_ sky130_fd_sc_hd__inv_2
XFILLER_0_78_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_2428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_2439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11602_ net269 net2413 net450 vssd1 vssd1 vccd1 vccd1 _01927_ sky130_fd_sc_hd__mux2_1
XANTENNA__08456__C1 net1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12582_ net1299 vssd1 vssd1 vccd1 vccd1 _00346_ sky130_fd_sc_hd__inv_2
XFILLER_0_93_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_152_3506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10802__A1 net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14321_ clknet_leaf_143_wb_clk_i _02085_ _00686_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[675\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11533_ net2048 net485 _06784_ net515 vssd1 vssd1 vccd1 vccd1 _01979_ sky130_fd_sc_hd__a22o_1
XFILLER_0_68_1135 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08325__Y _04267_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_160 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12004__B1 net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11464_ net655 _06589_ vssd1 vssd1 vccd1 vccd1 _06768_ sky130_fd_sc_hd__nor2_1
X_14252_ clknet_leaf_19_wb_clk_i _02016_ _00617_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[606\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11358__A2 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10415_ team_03_WB.instance_to_wrap.core.pc.current_pc\[11\] _06139_ team_03_WB.instance_to_wrap.core.pc.current_pc\[12\]
+ vssd1 vssd1 vccd1 vccd1 _06238_ sky130_fd_sc_hd__a21oi_1
X_13203_ net1267 vssd1 vssd1 vccd1 vccd1 _00967_ sky130_fd_sc_hd__inv_2
X_14183_ clknet_leaf_97_wb_clk_i _01947_ _00548_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[537\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07026__A3 net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11395_ net714 net266 net699 vssd1 vssd1 vccd1 vccd1 _06750_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_78_1976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10566__B1 net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_78_1987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12007__C net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10346_ _06179_ _06181_ net283 vssd1 vssd1 vccd1 vccd1 _06182_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13134_ net1303 vssd1 vssd1 vccd1 vccd1 _00898_ sky130_fd_sc_hd__inv_2
XANTENNA__07982__A1 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13065_ net1256 vssd1 vssd1 vccd1 vccd1 _00829_ sky130_fd_sc_hd__inv_2
X_10277_ _06115_ _06118_ vssd1 vssd1 vccd1 vccd1 _06119_ sky130_fd_sc_hd__or2_1
XFILLER_0_104_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1420 net1421 vssd1 vssd1 vccd1 vccd1 net1420 sky130_fd_sc_hd__buf_4
X_12016_ _06764_ net460 net360 net2215 vssd1 vssd1 vccd1 vccd1 _01529_ sky130_fd_sc_hd__a22o_1
XFILLER_0_104_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1431 net1435 vssd1 vssd1 vccd1 vccd1 net1431 sky130_fd_sc_hd__buf_4
XFILLER_0_139_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11530__A2 net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08931__B1 net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_124_2918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11818__B1 net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13967_ clknet_leaf_137_wb_clk_i _01731_ _00332_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[321\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10759__A _02774_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12086__A3 net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13135__A net1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11294__A1 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12918_ net1280 vssd1 vssd1 vccd1 vccd1 _00682_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_17_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08695__C1 net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13898_ clknet_leaf_1_wb_clk_i _01662_ _00263_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[252\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_75_206 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12849_ net1268 vssd1 vssd1 vccd1 vccd1 _00613_ sky130_fd_sc_hd__inv_2
XFILLER_0_75_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_150_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14519_ clknet_leaf_79_wb_clk_i _02283_ _00884_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[873\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_83_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_374 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08040_ net821 _03977_ _03979_ _03981_ net721 vssd1 vssd1 vccd1 vccd1 _03982_ sky130_fd_sc_hd__a41o_1
XFILLER_0_153_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_141_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold903 team_03_WB.instance_to_wrap.core.register_file.registers_state\[796\] vssd1
+ vssd1 vccd1 vccd1 net2396 sky130_fd_sc_hd__dlygate4sd3_1
Xhold914 team_03_WB.instance_to_wrap.core.register_file.registers_state\[667\] vssd1
+ vssd1 vccd1 vccd1 net2407 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10557__B1 net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold925 team_03_WB.instance_to_wrap.core.register_file.registers_state\[258\] vssd1
+ vssd1 vccd1 vccd1 net2418 sky130_fd_sc_hd__dlygate4sd3_1
Xhold936 team_03_WB.instance_to_wrap.core.register_file.registers_state\[852\] vssd1
+ vssd1 vccd1 vccd1 net2429 sky130_fd_sc_hd__dlygate4sd3_1
Xhold947 team_03_WB.instance_to_wrap.core.register_file.registers_state\[813\] vssd1
+ vssd1 vccd1 vccd1 net2440 sky130_fd_sc_hd__dlygate4sd3_1
Xhold958 team_03_WB.instance_to_wrap.core.register_file.registers_state\[397\] vssd1
+ vssd1 vccd1 vccd1 net2451 sky130_fd_sc_hd__dlygate4sd3_1
X_09991_ _05876_ net1791 net290 vssd1 vssd1 vccd1 vccd1 _02723_ sky130_fd_sc_hd__mux2_1
Xhold969 team_03_WB.instance_to_wrap.core.register_file.registers_state\[658\] vssd1
+ vssd1 vccd1 vccd1 net2462 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_86_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10941__B net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08942_ _04880_ _04883_ net1208 vssd1 vssd1 vccd1 vccd1 _04884_ sky130_fd_sc_hd__o21ai_1
X_08873_ _02944_ _02947_ vssd1 vssd1 vccd1 vccd1 _04815_ sky130_fd_sc_hd__nor2_1
XANTENNA__07725__A1 net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07824_ net1084 team_03_WB.instance_to_wrap.core.register_file.registers_state\[202\]
+ net792 team_03_WB.instance_to_wrap.core.register_file.registers_state\[234\] net726
+ vssd1 vssd1 vccd1 vccd1 _03766_ sky130_fd_sc_hd__a221o_1
XANTENNA__09190__A3 _04679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07755_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[428\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[396\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[300\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[268\]
+ net780 net1133 vssd1 vssd1 vccd1 vccd1 _03697_ sky130_fd_sc_hd__mux4_1
XANTENNA__12077__A3 net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout361_A _06817_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout459_A net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07489__B1 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07686_ _03626_ _03627_ net1160 vssd1 vssd1 vccd1 vccd1 _03628_ sky130_fd_sc_hd__a21o_1
XANTENNA__08139__A net1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08150__A1 net1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09425_ net564 _05366_ _05359_ net580 vssd1 vssd1 vccd1 vccd1 _05367_ sky130_fd_sc_hd__a211o_1
XFILLER_0_165_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10956__X _06538_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1270_A net1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout626_A net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1368_A net1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07978__A net1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09356_ net590 _05297_ vssd1 vssd1 vccd1 vccd1 _05298_ sky130_fd_sc_hd__or2_2
XANTENNA__11037__B2 net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06882__A team_03_WB.instance_to_wrap.core.decoder.inst\[29\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_139_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_139_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_35_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08989__B1 net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08307_ net1064 _04246_ _04247_ vssd1 vssd1 vccd1 vccd1 _04249_ sky130_fd_sc_hd__or3_1
XANTENNA__07697__B net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09287_ _03208_ _05223_ vssd1 vssd1 vccd1 vccd1 _05229_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_47_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10796__A0 net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout414_X net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1156_X net1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08238_ net550 _04179_ vssd1 vssd1 vccd1 vccd1 _04180_ sky130_fd_sc_hd__nand2_1
XFILLER_0_62_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout995_A net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_166_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08169_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[948\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[916\]
+ net958 vssd1 vssd1 vccd1 vccd1 _04111_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10200_ _02990_ _06041_ vssd1 vssd1 vccd1 vccd1 _06042_ sky130_fd_sc_hd__nor2_1
XFILLER_0_132_388 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07413__B1 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11180_ net1986 net414 _06670_ net503 vssd1 vssd1 vccd1 vccd1 _02218_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_56_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout783_X net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10131_ _03313_ _05972_ vssd1 vssd1 vccd1 vccd1 _05973_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_128_3007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11760__A2 net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_1884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10062_ net13 net1039 net911 team_03_WB.instance_to_wrap.CPU_DAT_O\[1\] vssd1 vssd1
+ vccd1 vccd1 _02669_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_145_3343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_3354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14870_ clknet_leaf_57_wb_clk_i net1588 _01235_ vssd1 vssd1 vccd1 vccd1 net127 sky130_fd_sc_hd__dfrtp_1
XANTENNA__10720__B1 net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13821_ clknet_leaf_27_wb_clk_i _01585_ _00186_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[175\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_106_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11276__A1 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09564__S1 net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13752_ clknet_leaf_186_wb_clk_i _01516_ _00117_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[106\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_74_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10964_ _06542_ _06543_ _06544_ _06399_ vssd1 vssd1 vccd1 vccd1 _06545_ sky130_fd_sc_hd__o211a_4
XANTENNA__11815__A3 net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_898 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08049__A net1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12703_ net1286 vssd1 vssd1 vccd1 vccd1 _00467_ sky130_fd_sc_hd__inv_2
X_13683_ clknet_leaf_109_wb_clk_i _01447_ _00048_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[37\]
+ sky130_fd_sc_hd__dfrtp_1
X_10895_ team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[14\] net306 vssd1
+ vssd1 vccd1 vccd1 _06488_ sky130_fd_sc_hd__and2_1
XFILLER_0_168_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11028__A1 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_959 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12634_ net1375 vssd1 vssd1 vccd1 vccd1 _00398_ sky130_fd_sc_hd__inv_2
XANTENNA__08483__S net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09641__A1 net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12565_ net1275 vssd1 vssd1 vccd1 vccd1 _00329_ sky130_fd_sc_hd__inv_2
XANTENNA__07101__C1 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_992 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14304_ clknet_leaf_187_wb_clk_i _02068_ _00669_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[658\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07652__B1 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11516_ net264 net2386 net390 vssd1 vssd1 vccd1 vccd1 _01990_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12496_ net1400 vssd1 vssd1 vccd1 vccd1 _00260_ sky130_fd_sc_hd__inv_2
XFILLER_0_103_7 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_2777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_2788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14235_ clknet_leaf_123_wb_clk_i _01999_ _00600_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[589\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11447_ net2649 net394 _06762_ net516 vssd1 vssd1 vccd1 vccd1 _02043_ sky130_fd_sc_hd__a22o_1
XFILLER_0_22_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10539__B1 net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_169_3844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08601__C1 net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11378_ net513 net640 _06741_ net403 net2022 vssd1 vssd1 vccd1 vccd1 _02091_ sky130_fd_sc_hd__a32o_1
X_14166_ clknet_leaf_153_wb_clk_i _01930_ _00531_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[520\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07955__A1 net1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11751__A2 net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10329_ _06167_ _06166_ net283 vssd1 vssd1 vccd1 vccd1 _06168_ sky130_fd_sc_hd__mux2_1
X_13117_ net1388 vssd1 vssd1 vccd1 vccd1 _00881_ sky130_fd_sc_hd__inv_2
XANTENNA__10106__X _05950_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14097_ clknet_leaf_138_wb_clk_i _01861_ _00462_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[451\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_147_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13048_ net1375 vssd1 vssd1 vccd1 vccd1 _00812_ sky130_fd_sc_hd__inv_2
XANTENNA__12969__A net1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1250 team_03_WB.instance_to_wrap.core.decoder.inst\[9\] vssd1 vssd1 vccd1 vccd1
+ net1250 sky130_fd_sc_hd__buf_4
Xfanout1261 net1263 vssd1 vssd1 vccd1 vccd1 net1261 sky130_fd_sc_hd__buf_2
Xfanout1272 net1273 vssd1 vssd1 vccd1 vccd1 net1272 sky130_fd_sc_hd__buf_4
XANTENNA__06967__A net1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1283 net1302 vssd1 vssd1 vccd1 vccd1 net1283 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_1_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1294 net1295 vssd1 vssd1 vccd1 vccd1 net1294 sky130_fd_sc_hd__buf_2
XANTENNA__08380__A1 net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14999_ clknet_leaf_10_wb_clk_i net47 _01364_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[18\]
+ sky130_fd_sc_hd__dfrtp_2
X_07540_ net1102 team_03_WB.instance_to_wrap.core.register_file.registers_state\[454\]
+ vssd1 vssd1 vccd1 vccd1 _03482_ sky130_fd_sc_hd__and2_1
XFILLER_0_159_731 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07471_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[533\] net772
+ net744 _03412_ vssd1 vssd1 vccd1 vccd1 _03413_ sky130_fd_sc_hd__a211o_1
XANTENNA__10776__X _06386_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09210_ net431 _05146_ vssd1 vssd1 vccd1 vccd1 _05152_ sky130_fd_sc_hd__nor2_1
XANTENNA__07798__A net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10490__A2 net1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10936__B net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09141_ net543 _04208_ vssd1 vssd1 vccd1 vccd1 _05083_ sky130_fd_sc_hd__nor2_1
XFILLER_0_174_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_5 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11113__A net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09072_ net550 _04985_ _05013_ vssd1 vssd1 vccd1 vccd1 _05014_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_16_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08840__C1 net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08023_ net1085 net894 team_03_WB.instance_to_wrap.core.register_file.registers_state\[145\]
+ vssd1 vssd1 vccd1 vccd1 _03965_ sky130_fd_sc_hd__o21a_1
XFILLER_0_115_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold700 team_03_WB.instance_to_wrap.core.register_file.registers_state\[369\] vssd1
+ vssd1 vccd1 vccd1 net2193 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_331 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold711 team_03_WB.instance_to_wrap.core.register_file.registers_state\[752\] vssd1
+ vssd1 vccd1 vccd1 net2204 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold722 team_03_WB.instance_to_wrap.core.register_file.registers_state\[119\] vssd1
+ vssd1 vccd1 vccd1 net2215 sky130_fd_sc_hd__dlygate4sd3_1
Xhold733 team_03_WB.instance_to_wrap.core.register_file.registers_state\[571\] vssd1
+ vssd1 vccd1 vccd1 net2226 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08738__A3 _04679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold744 team_03_WB.instance_to_wrap.core.register_file.registers_state\[337\] vssd1
+ vssd1 vccd1 vccd1 net2237 sky130_fd_sc_hd__dlygate4sd3_1
Xhold755 team_03_WB.instance_to_wrap.core.register_file.registers_state\[372\] vssd1
+ vssd1 vccd1 vccd1 net2248 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07964__C net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10671__B _05583_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_39_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_97_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold766 team_03_WB.instance_to_wrap.core.register_file.registers_state\[420\] vssd1
+ vssd1 vccd1 vccd1 net2259 sky130_fd_sc_hd__dlygate4sd3_1
Xhold777 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[8\] vssd1 vssd1 vccd1
+ vccd1 net2270 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10163__S net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold788 team_03_WB.instance_to_wrap.core.register_file.registers_state\[499\] vssd1
+ vssd1 vccd1 vccd1 net2281 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09974_ _03488_ net2668 net293 vssd1 vssd1 vccd1 vccd1 _02739_ sky130_fd_sc_hd__mux2_1
Xhold799 team_03_WB.instance_to_wrap.core.register_file.registers_state\[104\] vssd1
+ vssd1 vccd1 vccd1 net2292 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11486__C _06557_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1116_A net1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09952__S net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08925_ _04865_ _04866_ net857 vssd1 vssd1 vccd1 vccd1 _04867_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_51_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09699__A1 _04816_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12879__A net1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08856_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[672\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[640\]
+ net990 vssd1 vssd1 vccd1 vccd1 _04798_ sky130_fd_sc_hd__mux2_1
XANTENNA__10702__B1 net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11029__C_N _06495_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_1134 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07807_ net1096 team_03_WB.instance_to_wrap.core.register_file.registers_state\[331\]
+ net796 team_03_WB.instance_to_wrap.core.register_file.registers_state\[363\] net1154
+ vssd1 vssd1 vccd1 vccd1 _03749_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_98_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08787_ net1051 team_03_WB.instance_to_wrap.core.register_file.registers_state\[962\]
+ net1001 team_03_WB.instance_to_wrap.core.register_file.registers_state\[994\] net1075
+ vssd1 vssd1 vccd1 vccd1 _04729_ sky130_fd_sc_hd__a221o_1
XFILLER_0_58_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout743_A net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout364_X net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_140_3240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_3251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11258__A1 net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07738_ net611 _03679_ vssd1 vssd1 vccd1 vccd1 _03680_ sky130_fd_sc_hd__and2_1
XFILLER_0_79_375 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_904 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout531_X net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_49_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07669_ net1085 team_03_WB.instance_to_wrap.core.register_file.registers_state\[254\]
+ net890 vssd1 vssd1 vccd1 vccd1 _03611_ sky130_fd_sc_hd__or3_1
XFILLER_0_138_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout629_X net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1273_X net1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_9_Left_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13503__A net1328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09408_ _05348_ _05349_ _03064_ vssd1 vssd1 vccd1 vccd1 _05350_ sky130_fd_sc_hd__mux2_1
XANTENNA__10481__A2 net1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10680_ _06307_ net527 vssd1 vssd1 vccd1 vccd1 _06322_ sky130_fd_sc_hd__nor2_4
XFILLER_0_54_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09339_ _05204_ _05207_ _05279_ _05280_ _05201_ vssd1 vssd1 vccd1 vccd1 _05281_ sky130_fd_sc_hd__o311a_2
XFILLER_0_118_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_109_Right_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10769__B1 net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_78_wb_clk_i_A clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_8_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07634__B1 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11430__A1 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12350_ net1414 vssd1 vssd1 vccd1 vccd1 _00114_ sky130_fd_sc_hd__inv_2
XFILLER_0_62_264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout998_X net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11301_ _06611_ net2533 net405 vssd1 vssd1 vccd1 vccd1 _02144_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12281_ net1365 vssd1 vssd1 vccd1 vccd1 _00045_ sky130_fd_sc_hd__inv_2
XFILLER_0_160_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08809__S0 net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_1913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11232_ net267 net2311 net488 vssd1 vssd1 vccd1 vccd1 _02179_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_75_1924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14020_ clknet_leaf_29_wb_clk_i _01784_ _00385_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[374\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07398__C1 net1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_2674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11163_ net503 net653 _06659_ net414 net1664 vssd1 vssd1 vccd1 vccd1 _02224_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_112_2685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_36_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_36_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_101_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10114_ _05952_ _05953_ _05956_ vssd1 vssd1 vccd1 vccd1 _05958_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_164_3741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11094_ _06623_ net2465 net417 vssd1 vssd1 vccd1 vccd1 _02257_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_164_3752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10045_ net11 net1039 net911 net2745 vssd1 vssd1 vccd1 vccd1 _02686_ sky130_fd_sc_hd__a22o_1
X_14922_ clknet_leaf_42_wb_clk_i _02677_ _01287_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_O\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09154__A3 _04354_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10801__S net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08898__C1 net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold60 team_03_WB.instance_to_wrap.core.register_file.registers_state\[8\] vssd1
+ vssd1 vccd1 vccd1 net1553 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08362__A1 net1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold71 team_03_WB.instance_to_wrap.ADR_I\[20\] vssd1 vssd1 vccd1 vccd1 net1564 sky130_fd_sc_hd__dlygate4sd3_1
Xhold82 team_03_WB.instance_to_wrap.core.register_file.registers_state\[985\] vssd1
+ vssd1 vccd1 vccd1 net1575 sky130_fd_sc_hd__dlygate4sd3_1
X_14853_ clknet_leaf_66_wb_clk_i net1659 _01218_ vssd1 vssd1 vccd1 vccd1 net108 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold93 team_03_WB.instance_to_wrap.core.register_file.registers_state\[18\] vssd1
+ vssd1 vccd1 vccd1 net1586 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13804_ clknet_leaf_5_wb_clk_i _01568_ _00169_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[158\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10102__A net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14784_ clknet_leaf_104_wb_clk_i _02548_ _01149_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_I\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_11996_ _06509_ net2448 net443 vssd1 vssd1 vccd1 vccd1 _01548_ sky130_fd_sc_hd__mux2_1
XANTENNA__08114__A1 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13735_ clknet_leaf_107_wb_clk_i _01499_ _00100_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[89\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_156_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10596__X _06304_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10947_ net693 _05757_ _06399_ vssd1 vssd1 vccd1 vccd1 _06531_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_129_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_200 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13666_ clknet_leaf_172_wb_clk_i _01430_ _00031_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07873__B1 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10878_ net692 _05632_ net586 vssd1 vssd1 vccd1 vccd1 _06474_ sky130_fd_sc_hd__o21ai_2
XTAP_TAPCELL_ROW_119_2817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07411__A net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_2828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12617_ net1254 vssd1 vssd1 vccd1 vccd1 _00381_ sky130_fd_sc_hd__inv_2
XFILLER_0_54_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10248__S net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13597_ net1340 vssd1 vssd1 vccd1 vccd1 _01361_ sky130_fd_sc_hd__inv_2
XFILLER_0_171_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_170_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08822__C1 net1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12548_ net1366 vssd1 vssd1 vccd1 vccd1 _00312_ sky130_fd_sc_hd__inv_2
XANTENNA__11421__B2 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_415 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_990 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09609__Y _05551_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_686 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10772__A team_03_WB.instance_to_wrap.core.decoder.inst\[10\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12479_ net1285 vssd1 vssd1 vccd1 vccd1 _00243_ sky130_fd_sc_hd__inv_2
XANTENNA_2 net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14218_ clknet_leaf_5_wb_clk_i _01982_ _00583_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[572\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07928__A1 net1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11079__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14149_ clknet_leaf_11_wb_clk_i _01913_ _00514_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[503\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08050__B1 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout509 net510 vssd1 vssd1 vccd1 vccd1 net509 sky130_fd_sc_hd__buf_2
X_06971_ net1148 _02912_ net719 vssd1 vssd1 vccd1 vccd1 _02913_ sky130_fd_sc_hd__a21o_1
XANTENNA__11807__S net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08710_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[4\] net1013
+ net928 _04651_ vssd1 vssd1 vccd1 vccd1 _04652_ sky130_fd_sc_hd__o211a_1
XANTENNA__10711__S net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09145__A3 _04323_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09690_ net581 _05624_ _05625_ _05631_ vssd1 vssd1 vccd1 vccd1 _05632_ sky130_fd_sc_hd__a31o_2
Xfanout1080 _02789_ vssd1 vssd1 vccd1 vccd1 net1080 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07156__A2 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08641_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[934\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[902\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[806\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[774\]
+ net983 net1077 vssd1 vssd1 vccd1 vccd1 _04583_ sky130_fd_sc_hd__mux4_1
Xfanout1091 net1092 vssd1 vssd1 vccd1 vccd1 net1091 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_83_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_1070 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08572_ net1234 team_03_WB.instance_to_wrap.core.register_file.registers_state\[477\]
+ net966 team_03_WB.instance_to_wrap.core.register_file.registers_state\[509\] net1212
+ vssd1 vssd1 vccd1 vccd1 _04514_ sky130_fd_sc_hd__o221a_1
X_07523_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[550\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[518\]
+ net779 vssd1 vssd1 vccd1 vccd1 _03465_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_112_wb_clk_i_A clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_49_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13323__A net1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07454_ net744 _03392_ _03393_ _03394_ _03395_ vssd1 vssd1 vccd1 vccd1 _03396_ sky130_fd_sc_hd__o32a_1
XFILLER_0_14_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11660__A1 _06623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07321__A net1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_79_2002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07385_ _03325_ _03326_ net1160 vssd1 vssd1 vccd1 vccd1 _03327_ sky130_fd_sc_hd__o21a_1
XFILLER_0_29_283 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08136__B _03391_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout324_A _06811_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_231 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1066_A net1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07616__B1 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09124_ net868 _05065_ net848 vssd1 vssd1 vccd1 vccd1 _05066_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_44_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08704__X _04646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_143_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07092__A1 net1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09055_ net1064 _04995_ _04996_ vssd1 vssd1 vccd1 vccd1 _04997_ sky130_fd_sc_hd__a21o_1
XFILLER_0_5_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_612 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1233_A net1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08006_ net1178 team_03_WB.instance_to_wrap.core.register_file.registers_state\[977\]
+ vssd1 vssd1 vccd1 vccd1 _03948_ sky130_fd_sc_hd__or2_1
XANTENNA__09248__A _04294_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold530 team_03_WB.instance_to_wrap.core.register_file.registers_state\[841\] vssd1
+ vssd1 vccd1 vccd1 net2023 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_2257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08152__A net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold541 team_03_WB.instance_to_wrap.core.register_file.registers_state\[825\] vssd1
+ vssd1 vccd1 vccd1 net2034 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_2268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold552 team_03_WB.instance_to_wrap.core.register_file.registers_state\[63\] vssd1
+ vssd1 vccd1 vccd1 net2045 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold563 team_03_WB.instance_to_wrap.core.register_file.registers_state\[782\] vssd1
+ vssd1 vccd1 vccd1 net2056 sky130_fd_sc_hd__dlygate4sd3_1
Xhold574 team_03_WB.instance_to_wrap.core.register_file.registers_state\[712\] vssd1
+ vssd1 vccd1 vccd1 net2067 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1024 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1400_A net1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold585 team_03_WB.instance_to_wrap.core.register_file.registers_state\[257\] vssd1
+ vssd1 vccd1 vccd1 net2078 sky130_fd_sc_hd__dlygate4sd3_1
Xhold596 team_03_WB.instance_to_wrap.ADR_I\[21\] vssd1 vssd1 vccd1 vccd1 net2089 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1119_X net1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09535__X _05477_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09957_ _03844_ _03863_ net663 vssd1 vssd1 vccd1 vccd1 _05883_ sky130_fd_sc_hd__nor3_1
XANTENNA_fanout481_X net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout860_A net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout958_A net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11717__S net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11479__A1 net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08908_ _04848_ _04849_ net1221 vssd1 vssd1 vccd1 vccd1 _04850_ sky130_fd_sc_hd__o21a_1
XANTENNA__10621__S net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09888_ net1021 _03109_ _04820_ _05827_ _05829_ vssd1 vssd1 vccd1 vccd1 _05830_ sky130_fd_sc_hd__a221o_1
XANTENNA_clkbuf_leaf_151_wb_clk_i_A clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold1230 team_03_WB.instance_to_wrap.core.register_file.registers_state\[197\] vssd1
+ vssd1 vccd1 vccd1 net2723 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1241 net225 vssd1 vssd1 vccd1 vccd1 net2734 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1252 team_03_WB.instance_to_wrap.CPU_DAT_O\[18\] vssd1 vssd1 vccd1 vccd1 net2745
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08839_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[0\] net1010
+ net930 _04780_ vssd1 vssd1 vccd1 vccd1 _04781_ sky130_fd_sc_hd__o211a_1
Xhold1263 team_03_WB.instance_to_wrap.core.register_file.registers_state\[474\] vssd1
+ vssd1 vccd1 vccd1 net2756 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout746_X net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1274 team_03_WB.instance_to_wrap.core.register_file.registers_state\[198\] vssd1
+ vssd1 vccd1 vccd1 net2767 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1285 team_03_WB.instance_to_wrap.CPU_DAT_O\[16\] vssd1 vssd1 vccd1 vccd1 net2778
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_135_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11850_ net276 net2029 net376 vssd1 vssd1 vccd1 vccd1 _01690_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_154_wb_clk_i clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_154_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_169_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_68_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10801_ _06409_ net2294 net519 vssd1 vssd1 vccd1 vccd1 _02336_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_68_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11781_ net2375 _06614_ net329 vssd1 vssd1 vccd1 vccd1 _01757_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_1153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13520_ net1307 vssd1 vssd1 vccd1 vccd1 _01284_ sky130_fd_sc_hd__inv_2
X_10732_ team_03_WB.instance_to_wrap.core.pc.current_pc\[15\] _05646_ net603 vssd1
+ vssd1 vccd1 vccd1 _06358_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_24_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13451_ net1405 vssd1 vssd1 vccd1 vccd1 _01215_ sky130_fd_sc_hd__inv_2
XFILLER_0_125_406 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10663_ _06300_ net606 net1145 vssd1 vssd1 vccd1 vccd1 _06305_ sky130_fd_sc_hd__and3b_1
XFILLER_0_119_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09057__C1 net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08046__B _03987_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12402_ net1336 vssd1 vssd1 vccd1 vccd1 _00166_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07607__B1 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13382_ net1431 vssd1 vssd1 vccd1 vccd1 _01146_ sky130_fd_sc_hd__inv_2
X_10594_ team_03_WB.instance_to_wrap.core.ru.prev_busy team_03_WB.instance_to_wrap.core.ru.state\[3\]
+ _06281_ vssd1 vssd1 vccd1 vccd1 _06303_ sky130_fd_sc_hd__and3_1
XANTENNA__08804__C1 net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input87_A wbs_adr_i[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15121_ net915 vssd1 vssd1 vccd1 vccd1 net252 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_114_2714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12333_ net1332 vssd1 vssd1 vccd1 vccd1 _00097_ sky130_fd_sc_hd__inv_2
XFILLER_0_133_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_114_2725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09158__A net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15052_ net1493 vssd1 vssd1 vccd1 vccd1 gpio_oeb[4] sky130_fd_sc_hd__buf_2
X_12264_ net1292 vssd1 vssd1 vccd1 vccd1 _00028_ sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_190_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_14003_ clknet_leaf_103_wb_clk_i _01767_ _00368_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[357\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11706__A2 net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11215_ net272 net2380 net489 vssd1 vssd1 vccd1 vccd1 _02194_ sky130_fd_sc_hd__mux2_1
X_12195_ net1501 vssd1 vssd1 vccd1 vccd1 _02358_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_128_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11146_ net275 net704 net696 vssd1 vssd1 vccd1 vccd1 _06650_ sky130_fd_sc_hd__and3_1
XANTENNA__10390__A1 net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11077_ _06616_ net2534 net419 vssd1 vssd1 vccd1 vccd1 _02267_ sky130_fd_sc_hd__mux2_1
XFILLER_0_170_7 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14905_ clknet_leaf_53_wb_clk_i _00010_ _01270_ vssd1 vssd1 vccd1 vccd1 net238 sky130_fd_sc_hd__dfrtp_1
X_10028_ team_03_WB.instance_to_wrap.wb.curr_state\[1\] net1 vssd1 vssd1 vccd1 vccd1
+ _05904_ sky130_fd_sc_hd__and2_1
XANTENNA__09532__B1 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14836_ clknet_leaf_87_wb_clk_i net1856 _01201_ vssd1 vssd1 vccd1 vccd1 net157 sky130_fd_sc_hd__dfrtp_1
XANTENNA__10693__A2 net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11890__A1 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07840__S net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08099__B1 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14767_ clknet_leaf_54_wb_clk_i _02531_ _01132_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.d_hit
+ sky130_fd_sc_hd__dfrtp_4
X_11979_ net302 net2588 net444 vssd1 vssd1 vccd1 vccd1 _01565_ sky130_fd_sc_hd__mux2_1
XANTENNA__10445__A2 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13718_ clknet_leaf_179_wb_clk_i _01482_ _00083_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[72\]
+ sky130_fd_sc_hd__dfrtp_1
X_14698_ clknet_leaf_58_wb_clk_i _02462_ _01063_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.ADR_I\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07310__A2 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_171_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13649_ clknet_leaf_141_wb_clk_i _01413_ _00014_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_615 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09048__C1 net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07170_ _03110_ _03111_ net741 vssd1 vssd1 vccd1 vccd1 _03112_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06980__A net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10706__S net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11158__B1 net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11110__B net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10905__B1 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06979__X _02921_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout306 _06397_ vssd1 vssd1 vccd1 vccd1 net306 sky130_fd_sc_hd__buf_2
X_09811_ net572 _04650_ vssd1 vssd1 vccd1 vccd1 _05753_ sky130_fd_sc_hd__nand2_1
Xfanout317 net318 vssd1 vssd1 vccd1 vccd1 net317 sky130_fd_sc_hd__buf_2
Xfanout328 _06810_ vssd1 vssd1 vccd1 vccd1 net328 sky130_fd_sc_hd__buf_4
Xfanout339 _06806_ vssd1 vssd1 vccd1 vccd1 net339 sky130_fd_sc_hd__buf_4
X_09742_ _05527_ _05654_ _05683_ _04777_ vssd1 vssd1 vccd1 vccd1 _05684_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__13318__A net1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06954_ _02894_ _02895_ net736 vssd1 vssd1 vccd1 vccd1 _02896_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_1131 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09673_ net575 _05570_ vssd1 vssd1 vccd1 vccd1 _05615_ sky130_fd_sc_hd__nor2_1
XANTENNA__08877__A2 _04770_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06885_ _02808_ _02817_ _02820_ _02826_ vssd1 vssd1 vccd1 vccd1 _02827_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_118_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08624_ net435 net430 _04565_ net551 vssd1 vssd1 vccd1 vccd1 _04566_ sky130_fd_sc_hd__o31a_1
XANTENNA__11881__A1 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10948__Y _06532_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08555_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[446\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[414\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[318\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[286\]
+ net965 net1072 vssd1 vssd1 vccd1 vccd1 _04497_ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout441_A _06819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1183_A net1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout539_A net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_356 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07506_ net1109 team_03_WB.instance_to_wrap.core.register_file.registers_state\[199\]
+ net803 team_03_WB.instance_to_wrap.core.register_file.registers_state\[231\] net735
+ vssd1 vssd1 vccd1 vccd1 _03448_ sky130_fd_sc_hd__a221o_1
XANTENNA__10436__A2 _05945_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08486_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[1019\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[987\]
+ net986 vssd1 vssd1 vccd1 vccd1 _04428_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10841__C1 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07437_ net1175 team_03_WB.instance_to_wrap.core.register_file.registers_state\[84\]
+ net764 team_03_WB.instance_to_wrap.core.register_file.registers_state\[116\] net726
+ vssd1 vssd1 vccd1 vccd1 _03379_ sky130_fd_sc_hd__o221a_1
XANTENNA__10964__X _06545_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout706_A net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout327_X net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1069_X net1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07986__A net1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_3150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_787 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_99_Left_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06890__A team_03_WB.instance_to_wrap.core.decoder.inst\[12\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07368_ net725 _03299_ _03300_ net1146 vssd1 vssd1 vccd1 vccd1 _03310_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_94_2308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09107_ net862 _05047_ _05048_ _05046_ vssd1 vssd1 vccd1 vccd1 _05049_ sky130_fd_sc_hd__a31o_1
XFILLER_0_162_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_150_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10616__S net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07299_ _03217_ _03224_ _03233_ _03240_ vssd1 vssd1 vccd1 vccd1 _03241_ sky130_fd_sc_hd__o2bb2a_2
XTAP_TAPCELL_ROW_131_3058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1236_X net1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_3069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09038_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[1008\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[976\]
+ net984 vssd1 vssd1 vccd1 vccd1 _04980_ sky130_fd_sc_hd__mux2_1
XANTENNA__11149__B1 net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout696_X net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold360 _02616_ vssd1 vssd1 vccd1 vccd1 net1853 sky130_fd_sc_hd__dlygate4sd3_1
Xhold371 _02608_ vssd1 vssd1 vccd1 vccd1 net1864 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08565__A1 net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold382 team_03_WB.instance_to_wrap.core.register_file.registers_state\[548\] vssd1
+ vssd1 vccd1 vccd1 net1875 sky130_fd_sc_hd__dlygate4sd3_1
X_11000_ net497 net649 _06572_ net420 net1993 vssd1 vssd1 vccd1 vccd1 _02300_ sky130_fd_sc_hd__a32o_1
Xhold393 team_03_WB.instance_to_wrap.core.register_file.registers_state\[695\] vssd1
+ vssd1 vccd1 vccd1 net1886 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08565__B2 net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout863_X net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1042 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07773__C1 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout840 net841 vssd1 vssd1 vccd1 vccd1 net840 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10911__A3 net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13228__A net1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout851 _04096_ vssd1 vssd1 vccd1 vccd1 net851 sky130_fd_sc_hd__buf_4
XANTENNA__10351__S net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout862 net866 vssd1 vssd1 vccd1 vccd1 net862 sky130_fd_sc_hd__clkbuf_8
Xfanout873 net875 vssd1 vssd1 vccd1 vccd1 net873 sky130_fd_sc_hd__clkbuf_8
XANTENNA__08317__A1 net1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout884 net887 vssd1 vssd1 vccd1 vccd1 net884 sky130_fd_sc_hd__clkbuf_4
Xfanout895 net904 vssd1 vssd1 vccd1 vccd1 net895 sky130_fd_sc_hd__clkbuf_4
X_12951_ net1390 vssd1 vssd1 vccd1 vccd1 _00715_ sky130_fd_sc_hd__inv_2
XANTENNA__07525__C1 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1060 team_03_WB.instance_to_wrap.core.register_file.registers_state\[152\] vssd1
+ vssd1 vccd1 vccd1 net2553 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_172_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1071 team_03_WB.instance_to_wrap.core.register_file.registers_state\[834\] vssd1
+ vssd1 vccd1 vccd1 net2564 sky130_fd_sc_hd__dlygate4sd3_1
X_11902_ net643 _06711_ net479 net374 net2571 vssd1 vssd1 vccd1 vccd1 _01639_ sky130_fd_sc_hd__a32o_1
Xhold1082 team_03_WB.instance_to_wrap.core.register_file.registers_state\[148\] vssd1
+ vssd1 vccd1 vccd1 net2575 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_107_2573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1093 team_03_WB.instance_to_wrap.core.register_file.registers_state\[643\] vssd1
+ vssd1 vccd1 vccd1 net2586 sky130_fd_sc_hd__dlygate4sd3_1
X_12882_ net1395 vssd1 vssd1 vccd1 vccd1 _00646_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_29_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14621_ clknet_leaf_166_wb_clk_i _02385_ _00986_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[975\]
+ sky130_fd_sc_hd__dfstp_1
X_11833_ _06670_ net464 net325 net1800 vssd1 vssd1 vccd1 vccd1 _01706_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_159_3640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10427__A2 net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_518 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07828__B1 net1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14552_ clknet_leaf_3_wb_clk_i _02316_ _00917_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[906\]
+ sky130_fd_sc_hd__dfrtp_1
X_11764_ _06594_ net464 net333 net2274 vssd1 vssd1 vccd1 vccd1 _01773_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_161_Right_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13503_ net1328 vssd1 vssd1 vccd1 vccd1 _01267_ sky130_fd_sc_hd__inv_2
X_10715_ team_03_WB.instance_to_wrap.core.pc.current_pc\[22\] net603 vssd1 vssd1 vccd1
+ vccd1 _06348_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_155_3548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_155_3559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14483_ clknet_leaf_100_wb_clk_i _02247_ _00848_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[837\]
+ sky130_fd_sc_hd__dfrtp_1
X_11695_ _06737_ net383 net340 net1990 vssd1 vssd1 vccd1 vccd1 _01839_ sky130_fd_sc_hd__a22o_1
XANTENNA__11910__S net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13434_ net1423 vssd1 vssd1 vccd1 vccd1 _01198_ sky130_fd_sc_hd__inv_2
XFILLER_0_153_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10646_ net1235 net1849 net844 vssd1 vssd1 vccd1 vccd1 _02482_ sky130_fd_sc_hd__mux2_1
XANTENNA__09045__A2 net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11388__B1 net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13365_ net1326 vssd1 vssd1 vccd1 vccd1 _01129_ sky130_fd_sc_hd__inv_2
X_10577_ net1754 net532 net599 _05887_ vssd1 vssd1 vccd1 vccd1 _02546_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_51_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_51_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_23_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08504__B _04444_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15104_ net912 vssd1 vssd1 vccd1 vccd1 net262 sky130_fd_sc_hd__clkbuf_1
X_12316_ net1419 vssd1 vssd1 vccd1 vccd1 _00080_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13296_ net1341 vssd1 vssd1 vccd1 vccd1 _01060_ sky130_fd_sc_hd__inv_2
X_15035_ clknet_leaf_82_wb_clk_i _02755_ _01400_ vssd1 vssd1 vccd1 vccd1 net191 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12247_ net1762 vssd1 vssd1 vccd1 vccd1 _01410_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08556__A1 net1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09753__B1 _04820_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10363__A1 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12178_ net1603 vssd1 vssd1 vccd1 vccd1 _02375_ sky130_fd_sc_hd__clkbuf_1
X_15079__1465 vssd1 vssd1 vccd1 vccd1 _15079__1465/HI net1465 sky130_fd_sc_hd__conb_1
X_11129_ net1044 net836 net279 net668 vssd1 vssd1 vccd1 vccd1 _06640_ sky130_fd_sc_hd__and4_1
XFILLER_0_3_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08308__A1 net1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12104__A2 net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09903__X _05845_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09351__A _04178_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07531__A2 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14819_ clknet_leaf_95_wb_clk_i net1822 _01184_ vssd1 vssd1 vccd1 vccd1 net139 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_153_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11092__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08340_ net1235 team_03_WB.instance_to_wrap.core.register_file.registers_state\[181\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[149\] net968 net920
+ vssd1 vssd1 vccd1 vccd1 _04282_ sky130_fd_sc_hd__a221o_1
XANTENNA__07819__B1 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_698 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_123 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08271_ net1234 team_03_WB.instance_to_wrap.core.register_file.registers_state\[183\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[151\] net963 net920
+ vssd1 vssd1 vccd1 vccd1 _04213_ sky130_fd_sc_hd__a221o_1
XFILLER_0_156_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08492__B1 net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_15_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07222_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[946\] net757
+ net1014 _03163_ vssd1 vssd1 vccd1 vccd1 _03164_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_41_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_707 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07047__A1 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07153_ net1204 team_03_WB.instance_to_wrap.core.register_file.registers_state\[480\]
+ net885 _03094_ net1134 vssd1 vssd1 vccd1 vccd1 _03095_ sky130_fd_sc_hd__a311o_1
XFILLER_0_144_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10051__B1 net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07084_ net1102 team_03_WB.instance_to_wrap.core.register_file.registers_state\[545\]
+ net899 vssd1 vssd1 vccd1 vccd1 _03026_ sky130_fd_sc_hd__or3_1
XFILLER_0_70_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_39_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08547__A1 net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1029_A net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_39_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout391_A _06778_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout489_A _06680_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10024__X net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07986_ net1201 team_03_WB.instance_to_wrap.core.register_file.registers_state\[976\]
+ vssd1 vssd1 vccd1 vccd1 _03928_ sky130_fd_sc_hd__or2_1
XANTENNA__09960__S net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09725_ _03759_ _04893_ _05666_ vssd1 vssd1 vccd1 vccd1 _05667_ sky130_fd_sc_hd__a21oi_1
X_06937_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[740\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[708\]
+ net775 vssd1 vssd1 vccd1 vccd1 _02879_ sky130_fd_sc_hd__mux2_1
XANTENNA__10959__X _06541_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_2156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout277_X net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout656_A net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_2167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1398_A net1408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09656_ _05296_ _05597_ _05303_ _05285_ vssd1 vssd1 vccd1 vccd1 _05598_ sky130_fd_sc_hd__o211a_1
X_06868_ team_03_WB.instance_to_wrap.core.control_logic.instruction\[4\] team_03_WB.instance_to_wrap.core.control_logic.instruction\[5\]
+ team_03_WB.instance_to_wrap.core.control_logic.instruction\[6\] vssd1 vssd1 vccd1
+ vccd1 _02810_ sky130_fd_sc_hd__and3b_1
XFILLER_0_69_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08576__S net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14875__Q team_03_WB.instance_to_wrap.core.pc.current_pc\[4\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08607_ _04545_ _04546_ _04547_ _04548_ net865 net947 vssd1 vssd1 vccd1 vccd1 _04549_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_26_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09587_ net538 _05528_ vssd1 vssd1 vccd1 vccd1 _05529_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_65_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout823_A net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout444_X net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08158__S0 net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1186_X net1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08538_ net1234 team_03_WB.instance_to_wrap.core.register_file.registers_state\[862\]
+ net965 team_03_WB.instance_to_wrap.core.register_file.registers_state\[894\] net1072
+ vssd1 vssd1 vccd1 vccd1 _04480_ sky130_fd_sc_hd__o221a_1
XANTENNA__10200__A _02990_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_102_2470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_350 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_2481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11015__B _06468_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout611_X net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08469_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[444\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[412\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[316\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[284\]
+ net951 net1070 vssd1 vssd1 vccd1 vccd1 _04411_ sky130_fd_sc_hd__mux4_1
XANTENNA__11730__S net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout709_X net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10500_ net1686 net1035 net908 net1680 vssd1 vssd1 vccd1 vccd1 _02609_ sky130_fd_sc_hd__a22o_1
XANTENNA__10290__B1 net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_3109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11480_ net511 net639 _06604_ net394 net1887 vssd1 vssd1 vccd1 vccd1 _02022_ sky130_fd_sc_hd__a32o_1
XANTENNA__07038__A1 net1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10431_ _06020_ _06022_ _06061_ vssd1 vssd1 vccd1 vccd1 _06251_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_123_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10346__S net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_150_3445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_150_3456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09983__A0 _05868_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07589__A2 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08786__A1 net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13150_ net1410 vssd1 vssd1 vccd1 vccd1 _00914_ sky130_fd_sc_hd__inv_2
X_10362_ team_03_WB.instance_to_wrap.core.pc.current_pc\[22\] _06146_ vssd1 vssd1
+ vccd1 vccd1 _06195_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout980_X net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12101_ net639 _06675_ net473 net442 net1947 vssd1 vssd1 vccd1 vccd1 _01446_ sky130_fd_sc_hd__a32o_1
XANTENNA__07994__C1 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10293_ team_03_WB.instance_to_wrap.core.pc.current_pc\[5\] team_03_WB.instance_to_wrap.core.pc.current_pc\[4\]
+ team_03_WB.instance_to_wrap.core.pc.current_pc\[3\] team_03_WB.instance_to_wrap.core.pc.current_pc\[2\]
+ vssd1 vssd1 vccd1 vccd1 _06135_ sky130_fd_sc_hd__and4_1
X_13081_ net1352 vssd1 vssd1 vccd1 vccd1 _00845_ sky130_fd_sc_hd__inv_2
XANTENNA__08538__A1 net1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12032_ _06773_ net478 net362 net2408 vssd1 vssd1 vccd1 vccd1 _01513_ sky130_fd_sc_hd__a22o_1
Xhold190 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[30\] vssd1 vssd1 vccd1
+ vccd1 net1683 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07882__C net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07746__C1 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11542__B1 net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10896__A2 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_2613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_2624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout670 _06563_ vssd1 vssd1 vccd1 vccd1 net670 sky130_fd_sc_hd__clkbuf_4
Xfanout681 _05915_ vssd1 vssd1 vccd1 vccd1 net681 sky130_fd_sc_hd__buf_2
Xfanout692 net693 vssd1 vssd1 vccd1 vccd1 net692 sky130_fd_sc_hd__clkbuf_4
X_13983_ clknet_leaf_169_wb_clk_i _01747_ _00348_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[337\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_705 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_126_2960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12934_ net1300 vssd1 vssd1 vccd1 vccd1 _00698_ sky130_fd_sc_hd__inv_2
XANTENNA__08486__S net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_16_Right_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08171__C1 net1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12865_ net1262 vssd1 vssd1 vccd1 vccd1 _00629_ sky130_fd_sc_hd__inv_2
XFILLER_0_84_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_140_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_122_2879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14604_ clknet_leaf_15_wb_clk_i _02368_ _00969_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[958\]
+ sky130_fd_sc_hd__dfstp_1
X_11816_ _06644_ net478 net326 net1794 vssd1 vssd1 vccd1 vccd1 _01723_ sky130_fd_sc_hd__a22o_1
X_12796_ net1411 vssd1 vssd1 vccd1 vccd1 _00560_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_174_3946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_174_3957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14535_ clknet_leaf_111_wb_clk_i _02299_ _00900_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[889\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07277__A1 net1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_174_3968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11747_ net646 _06569_ net451 net331 net2416 vssd1 vssd1 vccd1 vccd1 _01790_ sky130_fd_sc_hd__a32o_1
XFILLER_0_50_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14466_ clknet_leaf_174_wb_clk_i _02230_ _00831_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[820\]
+ sky130_fd_sc_hd__dfrtp_1
X_11678_ _06720_ net381 net339 net1987 vssd1 vssd1 vccd1 vccd1 _01856_ sky130_fd_sc_hd__a22o_1
X_13417_ net1432 vssd1 vssd1 vccd1 vccd1 _01181_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09569__A3 _04820_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10629_ net2323 team_03_WB.instance_to_wrap.CPU_DAT_O\[0\] net843 vssd1 vssd1 vccd1
+ vccd1 _02499_ sky130_fd_sc_hd__mux2_1
XANTENNA__08226__B1 net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_25_Right_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14397_ clknet_leaf_24_wb_clk_i _02161_ _00762_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[751\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_144_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09974__A0 _03488_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08777__A1 net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13348_ net1326 vssd1 vssd1 vccd1 vccd1 _01112_ sky130_fd_sc_hd__inv_2
XFILLER_0_109_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10584__B2 _02888_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13279_ net1407 vssd1 vssd1 vccd1 vccd1 _01043_ sky130_fd_sc_hd__inv_2
XFILLER_0_121_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15018_ clknet_leaf_92_wb_clk_i _02738_ _01383_ vssd1 vssd1 vccd1 vccd1 net205 sky130_fd_sc_hd__dfrtp_1
XANTENNA__09346__A _04148_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10336__B2 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11087__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07201__A1 net1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07840_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[682\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[650\]
+ net760 vssd1 vssd1 vccd1 vccd1 _03782_ sky130_fd_sc_hd__mux2_1
XANTENNA__12089__A1 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07771_ net1098 team_03_WB.instance_to_wrap.core.register_file.registers_state\[876\]
+ net897 _03710_ net1165 vssd1 vssd1 vccd1 vccd1 _03713_ sky130_fd_sc_hd__o311a_1
XPHY_EDGE_ROW_34_Right_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06960__B1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09510_ net580 _05451_ net351 vssd1 vssd1 vccd1 vccd1 _05452_ sky130_fd_sc_hd__o21a_1
XFILLER_0_79_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11836__A1 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10939__B net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09441_ _04826_ _05382_ net557 vssd1 vssd1 vccd1 vccd1 _05383_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_82_2053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11116__A net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_2064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09372_ _04382_ _05312_ vssd1 vssd1 vccd1 vccd1 _05314_ sky130_fd_sc_hd__and2_1
XFILLER_0_8_1096 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08323_ net856 _04261_ _04263_ _04264_ vssd1 vssd1 vccd1 vccd1 _04265_ sky130_fd_sc_hd__a31o_1
XFILLER_0_145_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_966 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13331__A net1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08254_ _04194_ _04195_ net859 vssd1 vssd1 vccd1 vccd1 _04196_ sky130_fd_sc_hd__o21a_1
XFILLER_0_89_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_43_Right_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07205_ net1170 team_03_WB.instance_to_wrap.core.register_file.registers_state\[338\]
+ net756 team_03_WB.instance_to_wrap.core.register_file.registers_state\[370\] net1123
+ vssd1 vssd1 vccd1 vccd1 _03147_ sky130_fd_sc_hd__o221a_1
XANTENNA__08217__B1 net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12013__A1 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_148 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08185_ net855 _04125_ _04126_ vssd1 vssd1 vccd1 vccd1 _04127_ sky130_fd_sc_hd__or3_1
XFILLER_0_144_397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_340 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout404_A _06717_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08768__A1 net1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1146_A net1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07136_ net1109 team_03_WB.instance_to_wrap.core.register_file.registers_state\[960\]
+ net803 team_03_WB.instance_to_wrap.core.register_file.registers_state\[992\] net1135
+ vssd1 vssd1 vccd1 vccd1 _03078_ sky130_fd_sc_hd__a221o_1
XANTENNA__11772__B1 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07976__C1 net1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10575__B2 _05885_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07067_ net1097 team_03_WB.instance_to_wrap.core.register_file.registers_state\[34\]
+ net899 vssd1 vssd1 vccd1 vccd1 _03009_ sky130_fd_sc_hd__or3_1
Xoutput240 net240 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[10] sky130_fd_sc_hd__buf_2
XANTENNA_fanout1313_A net1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11001__D net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput251 net251 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[25] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_101_957 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput262 net262 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[9] sky130_fd_sc_hd__buf_2
XANTENNA_fanout773_A _02851_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07728__C1 net1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_2207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout394_X net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10878__A2 _05632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1101_X net1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_52_Right_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07743__A2 net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08940__A1 net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout940_A net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07969_ net1107 team_03_WB.instance_to_wrap.core.register_file.registers_state\[240\]
+ net901 vssd1 vssd1 vccd1 vccd1 _03911_ sky130_fd_sc_hd__or3_1
XANTENNA_fanout659_X net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08379__S0 net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09708_ _04150_ _04210_ _05014_ _05071_ net555 net571 vssd1 vssd1 vccd1 vccd1 _05650_
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_96_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11827__A1 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10980_ net1251 net1252 net1018 vssd1 vssd1 vccd1 vccd1 _06558_ sky130_fd_sc_hd__and3_2
XFILLER_0_69_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_104_2510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_2521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09639_ _05356_ _05577_ _05578_ _05580_ _05575_ vssd1 vssd1 vccd1 vccd1 _05581_ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout826_X net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_434 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07223__B net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12650_ net1284 vssd1 vssd1 vccd1 vccd1 _00414_ sky130_fd_sc_hd__inv_2
XFILLER_0_168_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_2429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_139_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11601_ _06527_ net2496 net449 vssd1 vssd1 vccd1 vccd1 _01928_ sky130_fd_sc_hd__mux2_1
XFILLER_0_167_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_155_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12581_ net1356 vssd1 vssd1 vccd1 vccd1 _00345_ sky130_fd_sc_hd__inv_2
XANTENNA__10865__A net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_61_Right_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_154_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14320_ clknet_leaf_161_wb_clk_i _02084_ _00685_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[674\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_93_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15078__1464 vssd1 vssd1 vccd1 vccd1 _15078__1464/HI net1464 sky130_fd_sc_hd__conb_1
X_11532_ _06430_ net643 net707 net699 vssd1 vssd1 vccd1 vccd1 _06784_ sky130_fd_sc_hd__and4_1
XANTENNA__10802__A2 net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14251_ clknet_leaf_42_wb_clk_i _02015_ _00616_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[605\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12004__A1 net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11463_ net504 net634 _06588_ net393 net1983 vssd1 vssd1 vccd1 vccd1 _02032_ sky130_fd_sc_hd__a32o_1
XFILLER_0_162_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13202_ net1398 vssd1 vssd1 vccd1 vccd1 _00966_ sky130_fd_sc_hd__inv_2
XANTENNA__09956__A0 _05882_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08759__A1 net1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10414_ _06236_ _06237_ team_03_WB.instance_to_wrap.core.pc.current_pc\[13\] net681
+ vssd1 vssd1 vccd1 vccd1 _02647_ sky130_fd_sc_hd__o2bb2a_1
X_14182_ clknet_leaf_117_wb_clk_i _01946_ _00547_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[536\]
+ sky130_fd_sc_hd__dfrtp_1
X_11394_ net508 net636 _06749_ net402 net2133 vssd1 vssd1 vccd1 vccd1 _02083_ sky130_fd_sc_hd__a32o_1
XANTENNA__09420__A2 _02804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_1977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10566__B2 _05876_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11763__B1 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_1988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07431__A1 net1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13133_ net1292 vssd1 vssd1 vccd1 vccd1 _00897_ sky130_fd_sc_hd__inv_2
X_10345_ _06110_ _06180_ vssd1 vssd1 vccd1 vccd1 _06181_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_29_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13064_ net1299 vssd1 vssd1 vccd1 vccd1 _00828_ sky130_fd_sc_hd__inv_2
X_10276_ _03822_ _06117_ vssd1 vssd1 vccd1 vccd1 _06118_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07719__C1 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_70_Right_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_167_3794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1410 net1413 vssd1 vssd1 vccd1 vccd1 net1410 sky130_fd_sc_hd__buf_4
X_12015_ _06763_ net463 net360 net2415 vssd1 vssd1 vccd1 vccd1 _01530_ sky130_fd_sc_hd__a22o_1
Xfanout1421 net1422 vssd1 vssd1 vccd1 vccd1 net1421 sky130_fd_sc_hd__buf_4
Xfanout1432 net1434 vssd1 vssd1 vccd1 vccd1 net1432 sky130_fd_sc_hd__buf_4
XFILLER_0_136_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08931__A1 net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07734__A2 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_2919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13966_ clknet_leaf_130_wb_clk_i _01730_ _00331_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[320\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10759__B _06294_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08144__C1 net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_535 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12917_ net1274 vssd1 vssd1 vccd1 vccd1 _00681_ sky130_fd_sc_hd__inv_2
XANTENNA__08695__B1 net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11294__A2 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13897_ clknet_leaf_74_wb_clk_i _01661_ _00262_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[251\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09892__C1 net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12848_ net1410 vssd1 vssd1 vccd1 vccd1 _00612_ sky130_fd_sc_hd__inv_2
XFILLER_0_57_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12779_ net1281 vssd1 vssd1 vccd1 vccd1 _00543_ sky130_fd_sc_hd__inv_2
XFILLER_0_57_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13151__A net1347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08998__A1 net1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14518_ clknet_leaf_178_wb_clk_i _02282_ _00883_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[872\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14449_ clknet_leaf_141_wb_clk_i _02213_ _00814_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[803\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_142_835 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10006__A0 _03458_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09628__X _05570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold904 team_03_WB.instance_to_wrap.core.register_file.registers_state\[651\] vssd1
+ vssd1 vccd1 vccd1 net2397 sky130_fd_sc_hd__dlygate4sd3_1
Xhold915 team_03_WB.instance_to_wrap.core.register_file.registers_state\[103\] vssd1
+ vssd1 vccd1 vccd1 net2408 sky130_fd_sc_hd__dlygate4sd3_1
Xhold926 team_03_WB.instance_to_wrap.core.register_file.registers_state\[527\] vssd1
+ vssd1 vccd1 vccd1 net2419 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11754__B1 net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold937 team_03_WB.instance_to_wrap.core.register_file.registers_state\[901\] vssd1
+ vssd1 vccd1 vccd1 net2430 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_29_wb_clk_i_A clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__07422__A1 net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold948 team_03_WB.instance_to_wrap.core.register_file.registers_state\[845\] vssd1
+ vssd1 vccd1 vccd1 net2441 sky130_fd_sc_hd__dlygate4sd3_1
X_09990_ _05875_ net1738 net290 vssd1 vssd1 vccd1 vccd1 _02724_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold959 team_03_WB.instance_to_wrap.core.register_file.registers_state\[918\] vssd1
+ vssd1 vccd1 vccd1 net2452 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_86_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08941_ net1217 _04881_ _04882_ net1071 vssd1 vssd1 vccd1 vccd1 _04883_ sky130_fd_sc_hd__o211a_1
XANTENNA__11506__A0 _06624_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_0_wb_clk_i_A wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08872_ _04808_ _04811_ _04812_ net595 vssd1 vssd1 vccd1 vccd1 _04814_ sky130_fd_sc_hd__a31o_1
XANTENNA__07186__B1 net1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07823_ net1082 team_03_WB.instance_to_wrap.core.register_file.registers_state\[74\]
+ net792 team_03_WB.instance_to_wrap.core.register_file.registers_state\[106\] net739
+ vssd1 vssd1 vccd1 vccd1 _03765_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_84_2104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10302__X _06144_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07754_ net1101 team_03_WB.instance_to_wrap.core.register_file.registers_state\[492\]
+ net898 _03695_ net1155 vssd1 vssd1 vccd1 vccd1 _03696_ sky130_fd_sc_hd__o311a_1
XANTENNA__09478__A2 _04476_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09015__S net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_149_412 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07685_ net1174 team_03_WB.instance_to_wrap.core.register_file.registers_state\[702\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[670\] net760 net728
+ vssd1 vssd1 vccd1 vccd1 _03627_ sky130_fd_sc_hd__a221o_1
XFILLER_0_17_1024 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1096_A net1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10493__B1 net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09424_ _05360_ _05365_ net553 vssd1 vssd1 vccd1 vccd1 _05366_ sky130_fd_sc_hd__mux2_1
XANTENNA__08781__S0 net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_165_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09355_ _03947_ _05148_ vssd1 vssd1 vccd1 vccd1 _05297_ sky130_fd_sc_hd__xor2_1
XFILLER_0_118_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11037__A2 net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout521_A _06395_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06882__B team_03_WB.instance_to_wrap.core.decoder.inst\[26\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1263_A net1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout619_A net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08306_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[440\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[408\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[312\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[280\]
+ net973 net1073 vssd1 vssd1 vccd1 vccd1 _04248_ sky130_fd_sc_hd__mux4_1
XANTENNA_clkbuf_leaf_68_wb_clk_i_A clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09286_ _04922_ _05225_ vssd1 vssd1 vccd1 vccd1 _05228_ sky130_fd_sc_hd__or2_1
XANTENNA__08155__A team_03_WB.instance_to_wrap.core.decoder.inst\[19\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07110__B1 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11993__A0 net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09650__A2 _05547_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_173_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08237_ net432 net427 _04178_ vssd1 vssd1 vccd1 vccd1 _04179_ sky130_fd_sc_hd__or3b_2
XFILLER_0_16_852 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1430_A net1435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_595 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1051_X net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout407_X net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_179_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_179_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_43_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1149_X net1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08168_ net1061 _04108_ _04109_ _04107_ vssd1 vssd1 vccd1 vccd1 _04110_ sky130_fd_sc_hd__o31a_1
XFILLER_0_15_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout890_A net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_108_wb_clk_i clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_108_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__11745__B1 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07949__C1 net1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout988_A net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07119_ net614 _03060_ vssd1 vssd1 vccd1 vccd1 _03061_ sky130_fd_sc_hd__nor2_1
XANTENNA__07413__A1 net1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10624__S net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08099_ _04037_ _04040_ net821 vssd1 vssd1 vccd1 vccd1 _04041_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_24_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10130_ _04415_ _02767_ net672 vssd1 vssd1 vccd1 vccd1 _05972_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_128_3008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07335__A1_N net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_73_1874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10061_ net24 net1039 net911 net2770 vssd1 vssd1 vccd1 vccd1 _02670_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_73_1885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_3344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_3355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07716__A2 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout943_X net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10720__A1 net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06924__B1 net1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13820_ clknet_leaf_149_wb_clk_i _01584_ _00185_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[174\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_98_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_162_3691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07234__A net1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13751_ clknet_leaf_115_wb_clk_i _01515_ _00116_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[105\]
+ sky130_fd_sc_hd__dfrtp_1
X_10963_ net689 _05798_ vssd1 vssd1 vccd1 vccd1 _06544_ sky130_fd_sc_hd__nand2_1
XANTENNA__11276__A2 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12702_ net1391 vssd1 vssd1 vccd1 vccd1 _00466_ sky130_fd_sc_hd__inv_2
XANTENNA__10484__B1 net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08764__S net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13682_ clknet_leaf_117_wb_clk_i _01446_ _00047_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[36\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10894_ net299 net2580 net521 vssd1 vssd1 vccd1 vccd1 _02321_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11028__A2 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12633_ net1365 vssd1 vssd1 vccd1 vccd1 _00397_ sky130_fd_sc_hd__inv_2
XFILLER_0_38_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08429__B1 net1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10236__A0 net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12564_ net1310 vssd1 vssd1 vccd1 vccd1 _00328_ sky130_fd_sc_hd__inv_2
XFILLER_0_109_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08065__A net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11984__A0 net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14303_ clknet_leaf_25_wb_clk_i _02067_ _00668_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[657\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11515_ _06630_ net2617 net391 vssd1 vssd1 vccd1 vccd1 _01991_ sky130_fd_sc_hd__mux2_1
XANTENNA__10882__X _06478_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07652__A1 net1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07400__C net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12495_ net1336 vssd1 vssd1 vccd1 vccd1 _00259_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_117_2778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14234_ clknet_leaf_142_wb_clk_i _01998_ _00599_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[588\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_44_Left_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input72_X net72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11446_ net277 net643 net707 net830 vssd1 vssd1 vccd1 vccd1 _06762_ sky130_fd_sc_hd__and4_1
XANTENNA__08352__X _04294_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11736__B1 _06808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_141_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07404__A1 net1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_169_3845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14165_ clknet_leaf_106_wb_clk_i _01929_ _00530_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[519\]
+ sky130_fd_sc_hd__dfrtp_1
X_11377_ net714 net296 net699 vssd1 vssd1 vccd1 vccd1 _06741_ sky130_fd_sc_hd__and3_1
XFILLER_0_22_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13116_ net1419 vssd1 vssd1 vccd1 vccd1 _00880_ sky130_fd_sc_hd__inv_2
X_10328_ _02767_ _06151_ vssd1 vssd1 vccd1 vccd1 _06167_ sky130_fd_sc_hd__xnor2_1
X_14096_ clknet_leaf_158_wb_clk_i _01860_ _00461_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[450\]
+ sky130_fd_sc_hd__dfrtp_1
X_13047_ net1387 vssd1 vssd1 vccd1 vccd1 _00811_ sky130_fd_sc_hd__inv_2
X_10259_ _04030_ _06099_ vssd1 vssd1 vccd1 vccd1 _06101_ sky130_fd_sc_hd__xor2_1
XANTENNA__08939__S net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09183__X _05125_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08904__A1 net1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1240 net1241 vssd1 vssd1 vccd1 vccd1 net1240 sky130_fd_sc_hd__clkbuf_4
Xfanout1251 team_03_WB.instance_to_wrap.core.decoder.inst\[8\] vssd1 vssd1 vccd1 vccd1
+ net1251 sky130_fd_sc_hd__clkbuf_4
Xfanout1262 net1263 vssd1 vssd1 vccd1 vccd1 net1262 sky130_fd_sc_hd__buf_4
Xfanout1273 net1278 vssd1 vssd1 vccd1 vccd1 net1273 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06915__B1 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1284 net1286 vssd1 vssd1 vccd1 vccd1 net1284 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_1_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_53_Left_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13146__A net1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1295 net1302 vssd1 vssd1 vccd1 vccd1 net1295 sky130_fd_sc_hd__buf_2
XFILLER_0_163_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14998_ clknet_leaf_65_wb_clk_i net46 _01363_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08117__C1 net1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13949_ clknet_leaf_26_wb_clk_i _01713_ _00314_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[303\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_102_wb_clk_i_A clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_88_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_159_743 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10475__B1 net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07470_ net1184 team_03_WB.instance_to_wrap.core.register_file.registers_state\[565\]
+ net876 vssd1 vssd1 vccd1 vccd1 _03412_ sky130_fd_sc_hd__and3_1
XFILLER_0_5_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_147_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07891__A1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_173_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09140_ _04538_ _05074_ _04779_ vssd1 vssd1 vccd1 vccd1 _05082_ sky130_fd_sc_hd__or3b_4
XANTENNA__10936__C _05845_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_6_wb_clk_i clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_6_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__11975__A0 _06405_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_62_Left_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09071_ net433 net427 net589 net550 vssd1 vssd1 vccd1 vccd1 _05013_ sky130_fd_sc_hd__o31a_1
XFILLER_0_112_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11113__B _06541_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08840__B1 net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08022_ net1177 team_03_WB.instance_to_wrap.core.register_file.registers_state\[49\]
+ net877 vssd1 vssd1 vccd1 vccd1 _03964_ sky130_fd_sc_hd__and3_1
XFILLER_0_31_118 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold701 net237 vssd1 vssd1 vccd1 vccd1 net2194 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10952__B _05768_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold712 team_03_WB.instance_to_wrap.core.register_file.registers_state\[482\] vssd1
+ vssd1 vccd1 vccd1 net2205 sky130_fd_sc_hd__dlygate4sd3_1
Xhold723 team_03_WB.instance_to_wrap.core.register_file.registers_state\[876\] vssd1
+ vssd1 vccd1 vccd1 net2216 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_343 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold734 team_03_WB.instance_to_wrap.core.register_file.registers_state\[624\] vssd1
+ vssd1 vccd1 vccd1 net2227 sky130_fd_sc_hd__dlygate4sd3_1
Xhold745 team_03_WB.instance_to_wrap.core.register_file.registers_state\[774\] vssd1
+ vssd1 vccd1 vccd1 net2238 sky130_fd_sc_hd__dlygate4sd3_1
Xhold756 team_03_WB.instance_to_wrap.core.register_file.registers_state\[520\] vssd1
+ vssd1 vccd1 vccd1 net2249 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold767 team_03_WB.instance_to_wrap.core.register_file.registers_state\[547\] vssd1
+ vssd1 vccd1 vccd1 net2260 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07319__A net1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold778 team_03_WB.instance_to_wrap.core.register_file.registers_state\[475\] vssd1
+ vssd1 vccd1 vccd1 net2271 sky130_fd_sc_hd__dlygate4sd3_1
X_09973_ _03458_ net1830 net292 vssd1 vssd1 vccd1 vccd1 _02740_ sky130_fd_sc_hd__mux2_1
Xhold789 team_03_WB.instance_to_wrap.core.register_file.registers_state\[661\] vssd1
+ vssd1 vccd1 vccd1 net2282 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11486__D net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08924_ net1241 team_03_WB.instance_to_wrap.core.register_file.registers_state\[139\]
+ net977 team_03_WB.instance_to_wrap.core.register_file.registers_state\[171\] net940
+ vssd1 vssd1 vccd1 vccd1 _04866_ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout1011_A net1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07159__B1 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08356__C1 net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_141_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout1109_A net1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_71_Left_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08855_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[544\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[512\]
+ net990 vssd1 vssd1 vccd1 vccd1 _04797_ sky130_fd_sc_hd__mux2_1
X_15077__1463 vssd1 vssd1 vccd1 vccd1 _15077__1463/HI net1463 sky130_fd_sc_hd__conb_1
XANTENNA_fanout471_A net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07980__C net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_157_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout569_A _03024_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_107 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_2_Right_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07806_ _03744_ _03747_ net818 vssd1 vssd1 vccd1 vccd1 _03748_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_58_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08786_ net1051 team_03_WB.instance_to_wrap.core.register_file.registers_state\[834\]
+ net1001 team_03_WB.instance_to_wrap.core.register_file.registers_state\[866\] net1214
+ vssd1 vssd1 vccd1 vccd1 _04728_ sky130_fd_sc_hd__a221o_1
XFILLER_0_93_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08108__C1 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_140_3241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_3252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07737_ team_03_WB.instance_to_wrap.core.decoder.inst\[13\] net1015 _03107_ vssd1
+ vssd1 vccd1 vccd1 _03679_ sky130_fd_sc_hd__a21oi_4
XANTENNA__11258__A2 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1380_A net1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout736_A net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout357_X net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1099_X net1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_49_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07668_ net1174 team_03_WB.instance_to_wrap.core.register_file.registers_state\[94\]
+ net761 team_03_WB.instance_to_wrap.core.register_file.registers_state\[126\] net725
+ vssd1 vssd1 vccd1 vccd1 _03610_ sky130_fd_sc_hd__o221a_1
XFILLER_0_95_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09407_ net547 _04237_ _04325_ vssd1 vssd1 vccd1 vccd1 _05349_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10619__S net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout524_X net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout903_A net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07599_ net1203 team_03_WB.instance_to_wrap.core.register_file.registers_state\[473\]
+ vssd1 vssd1 vccd1 vccd1 _03541_ sky130_fd_sc_hd__or2_1
XFILLER_0_36_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09338_ _05196_ _05202_ vssd1 vssd1 vccd1 vccd1 _05280_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_80_Left_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10769__A1 net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12119__B net99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11966__B1 net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07634__A1 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09269_ net591 _05210_ vssd1 vssd1 vccd1 vccd1 _05211_ sky130_fd_sc_hd__or2_1
XFILLER_0_51_917 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09859__D_N _05757_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11300_ _06609_ net2731 net404 vssd1 vssd1 vccd1 vccd1 _02145_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12280_ net1375 vssd1 vssd1 vccd1 vccd1 _00044_ sky130_fd_sc_hd__inv_2
XFILLER_0_44_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout893_X net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08809__S1 net1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_75_1914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_180_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_11231_ _06545_ net2222 net488 vssd1 vssd1 vccd1 vccd1 _02180_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_75_1925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07229__A net1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_140_1020 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11162_ net706 net271 net698 vssd1 vssd1 vccd1 vccd1 _06659_ sky130_fd_sc_hd__and3_2
XTAP_TAPCELL_ROW_112_2675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10113_ _05952_ _05953_ _05956_ vssd1 vssd1 vccd1 vccd1 _05957_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_164_3742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11093_ net833 net299 vssd1 vssd1 vccd1 vccd1 _06623_ sky130_fd_sc_hd__and2_2
XANTENNA__08347__C1 net1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input32_A DAT_I[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07516__X _03458_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10044_ net12 net1039 net911 net2776 vssd1 vssd1 vccd1 vccd1 _02687_ sky130_fd_sc_hd__a22o_1
X_14921_ clknet_leaf_43_wb_clk_i _02676_ _01286_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_O\[8\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__08898__B1 net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_76_wb_clk_i clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_76_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xhold50 team_03_WB.instance_to_wrap.core.register_file.registers_state\[977\] vssd1
+ vssd1 vccd1 vccd1 net1543 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold61 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1009\] vssd1
+ vssd1 vccd1 vccd1 net1554 sky130_fd_sc_hd__dlygate4sd3_1
Xhold72 _02623_ vssd1 vssd1 vccd1 vccd1 net1565 sky130_fd_sc_hd__dlygate4sd3_1
X_14852_ clknet_leaf_66_wb_clk_i net1853 _01217_ vssd1 vssd1 vccd1 vccd1 net107 sky130_fd_sc_hd__dfrtp_1
Xhold83 team_03_WB.instance_to_wrap.core.register_file.registers_state\[978\] vssd1
+ vssd1 vccd1 vccd1 net1576 sky130_fd_sc_hd__dlygate4sd3_1
Xhold94 team_03_WB.instance_to_wrap.ADR_I\[31\] vssd1 vssd1 vccd1 vccd1 net1587 sky130_fd_sc_hd__dlygate4sd3_1
X_13803_ clknet_leaf_38_wb_clk_i _01567_ _00168_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[157\]
+ sky130_fd_sc_hd__dfrtp_1
X_14783_ clknet_leaf_95_wb_clk_i _02547_ _01148_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_I\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10102__B net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11995_ _06754_ net466 net444 net2317 vssd1 vssd1 vccd1 vccd1 _01549_ sky130_fd_sc_hd__a22o_1
XFILLER_0_58_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11913__S net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13734_ clknet_leaf_73_wb_clk_i _01498_ _00099_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[88\]
+ sky130_fd_sc_hd__dfrtp_1
X_10946_ team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[5\] net308 net689 vssd1
+ vssd1 vccd1 vccd1 _06530_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07322__B1 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_119_Left_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13665_ clknet_leaf_181_wb_clk_i _01429_ _00030_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_10877_ net273 net2187 net518 vssd1 vssd1 vccd1 vccd1 _02324_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_155_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_119_2818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12616_ net1297 vssd1 vssd1 vccd1 vccd1 _00380_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_119_2829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13596_ net1340 vssd1 vssd1 vccd1 vccd1 _01360_ sky130_fd_sc_hd__inv_2
XFILLER_0_155_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_171_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11957__B1 net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_610 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12547_ net1356 vssd1 vssd1 vccd1 vccd1 _00311_ sky130_fd_sc_hd__inv_2
XANTENNA__11421__A2 net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_427 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08888__C_N net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11972__A3 net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_451 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12478_ net1392 vssd1 vssd1 vccd1 vccd1 _00242_ sky130_fd_sc_hd__inv_2
XANTENNA_3 team_03_WB.instance_to_wrap.core.decoder.inst\[12\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__10772__B net1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14217_ clknet_leaf_77_wb_clk_i _01981_ _00582_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[571\]
+ sky130_fd_sc_hd__dfrtp_1
X_11429_ net269 net2755 net399 vssd1 vssd1 vccd1 vccd1 _02055_ sky130_fd_sc_hd__mux2_1
XFILLER_0_112_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07389__B1 net1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11185__B2 net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14148_ clknet_leaf_29_wb_clk_i _01912_ _00513_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[502\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06970_ _02871_ _02910_ _02911_ _02869_ _02909_ vssd1 vssd1 vccd1 vccd1 _02912_ sky130_fd_sc_hd__a221o_1
X_14079_ clknet_leaf_171_wb_clk_i _01843_ _00444_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[433\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1070 net1074 vssd1 vssd1 vccd1 vccd1 net1070 sky130_fd_sc_hd__buf_4
Xfanout1081 _02788_ vssd1 vssd1 vccd1 vccd1 net1081 sky130_fd_sc_hd__buf_6
X_08640_ _04580_ _04581_ vssd1 vssd1 vccd1 vccd1 _04582_ sky130_fd_sc_hd__and2_1
XFILLER_0_174_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1092 net1093 vssd1 vssd1 vccd1 vccd1 net1092 sky130_fd_sc_hd__buf_2
XANTENNA__09641__X _05583_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08571_ net1234 team_03_WB.instance_to_wrap.core.register_file.registers_state\[349\]
+ net966 team_03_WB.instance_to_wrap.core.register_file.registers_state\[381\] net1073
+ vssd1 vssd1 vccd1 vccd1 _04513_ sky130_fd_sc_hd__o221a_1
XFILLER_0_156_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_156_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13604__A net1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07522_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[934\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[902\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[806\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[774\]
+ net778 net1134 vssd1 vssd1 vccd1 vccd1 _03464_ sky130_fd_sc_hd__mux4_1
XFILLER_0_9_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08510__C1 net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_147_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07864__A1 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07453_ net1184 team_03_WB.instance_to_wrap.core.register_file.registers_state\[181\]
+ net895 net1128 vssd1 vssd1 vccd1 vccd1 _03395_ sky130_fd_sc_hd__a211o_1
XFILLER_0_174_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11124__A net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_79_2003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07384_ net1180 team_03_WB.instance_to_wrap.core.register_file.registers_state\[479\]
+ net758 team_03_WB.instance_to_wrap.core.register_file.registers_state\[511\] net1149
+ vssd1 vssd1 vccd1 vccd1 _03326_ sky130_fd_sc_hd__o221a_1
XFILLER_0_9_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_44_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11948__B1 net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_44_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08136__C _03428_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09123_ _05061_ _05062_ _05063_ _05064_ net862 net924 vssd1 vssd1 vccd1 vccd1 _05065_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_45_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout317_A net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1059_A net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_96_2350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09054_ net1219 _04993_ _04994_ vssd1 vssd1 vccd1 vccd1 _04996_ sky130_fd_sc_hd__and3_1
XFILLER_0_103_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11963__A3 net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08433__A net1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_624 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08005_ _03945_ _03946_ vssd1 vssd1 vccd1 vccd1 _03947_ sky130_fd_sc_hd__or2_2
XFILLER_0_4_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold520 team_03_WB.instance_to_wrap.core.register_file.registers_state\[377\] vssd1
+ vssd1 vccd1 vccd1 net2013 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold531 team_03_WB.instance_to_wrap.core.register_file.registers_state\[281\] vssd1
+ vssd1 vccd1 vccd1 net2024 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_2258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1226_A net1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold542 team_03_WB.instance_to_wrap.core.register_file.registers_state\[431\] vssd1
+ vssd1 vccd1 vccd1 net2035 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_2269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08577__C1 net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07919__A2 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold553 team_03_WB.instance_to_wrap.core.register_file.registers_state\[179\] vssd1
+ vssd1 vccd1 vccd1 net2046 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08041__A1 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold564 team_03_WB.instance_to_wrap.core.register_file.registers_state\[299\] vssd1
+ vssd1 vccd1 vccd1 net2057 sky130_fd_sc_hd__dlygate4sd3_1
Xhold575 team_03_WB.instance_to_wrap.core.register_file.registers_state\[101\] vssd1
+ vssd1 vccd1 vccd1 net2068 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10923__A1 net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold586 team_03_WB.instance_to_wrap.core.register_file.registers_state\[747\] vssd1
+ vssd1 vccd1 vccd1 net2079 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout686_A net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold597 team_03_WB.instance_to_wrap.core.register_file.registers_state\[332\] vssd1
+ vssd1 vccd1 vccd1 net2090 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_70_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09956_ _05882_ net1647 net291 vssd1 vssd1 vccd1 vccd1 _02749_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_70_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1014_X net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07336__X _03278_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08907_ net1239 team_03_WB.instance_to_wrap.core.register_file.registers_state\[716\]
+ net981 team_03_WB.instance_to_wrap.core.register_file.registers_state\[748\] net942
+ vssd1 vssd1 vccd1 vccd1 _04849_ sky130_fd_sc_hd__o221a_1
X_09887_ _03137_ _04148_ _05828_ vssd1 vssd1 vccd1 vccd1 _05829_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11479__A2 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout853_A _04096_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1220 team_03_WB.instance_to_wrap.core.register_file.registers_state\[722\] vssd1
+ vssd1 vccd1 vccd1 net2713 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1231 team_03_WB.instance_to_wrap.core.register_file.registers_state\[204\] vssd1
+ vssd1 vccd1 vccd1 net2724 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10687__B1 net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08838_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[32\] net994
+ vssd1 vssd1 vccd1 vccd1 _04780_ sky130_fd_sc_hd__or2_1
Xhold1242 team_03_WB.instance_to_wrap.core.register_file.registers_state\[656\] vssd1
+ vssd1 vccd1 vccd1 net2735 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_142_Right_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1253 team_03_WB.instance_to_wrap.core.register_file.registers_state\[588\] vssd1
+ vssd1 vccd1 vccd1 net2746 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1264 team_03_WB.instance_to_wrap.core.register_file.registers_state\[327\] vssd1
+ vssd1 vccd1 vccd1 net2757 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1275 team_03_WB.instance_to_wrap.CPU_DAT_O\[12\] vssd1 vssd1 vccd1 vccd1 net2768
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1286 team_03_WB.instance_to_wrap.core.register_file.registers_state\[704\] vssd1
+ vssd1 vccd1 vccd1 net2779 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout641_X net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08769_ net852 _04693_ _04702_ _04710_ vssd1 vssd1 vccd1 vccd1 _04711_ sky130_fd_sc_hd__a2bb2o_4
XANTENNA__11733__S net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout739_X net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10439__B1 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10800_ _06406_ _06408_ net585 vssd1 vssd1 vccd1 vccd1 _06409_ sky130_fd_sc_hd__o21a_2
XTAP_TAPCELL_ROW_68_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1057 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11780_ net2764 _06613_ net327 vssd1 vssd1 vccd1 vccd1 _01758_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_4_3__f_wb_clk_i_A clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10731_ net1743 net528 net523 _06357_ vssd1 vssd1 vccd1 vccd1 _02450_ sky130_fd_sc_hd__a22o_1
XANTENNA__07855__A1 net1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout906_X net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13450_ net1405 vssd1 vssd1 vccd1 vccd1 _01214_ sky130_fd_sc_hd__inv_2
XFILLER_0_165_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_24_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10662_ net1143 net1495 vssd1 vssd1 vccd1 vccd1 _02466_ sky130_fd_sc_hd__or2_1
XFILLER_0_12_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09057__B1 net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_157_3590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_204 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_123_wb_clk_i clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_123_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_12401_ net1267 vssd1 vssd1 vccd1 vccd1 _00165_ sky130_fd_sc_hd__inv_2
XFILLER_0_119_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07607__A1 net1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13381_ net1432 vssd1 vssd1 vccd1 vccd1 _01145_ sky130_fd_sc_hd__inv_2
XANTENNA__08804__B1 net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10593_ team_03_WB.instance_to_wrap.core.ru.prev_busy _06281_ vssd1 vssd1 vccd1 vccd1
+ _06302_ sky130_fd_sc_hd__nand2_1
XFILLER_0_152_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15120_ net913 vssd1 vssd1 vccd1 vccd1 net251 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_69_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12332_ net1311 vssd1 vssd1 vccd1 vccd1 _00096_ sky130_fd_sc_hd__inv_2
XANTENNA__07083__A2 _03023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_114_2715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11954__A3 net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08280__A1 net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_2726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15051_ net1492 vssd1 vssd1 vccd1 vccd1 gpio_oeb[3] sky130_fd_sc_hd__buf_2
XFILLER_0_32_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12263_ net1368 vssd1 vssd1 vccd1 vccd1 _00027_ sky130_fd_sc_hd__inv_2
X_14002_ clknet_leaf_165_wb_clk_i _01766_ _00367_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[356\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08568__C1 net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11214_ net2268 net486 _06681_ net495 vssd1 vssd1 vccd1 vccd1 _02195_ sky130_fd_sc_hd__a22o_1
XFILLER_0_31_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08032__A1 net1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12194_ net1530 vssd1 vssd1 vccd1 vccd1 _02359_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_120_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09445__Y _05387_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07240__C1 net1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11145_ net2081 net413 _06649_ net497 vssd1 vssd1 vccd1 vccd1 _02232_ sky130_fd_sc_hd__a22o_1
XFILLER_0_101_370 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08489__S net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10812__S net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10390__A2 net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07393__S net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11076_ net834 net277 vssd1 vssd1 vccd1 vccd1 _06616_ sky130_fd_sc_hd__and2_2
X_10027_ net1143 net100 _05903_ vssd1 vssd1 vccd1 vccd1 _02700_ sky130_fd_sc_hd__mux2_1
X_14904_ clknet_leaf_86_wb_clk_i _02667_ _01269_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.pc.current_pc\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07543__B1 net1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09902__A _05563_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14835_ clknet_leaf_89_wb_clk_i net1877 _01200_ vssd1 vssd1 vccd1 vccd1 net156 sky130_fd_sc_hd__dfrtp_1
XANTENNA__07125__C net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_127_Left_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08718__S0 net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14766_ clknet_leaf_44_wb_clk_i net1709 _01131_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_11978_ net279 net2634 net443 vssd1 vssd1 vccd1 vccd1 _01566_ sky130_fd_sc_hd__mux2_1
XANTENNA__10767__B net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09113__S net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_666 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10929_ net314 _05846_ _05928_ team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[8\]
+ vssd1 vssd1 vccd1 vccd1 _06516_ sky130_fd_sc_hd__or4b_1
XFILLER_0_129_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13717_ clknet_leaf_129_wb_clk_i _01481_ _00082_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[71\]
+ sky130_fd_sc_hd__dfrtp_1
X_14697_ clknet_leaf_60_wb_clk_i _02461_ _01062_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.ADR_I\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_129_746 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11642__A2 net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09048__B1 net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13648_ clknet_leaf_159_wb_clk_i _01412_ _00013_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_156_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_627 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09599__A1 net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13579_ net1426 vssd1 vssd1 vccd1 vccd1 _01343_ sky130_fd_sc_hd__inv_2
XANTENNA__06980__B _02893_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15076__1462 vssd1 vssd1 vccd1 vccd1 _15076__1462/HI net1462 sky130_fd_sc_hd__conb_1
XFILLER_0_42_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11945__A3 net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08271__A1 net1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08271__B2 net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_136_Left_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_169_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_10_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11158__A1 net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08559__C1 net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_55 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08023__A1 net1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_99_Right_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09220__B1 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10905__A1 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09810_ _02923_ _04565_ net537 _05751_ vssd1 vssd1 vccd1 vccd1 _05752_ sky130_fd_sc_hd__o31a_1
Xfanout307 _06396_ vssd1 vssd1 vccd1 vccd1 net307 sky130_fd_sc_hd__buf_4
Xfanout318 _05927_ vssd1 vssd1 vccd1 vccd1 net318 sky130_fd_sc_hd__clkbuf_4
Xfanout329 _06810_ vssd1 vssd1 vccd1 vccd1 net329 sky130_fd_sc_hd__buf_8
X_09741_ _05086_ _05117_ _05119_ _05110_ net555 net570 vssd1 vssd1 vccd1 vccd1 _05683_
+ sky130_fd_sc_hd__mux4_1
X_06953_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[37\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[5\]
+ net787 vssd1 vssd1 vccd1 vccd1 _02895_ sky130_fd_sc_hd__mux2_1
XANTENNA__08326__A2 net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09672_ net575 _05613_ vssd1 vssd1 vccd1 vccd1 _05614_ sky130_fd_sc_hd__and2_1
XFILLER_0_118_61 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06884_ team_03_WB.instance_to_wrap.core.decoder.inst\[30\] team_03_WB.instance_to_wrap.core.decoder.inst\[28\]
+ team_03_WB.instance_to_wrap.core.decoder.inst\[27\] _02824_ vssd1 vssd1 vccd1 vccd1
+ _02826_ sky130_fd_sc_hd__or4_1
XANTENNA__06995__X _02937_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10023__A net91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07534__B1 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_145_Left_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08731__C1 net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08623_ net853 _04564_ _04551_ vssd1 vssd1 vccd1 vccd1 _04565_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_96_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout267_A _06550_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08554_ net859 _04492_ _04495_ vssd1 vssd1 vccd1 vccd1 _04496_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_46_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11094__A0 _06623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07505_ net1110 team_03_WB.instance_to_wrap.core.register_file.registers_state\[71\]
+ net803 team_03_WB.instance_to_wrap.core.register_file.registers_state\[103\] net752
+ vssd1 vssd1 vccd1 vccd1 _03447_ sky130_fd_sc_hd__a221o_1
X_08485_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[891\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[859\]
+ net986 vssd1 vssd1 vccd1 vccd1 _04427_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_368 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11633__A2 net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout434_A net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09958__S net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1176_A net1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07436_ _03375_ _03377_ net811 vssd1 vssd1 vccd1 vccd1 _03378_ sky130_fd_sc_hd__a21o_1
XFILLER_0_91_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_63_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_232 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_3140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_hold1284_A team_03_WB.instance_to_wrap.CPU_DAT_O\[9\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_3151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout601_A _06299_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07367_ net1124 _03308_ _03307_ net1138 vssd1 vssd1 vccd1 vccd1 _03309_ sky130_fd_sc_hd__a211o_1
XFILLER_0_162_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_799 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_94_2309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09106_ net1051 team_03_WB.instance_to_wrap.core.register_file.registers_state\[206\]
+ net1001 team_03_WB.instance_to_wrap.core.register_file.registers_state\[238\] net924
+ vssd1 vssd1 vccd1 vccd1 _05048_ sky130_fd_sc_hd__a221o_1
XANTENNA__09259__A net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07298_ net819 _03239_ net719 vssd1 vssd1 vccd1 vccd1 _03240_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_14_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_3059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09037_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[944\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[912\]
+ net988 vssd1 vssd1 vccd1 vccd1 _04979_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10980__X _06558_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1131_X net1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11149__A1 net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1229_X net1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold350 team_03_WB.instance_to_wrap.core.register_file.registers_state\[53\] vssd1
+ vssd1 vccd1 vccd1 net1843 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold361 net214 vssd1 vssd1 vccd1 vccd1 net1854 sky130_fd_sc_hd__dlygate4sd3_1
Xhold372 net232 vssd1 vssd1 vccd1 vccd1 net1865 sky130_fd_sc_hd__dlygate4sd3_1
Xhold383 team_03_WB.instance_to_wrap.CPU_DAT_I\[28\] vssd1 vssd1 vccd1 vccd1 net1876
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11728__S net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10632__S net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold394 team_03_WB.instance_to_wrap.core.register_file.registers_state\[612\] vssd1
+ vssd1 vccd1 vccd1 net1887 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08610__B net992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout830 net831 vssd1 vssd1 vccd1 vccd1 net830 sky130_fd_sc_hd__buf_4
Xfanout841 _06304_ vssd1 vssd1 vccd1 vccd1 net841 sky130_fd_sc_hd__buf_4
XANTENNA__08970__C1 net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout852 _04096_ vssd1 vssd1 vccd1 vccd1 net852 sky130_fd_sc_hd__buf_6
XANTENNA__07507__A net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10109__C1 _03060_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09939_ _03526_ net662 vssd1 vssd1 vccd1 vccd1 _05874_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout856_X net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout863 net866 vssd1 vssd1 vccd1 vccd1 net863 sky130_fd_sc_hd__clkbuf_4
Xfanout874 net875 vssd1 vssd1 vccd1 vccd1 net874 sky130_fd_sc_hd__buf_4
XANTENNA__11029__A net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout885 net886 vssd1 vssd1 vccd1 vccd1 net885 sky130_fd_sc_hd__clkbuf_4
X_12950_ net1280 vssd1 vssd1 vccd1 vccd1 _00714_ sky130_fd_sc_hd__inv_2
Xfanout896 net900 vssd1 vssd1 vccd1 vccd1 net896 sky130_fd_sc_hd__buf_2
Xhold1050 team_03_WB.instance_to_wrap.core.register_file.registers_state\[131\] vssd1
+ vssd1 vccd1 vccd1 net2543 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07525__B1 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1061 team_03_WB.instance_to_wrap.core.register_file.registers_state\[147\] vssd1
+ vssd1 vccd1 vccd1 net2554 sky130_fd_sc_hd__dlygate4sd3_1
X_11901_ net637 _06710_ net470 net373 net2289 vssd1 vssd1 vccd1 vccd1 _01640_ sky130_fd_sc_hd__a32o_1
Xhold1072 team_03_WB.instance_to_wrap.core.register_file.registers_state\[671\] vssd1
+ vssd1 vccd1 vccd1 net2565 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1083 team_03_WB.instance_to_wrap.core.register_file.registers_state\[669\] vssd1
+ vssd1 vccd1 vccd1 net2576 sky130_fd_sc_hd__dlygate4sd3_1
X_12881_ net1268 vssd1 vssd1 vccd1 vccd1 _00645_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_419 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1094 team_03_WB.instance_to_wrap.core.register_file.registers_state\[105\] vssd1
+ vssd1 vccd1 vccd1 net2587 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_107_2574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13244__A net1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11832_ _06668_ net476 net326 net1913 vssd1 vssd1 vccd1 vccd1 _01707_ sky130_fd_sc_hd__a22o_1
X_14620_ clknet_leaf_151_wb_clk_i _02384_ _00985_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[974\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_29_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_159_3630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_178 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_159_3641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09817__A2 _04679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07242__A net1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14551_ clknet_leaf_80_wb_clk_i _02315_ _00916_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[905\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07828__A1 net1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07289__C1 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11763_ _06592_ net468 net333 net2008 vssd1 vssd1 vccd1 vccd1 _01774_ sky130_fd_sc_hd__a22o_1
XFILLER_0_36_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11624__A2 net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10832__A0 _06434_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10714_ net1628 net528 net522 _06347_ vssd1 vssd1 vccd1 vccd1 _02457_ sky130_fd_sc_hd__a22o_1
XFILLER_0_165_340 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13502_ net1328 vssd1 vssd1 vccd1 vccd1 _01266_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_155_3549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14482_ clknet_leaf_161_wb_clk_i _02246_ _00847_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[836\]
+ sky130_fd_sc_hd__dfrtp_1
X_11694_ _06736_ net383 net340 net1988 vssd1 vssd1 vccd1 vccd1 _01840_ sky130_fd_sc_hd__a22o_1
XFILLER_0_153_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_727 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13433_ net1433 vssd1 vssd1 vccd1 vccd1 _01197_ sky130_fd_sc_hd__inv_2
X_10645_ net1220 team_03_WB.instance_to_wrap.CPU_DAT_O\[16\] net845 vssd1 vssd1 vccd1
+ vccd1 _02483_ sky130_fd_sc_hd__mux2_1
XANTENNA__10807__S net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11388__A1 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_172_3896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13364_ net1319 vssd1 vssd1 vccd1 vccd1 _01128_ sky130_fd_sc_hd__inv_2
XANTENNA__08253__A1 net1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10576_ net1821 net532 net599 _05886_ vssd1 vssd1 vccd1 vccd1 _02547_ sky130_fd_sc_hd__a22o_1
XFILLER_0_107_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_544 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15103_ net1483 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[8] sky130_fd_sc_hd__buf_2
X_12315_ net1362 vssd1 vssd1 vccd1 vccd1 _00079_ sky130_fd_sc_hd__inv_2
XANTENNA__07461__C1 net1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13295_ net1341 vssd1 vssd1 vccd1 vccd1 _01059_ sky130_fd_sc_hd__inv_2
XFILLER_0_107_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15034_ clknet_leaf_94_wb_clk_i _02754_ _01399_ vssd1 vssd1 vccd1 vccd1 net190 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_32_780 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12246_ net1772 vssd1 vssd1 vccd1 vccd1 _01411_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_91_wb_clk_i clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_91_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__09753__A1 net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10899__A0 net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12177_ net1778 vssd1 vssd1 vccd1 vccd1 _02376_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_20_wb_clk_i clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_20_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08961__C1 net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11560__B2 net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11128_ net2116 net412 _06639_ net499 vssd1 vssd1 vccd1 vccd1 _02239_ sky130_fd_sc_hd__a22o_1
XANTENNA__07417__A net1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11059_ net655 net705 net267 net829 vssd1 vssd1 vccd1 vccd1 _06607_ sky130_fd_sc_hd__and4_1
XANTENNA__10115__A2 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08713__C1 net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06975__B net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14818_ clknet_leaf_95_wb_clk_i net1755 _01183_ vssd1 vssd1 vccd1 vccd1 net138 sky130_fd_sc_hd__dfrtp_2
XFILLER_0_171_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09808__A2 _04565_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07152__A net1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14749_ clknet_leaf_68_wb_clk_i _02513_ _01114_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_129_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11615__A2 net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12993__A net1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08270_ net937 _04211_ vssd1 vssd1 vccd1 vccd1 _04212_ sky130_fd_sc_hd__or2_1
XFILLER_0_144_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06991__A net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08492__A1 net1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14981__Q team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[0\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07221_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[914\] net791
+ vssd1 vssd1 vccd1 vccd1 _03163_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_15_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_4_2__f_wb_clk_i_X clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_15_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_83 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_10 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_719 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07152_ net1109 team_03_WB.instance_to_wrap.core.register_file.registers_state\[448\]
+ vssd1 vssd1 vccd1 vccd1 _03094_ sky130_fd_sc_hd__and2_1
XFILLER_0_42_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11121__B net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07083_ net614 _03023_ _02995_ vssd1 vssd1 vccd1 vccd1 _03025_ sky130_fd_sc_hd__a21o_1
XFILLER_0_120_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_160_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_1132 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09744__A1 net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11000__B1 net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11551__B2 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07985_ net1201 team_03_WB.instance_to_wrap.core.register_file.registers_state\[848\]
+ vssd1 vssd1 vccd1 vccd1 _03927_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout384_A net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09724_ _04816_ _05665_ net666 vssd1 vssd1 vccd1 vccd1 _05666_ sky130_fd_sc_hd__o21a_1
X_06936_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[676\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[644\]
+ net781 vssd1 vssd1 vccd1 vccd1 _02878_ sky130_fd_sc_hd__mux2_1
XANTENNA__08857__S net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_2157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09655_ _05278_ _05281_ _05300_ vssd1 vssd1 vccd1 vccd1 _05597_ sky130_fd_sc_hd__a21o_2
XFILLER_0_9_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06867_ team_03_WB.instance_to_wrap.core.control_logic.instruction\[4\] _02807_ team_03_WB.instance_to_wrap.core.control_logic.instruction\[5\]
+ vssd1 vssd1 vccd1 vccd1 _02809_ sky130_fd_sc_hd__or3b_2
XANTENNA_fanout551_A net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08606_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[997\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[965\]
+ net993 vssd1 vssd1 vccd1 vccd1 _04548_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout649_A net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09586_ _04071_ _04382_ vssd1 vssd1 vccd1 vccd1 _05528_ sky130_fd_sc_hd__or2_1
XFILLER_0_139_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_26_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08158__S1 net1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08537_ net1234 team_03_WB.instance_to_wrap.core.register_file.registers_state\[990\]
+ net965 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1022\] net1212
+ vssd1 vssd1 vccd1 vccd1 _04479_ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout1081_X net1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout437_X net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1179_X net1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_2471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07286__A2 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11015__C net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08468_ net1226 team_03_WB.instance_to_wrap.core.register_file.registers_state\[476\]
+ net951 team_03_WB.instance_to_wrap.core.register_file.registers_state\[508\] net1210
+ vssd1 vssd1 vccd1 vccd1 _04410_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_61_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07419_ net741 _03357_ _03358_ _03359_ _03360_ vssd1 vssd1 vccd1 vccd1 _03361_ sky130_fd_sc_hd__o32a_1
XFILLER_0_64_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10290__B2 net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout604_X net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10627__S net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08399_ net1245 team_03_WB.instance_to_wrap.core.register_file.registers_state\[601\]
+ net992 team_03_WB.instance_to_wrap.core.register_file.registers_state\[633\] net931
+ vssd1 vssd1 vccd1 vccd1 _04341_ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout1346_X net1346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10430_ team_03_WB.instance_to_wrap.core.pc.current_pc\[9\] _06137_ vssd1 vssd1 vccd1
+ vccd1 _06250_ sky130_fd_sc_hd__nor2_1
XFILLER_0_162_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1020 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12031__A2 net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_150_3446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_150_3457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10042__A1 net15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10361_ net304 net303 _06188_ _06193_ vssd1 vssd1 vccd1 vccd1 _06194_ sky130_fd_sc_hd__a211o_1
XFILLER_0_115_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12100_ net644 _06674_ net479 net442 net1905 vssd1 vssd1 vccd1 vccd1 _01447_ sky130_fd_sc_hd__a32o_1
XANTENNA__07994__B1 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13080_ net1379 vssd1 vssd1 vccd1 vccd1 _00844_ sky130_fd_sc_hd__inv_2
X_10292_ team_03_WB.instance_to_wrap.core.pc.current_pc\[3\] team_03_WB.instance_to_wrap.core.pc.current_pc\[2\]
+ vssd1 vssd1 vccd1 vccd1 _06134_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout973_X net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12031_ _06772_ net454 net359 net2292 vssd1 vssd1 vccd1 vccd1 _01514_ sky130_fd_sc_hd__a22o_1
Xhold180 team_03_WB.instance_to_wrap.ADR_I\[11\] vssd1 vssd1 vccd1 vccd1 net1673 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10215__X _06057_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold191 team_03_WB.instance_to_wrap.CPU_DAT_I\[16\] vssd1 vssd1 vccd1 vccd1 net1684
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07746__B1 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11542__A1 net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08943__C1 net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_2614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout660 _05950_ vssd1 vssd1 vccd1 vccd1 net660 sky130_fd_sc_hd__clkbuf_4
Xfanout671 _06563_ vssd1 vssd1 vccd1 vccd1 net671 sky130_fd_sc_hd__buf_2
Xfanout682 _05915_ vssd1 vssd1 vccd1 vccd1 net682 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12098__A2 net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout693 _02839_ vssd1 vssd1 vccd1 vccd1 net693 sky130_fd_sc_hd__clkbuf_4
X_13982_ clknet_leaf_120_wb_clk_i _01746_ _00347_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[336\]
+ sky130_fd_sc_hd__dfrtp_1
X_15075__1461 vssd1 vssd1 vccd1 vccd1 _15075__1461/HI net1461 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_126_2961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12933_ net1355 vssd1 vssd1 vccd1 vccd1 _00697_ sky130_fd_sc_hd__inv_2
XFILLER_0_88_717 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_126_2972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08171__B1 net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08710__A2 net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12864_ net1401 vssd1 vssd1 vccd1 vccd1 _00628_ sky130_fd_sc_hd__inv_2
X_14603_ clknet_leaf_45_wb_clk_i _02367_ _00968_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[957\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__11058__B1 net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11815_ net649 _06643_ net460 net323 net1724 vssd1 vssd1 vccd1 vccd1 _01724_ sky130_fd_sc_hd__a32o_1
XFILLER_0_84_912 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10885__X _06480_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12795_ net1360 vssd1 vssd1 vccd1 vccd1 _00559_ sky130_fd_sc_hd__inv_2
XFILLER_0_69_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10110__B net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11921__S net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_174_3947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14534_ clknet_leaf_71_wb_clk_i _02298_ _00899_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[888\]
+ sky130_fd_sc_hd__dfrtp_1
X_11746_ _06568_ net458 net331 net2192 vssd1 vssd1 vccd1 vccd1 _01791_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_174_3958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_174_3969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_153_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_12_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11677_ _06719_ net379 net338 net2122 vssd1 vssd1 vccd1 vccd1 _01857_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_12_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14465_ clknet_leaf_181_wb_clk_i _02229_ _00830_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[819\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_50_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13416_ net1420 vssd1 vssd1 vccd1 vccd1 _01180_ sky130_fd_sc_hd__inv_2
X_10628_ net2349 team_03_WB.instance_to_wrap.CPU_DAT_O\[1\] net843 vssd1 vssd1 vccd1
+ vccd1 _02500_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_928 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08226__A1 net1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_516 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14396_ clknet_leaf_149_wb_clk_i _02160_ _00761_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[750\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12022__A2 net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_1120 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11230__A0 net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13347_ net1335 vssd1 vssd1 vccd1 vccd1 _01111_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10559_ net1855 net533 net600 _05869_ vssd1 vssd1 vccd1 vccd1 _02564_ sky130_fd_sc_hd__a22o_1
XFILLER_0_12_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_19_wb_clk_i_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__10584__A2 net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13278_ net1406 vssd1 vssd1 vccd1 vccd1 _01042_ sky130_fd_sc_hd__inv_2
XFILLER_0_122_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09726__A1 net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09726__B2 _04820_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15017_ clknet_leaf_101_wb_clk_i _02737_ _01382_ vssd1 vssd1 vccd1 vccd1 net204 sky130_fd_sc_hd__dfrtp_1
X_12229_ net1586 vssd1 vssd1 vccd1 vccd1 _01428_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_166_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11533__B2 net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07832__S0 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07770_ net1194 team_03_WB.instance_to_wrap.core.register_file.registers_state\[972\]
+ net780 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1004\] net1165
+ vssd1 vssd1 vccd1 vccd1 _03712_ sky130_fd_sc_hd__o221a_1
XANTENNA__08677__S net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06960__A1 net1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14976__Q net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1102 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09440_ net551 _04712_ _04740_ vssd1 vssd1 vccd1 vccd1 _05382_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_82_2054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09371_ _04382_ _05312_ vssd1 vssd1 vccd1 vccd1 _05313_ sky130_fd_sc_hd__nor2_1
XFILLER_0_148_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11116__B _06550_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_2065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10795__X _06405_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07313__C net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08322_ _04253_ _04254_ net864 vssd1 vssd1 vccd1 vccd1 _04264_ sky130_fd_sc_hd__o21a_1
XFILLER_0_129_351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_58_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__08265__X _04207_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_978 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08253_ net1226 team_03_WB.instance_to_wrap.core.register_file.registers_state\[722\]
+ net950 team_03_WB.instance_to_wrap.core.register_file.registers_state\[754\] net934
+ vssd1 vssd1 vccd1 vccd1 _04195_ sky130_fd_sc_hd__o221a_1
XANTENNA__07673__C1 net1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11132__A net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07204_ net811 _03142_ _03145_ vssd1 vssd1 vccd1 vccd1 _03146_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_55_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08217__A1 net1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08184_ net1231 team_03_WB.instance_to_wrap.core.register_file.registers_state\[211\]
+ net958 team_03_WB.instance_to_wrap.core.register_file.registers_state\[243\] net935
+ vssd1 vssd1 vccd1 vccd1 _04126_ sky130_fd_sc_hd__o221a_1
XFILLER_0_160_836 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07135_ net1121 _03076_ vssd1 vssd1 vccd1 vccd1 _03077_ sky130_fd_sc_hd__nand2_1
XFILLER_0_160_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1041_A _02871_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1139_A net1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10575__A2 net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_240 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07066_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[162\] net778
+ net749 _03007_ vssd1 vssd1 vccd1 vccd1 _03008_ sky130_fd_sc_hd__o211a_1
Xoutput230 net230 vssd1 vssd1 vccd1 vccd1 gpio_out[33] sky130_fd_sc_hd__clkbuf_4
XANTENNA__08441__A _04382_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_994 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput241 net241 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[11] sky130_fd_sc_hd__buf_2
XFILLER_0_140_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput252 net252 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[26] sky130_fd_sc_hd__buf_2
XANTENNA__13059__A net1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_969 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07728__B1 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1306_A net1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_2208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12898__A net1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout387_X net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout766_A net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08587__S net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07968_ net1193 team_03_WB.instance_to_wrap.core.register_file.registers_state\[80\]
+ net786 team_03_WB.instance_to_wrap.core.register_file.registers_state\[112\] net734
+ vssd1 vssd1 vccd1 vccd1 _03910_ sky130_fd_sc_hd__o221a_1
X_09707_ _05209_ _05211_ _05276_ net595 vssd1 vssd1 vccd1 vccd1 _05649_ sky130_fd_sc_hd__a31o_1
X_06919_ net813 _02859_ _02860_ vssd1 vssd1 vccd1 vccd1 _02861_ sky130_fd_sc_hd__and3_1
XANTENNA__08379__S1 net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11288__B1 net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout554_X net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_97_wb_clk_i_A clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout933_A net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07899_ net1187 team_03_WB.instance_to_wrap.core.register_file.registers_state\[303\]
+ net877 _02872_ vssd1 vssd1 vccd1 vccd1 _03841_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout1296_X net1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_2511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_2522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09638_ net564 _05579_ net321 vssd1 vssd1 vccd1 vccd1 _05580_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_97_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09569_ _03904_ _04235_ _04820_ net1020 net1148 vssd1 vssd1 vccd1 vccd1 _05511_ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout721_X net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout819_X net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11741__S net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11600_ net295 net2279 net450 vssd1 vssd1 vccd1 vccd1 _01929_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08456__A1 net1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12580_ net1382 vssd1 vssd1 vccd1 vccd1 _00344_ sky130_fd_sc_hd__inv_2
XFILLER_0_148_671 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10799__C1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_146 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10865__B net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11531_ net497 net626 _06643_ net483 net1841 vssd1 vssd1 vccd1 vccd1 _01980_ sky130_fd_sc_hd__a32o_1
XFILLER_0_81_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11460__B1 net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10802__A3 net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14250_ clknet_leaf_7_wb_clk_i _02014_ _00615_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[604\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08208__A1 net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11462_ net2514 net395 _06767_ net501 vssd1 vssd1 vccd1 vccd1 _02033_ sky130_fd_sc_hd__a22o_1
XANTENNA__09405__B1 net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12004__A2 _06756_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13201_ net1268 vssd1 vssd1 vccd1 vccd1 _00965_ sky130_fd_sc_hd__inv_2
X_10413_ net284 _06141_ _06233_ net680 vssd1 vssd1 vccd1 vccd1 _06237_ sky130_fd_sc_hd__o31a_1
XFILLER_0_34_886 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14181_ clknet_leaf_37_wb_clk_i _01945_ _00546_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[535\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11393_ net712 net267 net697 vssd1 vssd1 vccd1 vccd1 _06749_ sky130_fd_sc_hd__and3_1
XANTENNA__10566__A2 net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13132_ net1313 vssd1 vssd1 vccd1 vccd1 _00896_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_78_1978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input62_A gpio_in[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10344_ _05975_ _05977_ vssd1 vssd1 vccd1 vccd1 _06180_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_78_1989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_1040 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13063_ net1369 vssd1 vssd1 vccd1 vccd1 _00827_ sky130_fd_sc_hd__inv_2
XFILLER_0_104_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10275_ _04444_ _02768_ net673 vssd1 vssd1 vccd1 vccd1 _06117_ sky130_fd_sc_hd__mux2_1
Xfanout1400 net1401 vssd1 vssd1 vccd1 vccd1 net1400 sky130_fd_sc_hd__buf_4
X_12014_ _06762_ net478 net362 net2604 vssd1 vssd1 vccd1 vccd1 _01531_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_167_3795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09734__X _05676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1411 net1412 vssd1 vssd1 vccd1 vccd1 net1411 sky130_fd_sc_hd__buf_4
Xfanout1422 net1436 vssd1 vssd1 vccd1 vccd1 net1422 sky130_fd_sc_hd__buf_2
XANTENNA__07195__A1 _03136_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1433 net1434 vssd1 vssd1 vccd1 vccd1 net1433 sky130_fd_sc_hd__buf_4
XANTENNA__10105__B net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11916__S net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout490 net492 vssd1 vssd1 vccd1 vccd1 net490 sky130_fd_sc_hd__clkbuf_4
X_13965_ clknet_leaf_187_wb_clk_i _01729_ _00330_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[319\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11818__A2 net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12916_ net1313 vssd1 vssd1 vccd1 vccd1 _00680_ sky130_fd_sc_hd__inv_2
XFILLER_0_88_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08695__A1 net1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13896_ clknet_leaf_8_wb_clk_i _01660_ _00261_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[250\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_17_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_100_Left_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09910__A net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12847_ net1336 vssd1 vssd1 vccd1 vccd1 _00611_ sky130_fd_sc_hd__inv_2
XFILLER_0_111_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_271 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11651__S net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_139_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12778_ net1279 vssd1 vssd1 vccd1 vccd1 _00542_ sky130_fd_sc_hd__inv_2
XANTENNA__09121__S net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14517_ clknet_leaf_105_wb_clk_i _02281_ _00882_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[871\]
+ sky130_fd_sc_hd__dfrtp_1
X_11729_ net2451 net298 net336 vssd1 vssd1 vccd1 vccd1 _01807_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_142_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_302 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14448_ clknet_leaf_161_wb_clk_i _02212_ _00813_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[802\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_142_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11203__A0 net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14379_ clknet_leaf_43_wb_clk_i _02143_ _00744_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[733\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold905 team_03_WB.instance_to_wrap.core.register_file.registers_state\[228\] vssd1
+ vssd1 vccd1 vccd1 net2398 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10557__A2 net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold916 team_03_WB.instance_to_wrap.core.register_file.registers_state\[321\] vssd1
+ vssd1 vccd1 vccd1 net2409 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11754__A1 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold927 team_03_WB.instance_to_wrap.core.register_file.registers_state\[793\] vssd1
+ vssd1 vccd1 vccd1 net2420 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09357__A net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold938 team_03_WB.instance_to_wrap.core.register_file.registers_state\[551\] vssd1
+ vssd1 vccd1 vccd1 net2431 sky130_fd_sc_hd__dlygate4sd3_1
Xhold949 team_03_WB.instance_to_wrap.core.register_file.registers_state\[166\] vssd1
+ vssd1 vccd1 vccd1 net2442 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_1113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11098__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08940_ net1046 team_03_WB.instance_to_wrap.core.register_file.registers_state\[843\]
+ net997 team_03_WB.instance_to_wrap.core.register_file.registers_state\[875\] net1062
+ vssd1 vssd1 vccd1 vccd1 _04882_ sky130_fd_sc_hd__a221o_1
XANTENNA__08907__C1 net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08871_ _04811_ _04812_ _04808_ vssd1 vssd1 vccd1 vccd1 _04813_ sky130_fd_sc_hd__a21oi_1
XANTENNA_clkbuf_leaf_131_wb_clk_i_A clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__07186__A1 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10015__B net67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07822_ _03761_ _03763_ net806 vssd1 vssd1 vccd1 vccd1 _03764_ sky130_fd_sc_hd__o21a_1
XANTENNA__10730__S net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06933__A1 net1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07605__A net1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09092__A net1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07753_ net1195 team_03_WB.instance_to_wrap.core.register_file.registers_state\[460\]
+ vssd1 vssd1 vccd1 vccd1 _03695_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_84_2105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08200__S net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11127__A net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07684_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[542\] net761
+ net740 _03625_ vssd1 vssd1 vccd1 vccd1 _03626_ sky130_fd_sc_hd__a211o_1
X_09423_ net541 _04446_ _04385_ vssd1 vssd1 vccd1 vccd1 _05365_ sky130_fd_sc_hd__o21a_1
XFILLER_0_149_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11690__B1 net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08781__S1 net1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout347_A _06804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13342__A net1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09354_ _05293_ _05295_ vssd1 vssd1 vccd1 vccd1 _05296_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout1089_A net1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07978__C net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06882__C team_03_WB.instance_to_wrap.core.decoder.inst\[25\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07340__A net1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08305_ net1236 team_03_WB.instance_to_wrap.core.register_file.registers_state\[472\]
+ net972 team_03_WB.instance_to_wrap.core.register_file.registers_state\[504\] net1212
+ vssd1 vssd1 vccd1 vccd1 _04247_ sky130_fd_sc_hd__o221a_1
XANTENNA__11442__B1 net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09285_ _05226_ vssd1 vssd1 vccd1 vccd1 _05227_ sky130_fd_sc_hd__inv_2
XANTENNA__07646__C1 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout514_A net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1256_A net1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09966__S net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08236_ net849 _04163_ _04177_ vssd1 vssd1 vccd1 vccd1 _04178_ sky130_fd_sc_hd__a21o_4
XFILLER_0_105_516 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_190 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15074__1460 vssd1 vssd1 vccd1 vccd1 _15074__1460/HI net1460 sky130_fd_sc_hd__conb_1
X_08167_ net1230 team_03_WB.instance_to_wrap.core.register_file.registers_state\[596\]
+ net959 team_03_WB.instance_to_wrap.core.register_file.registers_state\[628\] net918
+ vssd1 vssd1 vccd1 vccd1 _04109_ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout302_X net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_170_wb_clk_i_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout1044_X net1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07118_ net1251 _02808_ _02818_ net1163 vssd1 vssd1 vccd1 vccd1 _03060_ sky130_fd_sc_hd__a22oi_4
XFILLER_0_160_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_56_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08098_ net806 _04038_ _04039_ vssd1 vssd1 vccd1 vccd1 _04040_ sky130_fd_sc_hd__or3_1
XFILLER_0_63_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout883_A net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_390 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07049_ net614 _02990_ vssd1 vssd1 vccd1 vccd1 _02991_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_128_3009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1211_X net1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1309_X net1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_148_wb_clk_i clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_148_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__09797__S0 net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10060_ net27 net1039 net911 net2782 vssd1 vssd1 vccd1 vccd1 _02671_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_73_1875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_1886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout671_X net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_3345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08374__B1 net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout769_X net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_3356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10181__A0 _04646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10640__S net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06924__A1 net1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07582__D1 net1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_162_3692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout936_X net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10962_ team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[2\] net308 net689 vssd1
+ vssd1 vccd1 vccd1 _06543_ sky130_fd_sc_hd__a21o_1
X_13750_ clknet_leaf_178_wb_clk_i _01514_ _00115_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[104\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_173_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_1136 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_901 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12701_ net1388 vssd1 vssd1 vccd1 vccd1 _00465_ sky130_fd_sc_hd__inv_2
XANTENNA__08049__C net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11681__B1 net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07885__C1 net1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10893_ _06485_ _06486_ _06484_ vssd1 vssd1 vccd1 vccd1 _06487_ sky130_fd_sc_hd__o21a_2
X_13681_ clknet_leaf_141_wb_clk_i _01445_ _00046_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[35\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_78_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_155_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13252__A net1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12632_ net1376 vssd1 vssd1 vccd1 vccd1 _00396_ sky130_fd_sc_hd__inv_2
XFILLER_0_167_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_155_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11433__A0 net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12563_ net1256 vssd1 vssd1 vccd1 vccd1 _00327_ sky130_fd_sc_hd__inv_2
XFILLER_0_38_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07101__A1 team_03_WB.instance_to_wrap.core.decoder.inst\[23\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11514_ net265 net2739 net390 vssd1 vssd1 vccd1 vccd1 _01992_ sky130_fd_sc_hd__mux2_1
X_14302_ clknet_leaf_117_wb_clk_i _02066_ _00667_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[656\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12494_ net1270 vssd1 vssd1 vccd1 vccd1 _00258_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_672 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14233_ clknet_leaf_155_wb_clk_i _01997_ _00598_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[587\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_62_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11445_ net497 net626 _06572_ net395 net2151 vssd1 vssd1 vccd1 vccd1 _02044_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_117_2779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11736__A1 net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10539__A2 net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07396__S net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_169_3835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14164_ clknet_leaf_124_wb_clk_i _01928_ _00529_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[518\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_169_3846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08601__A1 net1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11376_ net491 net620 _06740_ net400 net2241 vssd1 vssd1 vccd1 vccd1 _02092_ sky130_fd_sc_hd__a32o_1
XANTENNA__08081__A net1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08601__B2 net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10327_ _06123_ _06125_ vssd1 vssd1 vccd1 vccd1 _06166_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_156_Right_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13115_ net1364 vssd1 vssd1 vccd1 vccd1 _00879_ sky130_fd_sc_hd__inv_2
X_14095_ clknet_leaf_137_wb_clk_i _01859_ _00460_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[449\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09905__A net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13046_ net1257 vssd1 vssd1 vccd1 vccd1 _00810_ sky130_fd_sc_hd__inv_2
X_10258_ _04030_ _06099_ vssd1 vssd1 vccd1 vccd1 _06100_ sky130_fd_sc_hd__and2b_1
Xfanout1230 net1233 vssd1 vssd1 vccd1 vccd1 net1230 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11646__S net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1241 net1246 vssd1 vssd1 vccd1 vccd1 net1241 sky130_fd_sc_hd__buf_4
X_10189_ _03460_ _06029_ vssd1 vssd1 vccd1 vccd1 _06031_ sky130_fd_sc_hd__or2_1
Xfanout1252 team_03_WB.instance_to_wrap.core.decoder.inst\[7\] vssd1 vssd1 vccd1 vccd1
+ net1252 sky130_fd_sc_hd__buf_4
XANTENNA__12331__A net1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1263 net1264 vssd1 vssd1 vccd1 vccd1 net1263 sky130_fd_sc_hd__clkbuf_2
Xfanout1274 net1277 vssd1 vssd1 vccd1 vccd1 net1274 sky130_fd_sc_hd__buf_4
Xfanout1285 net1286 vssd1 vssd1 vccd1 vccd1 net1285 sky130_fd_sc_hd__buf_4
Xfanout1296 net1298 vssd1 vssd1 vccd1 vccd1 net1296 sky130_fd_sc_hd__buf_4
XFILLER_0_89_823 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14997_ clknet_leaf_66_wb_clk_i net45 _01362_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_13948_ clknet_leaf_146_wb_clk_i _01712_ _00313_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[302\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09865__B1 _03944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_46 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_755 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10786__A net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13879_ clknet_leaf_113_wb_clk_i _01643_ _00244_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[233\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11234__X _06684_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_174_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07798__C net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_904 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10936__D net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1001 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09070_ net851 _04998_ _05011_ vssd1 vssd1 vccd1 vccd1 _05012_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_127_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08690__S net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08840__A1 net1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08021_ net1085 net894 team_03_WB.instance_to_wrap.core.register_file.registers_state\[17\]
+ vssd1 vssd1 vccd1 vccd1 _03963_ sky130_fd_sc_hd__o21a_1
XFILLER_0_126_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_823 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11727__A1 _06487_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold702 team_03_WB.instance_to_wrap.core.register_file.registers_state\[263\] vssd1
+ vssd1 vccd1 vccd1 net2195 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold713 team_03_WB.instance_to_wrap.core.register_file.registers_state\[925\] vssd1
+ vssd1 vccd1 vccd1 net2206 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold724 team_03_WB.instance_to_wrap.core.register_file.registers_state\[54\] vssd1
+ vssd1 vccd1 vccd1 net2217 sky130_fd_sc_hd__dlygate4sd3_1
Xhold735 team_03_WB.instance_to_wrap.CPU_DAT_O\[31\] vssd1 vssd1 vccd1 vccd1 net2228
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold746 team_03_WB.instance_to_wrap.core.register_file.registers_state\[757\] vssd1
+ vssd1 vccd1 vccd1 net2239 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold757 team_03_WB.instance_to_wrap.core.register_file.registers_state\[756\] vssd1
+ vssd1 vccd1 vccd1 net2250 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold768 team_03_WB.instance_to_wrap.core.register_file.registers_state\[161\] vssd1
+ vssd1 vccd1 vccd1 net2261 sky130_fd_sc_hd__dlygate4sd3_1
X_09972_ _05890_ net1965 net291 vssd1 vssd1 vccd1 vccd1 _02741_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_123_Right_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold779 team_03_WB.instance_to_wrap.core.register_file.registers_state\[806\] vssd1
+ vssd1 vccd1 vccd1 net2272 sky130_fd_sc_hd__dlygate4sd3_1
X_08923_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[11\] net997
+ net925 _04864_ vssd1 vssd1 vccd1 vccd1 _04865_ sky130_fd_sc_hd__o211a_1
XFILLER_0_23_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07159__A1 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout297_A _06499_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08854_ _04794_ _04795_ net858 vssd1 vssd1 vccd1 vccd1 _04796_ sky130_fd_sc_hd__a21o_1
X_07805_ net815 _03745_ _03746_ vssd1 vssd1 vccd1 vccd1 _03747_ sky130_fd_sc_hd__and3_1
X_08785_ net868 _04720_ _04726_ net852 vssd1 vssd1 vccd1 vccd1 _04727_ sky130_fd_sc_hd__a211o_1
XFILLER_0_98_119 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08108__B1 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout464_A net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_140_3242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07736_ _03669_ _03677_ _03660_ vssd1 vssd1 vccd1 vccd1 _03678_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_140_3253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08203__S0 net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08659__A1 net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07867__C1 net1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07667_ net739 _03605_ _03606_ _03607_ _03608_ vssd1 vssd1 vccd1 vccd1 _03609_ sky130_fd_sc_hd__o32a_1
XANTENNA_fanout631_A _06458_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1373_A net1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout729_A net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09406_ net548 _04296_ _04121_ vssd1 vssd1 vccd1 vccd1 _05348_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_1_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07598_ net1203 team_03_WB.instance_to_wrap.core.register_file.registers_state\[345\]
+ vssd1 vssd1 vccd1 vccd1 _03540_ sky130_fd_sc_hd__or2_1
XFILLER_0_30_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11415__A0 net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09337_ _05208_ _05211_ vssd1 vssd1 vccd1 vccd1 _05279_ sky130_fd_sc_hd__and2_1
XFILLER_0_36_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09084__A1 net1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1161_X net1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout517_X net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10769__A2 _06378_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11966__A1 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09268_ _03727_ _05150_ vssd1 vssd1 vccd1 vccd1 _05210_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_35_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11430__A3 _06756_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10086__A_N _05718_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_929 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08219_ net1061 _04158_ _04159_ vssd1 vssd1 vccd1 vccd1 _04161_ sky130_fd_sc_hd__or3_1
XFILLER_0_44_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10635__S net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09199_ _05073_ _05120_ _05140_ _04777_ _05127_ vssd1 vssd1 vccd1 vccd1 _05141_ sky130_fd_sc_hd__a221o_2
XANTENNA__12416__A net1402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11718__A1 net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11230_ net268 net2170 net488 vssd1 vssd1 vccd1 vccd1 _02181_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_1915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_891 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07398__A1 net1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout886_X net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11161_ net2478 net413 _06658_ net502 vssd1 vssd1 vccd1 vccd1 _02225_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_112_2676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_8_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10112_ _04807_ net660 _05954_ _03065_ vssd1 vssd1 vccd1 vccd1 _05956_ sky130_fd_sc_hd__a211oi_1
XANTENNA__07944__S net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_164_3732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11974__B _06751_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11092_ _06622_ net2374 net419 vssd1 vssd1 vccd1 vccd1 _02258_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_164_3743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08347__B1 net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10043_ net14 net1037 net909 net1964 vssd1 vssd1 vccd1 vccd1 _02688_ sky130_fd_sc_hd__o22a_1
X_14920_ clknet_leaf_42_wb_clk_i _02675_ _01285_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_O\[7\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__13247__A net1347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08898__A1 net1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold40 team_03_WB.instance_to_wrap.core.register_file.registers_state\[935\] vssd1
+ vssd1 vccd1 vccd1 net1533 sky130_fd_sc_hd__dlygate4sd3_1
Xhold51 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1010\] vssd1
+ vssd1 vccd1 vccd1 net1544 sky130_fd_sc_hd__dlygate4sd3_1
Xhold62 team_03_WB.instance_to_wrap.core.register_file.registers_state\[22\] vssd1
+ vssd1 vccd1 vccd1 net1555 sky130_fd_sc_hd__dlygate4sd3_1
X_14851_ clknet_leaf_66_wb_clk_i net1527 _01216_ vssd1 vssd1 vccd1 vccd1 net106 sky130_fd_sc_hd__dfrtp_1
XANTENNA_input25_A DAT_I[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold73 team_03_WB.instance_to_wrap.core.register_file.registers_state\[930\] vssd1
+ vssd1 vccd1 vccd1 net1566 sky130_fd_sc_hd__dlygate4sd3_1
Xhold84 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1005\] vssd1
+ vssd1 vccd1 vccd1 net1577 sky130_fd_sc_hd__dlygate4sd3_1
Xhold95 _02634_ vssd1 vssd1 vccd1 vccd1 net1588 sky130_fd_sc_hd__dlygate4sd3_1
X_13802_ clknet_leaf_3_wb_clk_i _01566_ _00167_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[156\]
+ sky130_fd_sc_hd__dfrtp_1
X_14782_ clknet_leaf_95_wb_clk_i _02546_ _01147_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_I\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09847__B1 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11994_ net297 net2541 net445 vssd1 vssd1 vccd1 vccd1 _01550_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13733_ clknet_leaf_10_wb_clk_i _01497_ _00098_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[87\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_168_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10945_ team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[5\] net306 vssd1 vssd1
+ vccd1 vccd1 _06529_ sky130_fd_sc_hd__nand2_2
XFILLER_0_86_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_45_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_45_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_42_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13664_ clknet_leaf_190_wb_clk_i _01428_ _00029_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_168_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10876_ _06470_ _06471_ _06472_ vssd1 vssd1 vccd1 vccd1 _06473_ sky130_fd_sc_hd__a21oi_4
XANTENNA__08076__A net1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11406__A0 net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12615_ net1369 vssd1 vssd1 vccd1 vccd1 _00379_ sky130_fd_sc_hd__inv_2
XANTENNA__10893__X _06487_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_2819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07411__C net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09075__A1 net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13595_ net1269 vssd1 vssd1 vccd1 vccd1 _01359_ sky130_fd_sc_hd__inv_2
XANTENNA__11957__A1 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08822__A1 net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12546_ net1296 vssd1 vssd1 vccd1 vccd1 _00310_ sky130_fd_sc_hd__inv_2
XFILLER_0_124_622 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08822__B2 net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12477_ net1389 vssd1 vssd1 vccd1 vccd1 _00241_ sky130_fd_sc_hd__inv_2
XFILLER_0_34_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_151_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_4 team_03_WB.instance_to_wrap.core.decoder.inst\[23\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_14216_ clknet_leaf_13_wb_clk_i _01980_ _00581_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[570\]
+ sky130_fd_sc_hd__dfrtp_1
X_11428_ net508 net265 _06756_ net398 net2520 vssd1 vssd1 vccd1 vccd1 _02056_ sky130_fd_sc_hd__a32o_1
XANTENNA__08015__S net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11185__A2 net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11359_ net709 _06473_ net695 vssd1 vssd1 vccd1 vccd1 _06732_ sky130_fd_sc_hd__and3_1
X_14147_ clknet_leaf_35_wb_clk_i _01911_ _00512_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[501\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_158_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08050__A2 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14078_ clknet_leaf_118_wb_clk_i _01842_ _00443_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[432\]
+ sky130_fd_sc_hd__dfrtp_1
X_13029_ net1348 vssd1 vssd1 vccd1 vccd1 _00793_ sky130_fd_sc_hd__inv_2
Xfanout1060 _02791_ vssd1 vssd1 vccd1 vccd1 net1060 sky130_fd_sc_hd__buf_2
Xfanout1071 net1074 vssd1 vssd1 vccd1 vccd1 net1071 sky130_fd_sc_hd__buf_4
XANTENNA__09550__A2 _04267_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11893__B1 net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1082 net1093 vssd1 vssd1 vccd1 vccd1 net1082 sky130_fd_sc_hd__clkbuf_4
Xfanout1093 _02787_ vssd1 vssd1 vccd1 vccd1 net1093 sky130_fd_sc_hd__buf_4
XFILLER_0_83_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_174_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08570_ net861 _04508_ _04511_ vssd1 vssd1 vccd1 vccd1 _04512_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_107_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06994__A team_03_WB.instance_to_wrap.core.decoder.inst\[13\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14984__Q team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[3\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07521_ _03461_ _03462_ vssd1 vssd1 vccd1 vccd1 _03463_ sky130_fd_sc_hd__and2_1
XFILLER_0_49_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_159_563 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08510__B1 net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07452_ net1089 net895 team_03_WB.instance_to_wrap.core.register_file.registers_state\[149\]
+ vssd1 vssd1 vccd1 vccd1 _03394_ sky130_fd_sc_hd__o21a_1
XANTENNA__07161__Y _03103_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_174_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_40 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11124__B net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07383_ net1171 team_03_WB.instance_to_wrap.core.register_file.registers_state\[351\]
+ net758 team_03_WB.instance_to_wrap.core.register_file.registers_state\[383\] net1123
+ vssd1 vssd1 vccd1 vccd1 _03325_ sky130_fd_sc_hd__o221a_1
XFILLER_0_18_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_2004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11948__A1 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_959 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09122_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[622\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[590\]
+ net976 vssd1 vssd1 vccd1 vccd1 _05064_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_44_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_44_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12070__A0 net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_599 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07616__A2 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08274__C1 net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_161_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10963__B _05798_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_110 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_2340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10620__A1 team_03_WB.instance_to_wrap.CPU_DAT_O\[9\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_115_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09053_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[431\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[399\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[303\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[271\]
+ net985 net1073 vssd1 vssd1 vccd1 vccd1 _04995_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_96_2351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07092__A3 net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11140__A net1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08004_ _03934_ _03941_ net617 _03925_ vssd1 vssd1 vccd1 vccd1 _03946_ sky130_fd_sc_hd__o211a_2
XFILLER_0_114_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_170_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold510 team_03_WB.instance_to_wrap.core.register_file.registers_state\[427\] vssd1
+ vssd1 vccd1 vccd1 net2003 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08026__C1 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_962 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold521 team_03_WB.instance_to_wrap.core.register_file.registers_state\[916\] vssd1
+ vssd1 vccd1 vccd1 net2014 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold532 team_03_WB.instance_to_wrap.core.register_file.registers_state\[173\] vssd1
+ vssd1 vccd1 vccd1 net2025 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_2259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold543 team_03_WB.instance_to_wrap.core.register_file.registers_state\[465\] vssd1
+ vssd1 vccd1 vccd1 net2036 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07049__B _02990_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold554 team_03_WB.instance_to_wrap.core.register_file.registers_state\[460\] vssd1
+ vssd1 vccd1 vccd1 net2047 sky130_fd_sc_hd__dlygate4sd3_1
Xhold565 team_03_WB.instance_to_wrap.core.register_file.registers_state\[254\] vssd1
+ vssd1 vccd1 vccd1 net2058 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1121_A net1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10923__A2 net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold576 team_03_WB.instance_to_wrap.core.register_file.registers_state\[426\] vssd1
+ vssd1 vccd1 vccd1 net2069 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1219_A net1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold587 team_03_WB.instance_to_wrap.core.register_file.registers_state\[408\] vssd1
+ vssd1 vccd1 vccd1 net2080 sky130_fd_sc_hd__dlygate4sd3_1
Xhold598 team_03_WB.instance_to_wrap.core.register_file.registers_state\[823\] vssd1
+ vssd1 vccd1 vccd1 net2091 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_70_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09955_ _03942_ net661 vssd1 vssd1 vccd1 vccd1 _05882_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout581_A net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout679_A net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10136__A0 _04267_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08906_ net1239 team_03_WB.instance_to_wrap.core.register_file.registers_state\[588\]
+ net979 team_03_WB.instance_to_wrap.core.register_file.registers_state\[620\] net926
+ vssd1 vssd1 vccd1 vccd1 _04848_ sky130_fd_sc_hd__o221a_1
X_09886_ _04816_ _05827_ net665 vssd1 vssd1 vccd1 vccd1 _05828_ sky130_fd_sc_hd__o21a_1
Xhold1210 team_03_WB.instance_to_wrap.core.register_file.registers_state\[591\] vssd1
+ vssd1 vccd1 vccd1 net2703 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1221 team_03_WB.instance_to_wrap.CPU_DAT_O\[6\] vssd1 vssd1 vccd1 vccd1 net2714
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07065__A net1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1232 team_03_WB.instance_to_wrap.core.register_file.registers_state\[741\] vssd1
+ vssd1 vccd1 vccd1 net2725 sky130_fd_sc_hd__dlygate4sd3_1
X_08837_ net565 _04650_ _04774_ _04778_ vssd1 vssd1 vccd1 vccd1 _04779_ sky130_fd_sc_hd__a211o_1
Xhold1243 team_03_WB.instance_to_wrap.CPU_DAT_O\[21\] vssd1 vssd1 vccd1 vccd1 net2736
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11884__B1 net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10978__X _06557_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10203__B net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout846_A net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1254 team_03_WB.instance_to_wrap.core.register_file.registers_state\[346\] vssd1
+ vssd1 vccd1 vccd1 net2747 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1265 team_03_WB.instance_to_wrap.core.register_file.registers_state\[343\] vssd1
+ vssd1 vccd1 vccd1 net2758 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1276 team_03_WB.instance_to_wrap.core.register_file.registers_state\[71\] vssd1
+ vssd1 vccd1 vccd1 net2769 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1287 team_03_WB.instance_to_wrap.CPU_DAT_O\[30\] vssd1 vssd1 vccd1 vccd1 net2780
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08595__S _02992_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08768_ net1208 _04709_ net848 vssd1 vssd1 vccd1 vccd1 _04710_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10439__A1 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11636__B1 net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07719_ net1197 team_03_WB.instance_to_wrap.core.register_file.registers_state\[717\]
+ net779 team_03_WB.instance_to_wrap.core.register_file.registers_state\[749\] net747
+ vssd1 vssd1 vccd1 vccd1 _03661_ sky130_fd_sc_hd__o221a_1
XFILLER_0_79_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout634_X net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08699_ net1241 team_03_WB.instance_to_wrap.core.register_file.registers_state\[456\]
+ net976 team_03_WB.instance_to_wrap.core.register_file.registers_state\[488\] net1211
+ vssd1 vssd1 vccd1 vccd1 _04641_ sky130_fd_sc_hd__o221a_1
XFILLER_0_67_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_1069 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1376_X net1376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10730_ team_03_WB.instance_to_wrap.core.pc.current_pc\[16\] _05812_ net603 vssd1
+ vssd1 vccd1 vccd1 _06357_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10661_ team_03_WB.instance_to_wrap.core.control_logic.instruction\[0\] team_03_WB.instance_to_wrap.CPU_DAT_O\[0\]
+ net846 vssd1 vssd1 vccd1 vccd1 _02467_ sky130_fd_sc_hd__mux2_1
XANTENNA__09057__A1 net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout801_X net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_157_3591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12400_ net1409 vssd1 vssd1 vccd1 vccd1 _00164_ sky130_fd_sc_hd__inv_2
XANTENNA__12061__A0 _06505_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07068__B1 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13380_ net1420 vssd1 vssd1 vccd1 vccd1 _01144_ sky130_fd_sc_hd__inv_2
X_10592_ _06301_ _06292_ team_03_WB.instance_to_wrap.READ_I net1142 vssd1 vssd1 vccd1
+ vccd1 _02533_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_106_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08804__A1 net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12331_ net1282 vssd1 vssd1 vccd1 vccd1 _00095_ sky130_fd_sc_hd__inv_2
XFILLER_0_133_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_161_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_114_2716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_299 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_2727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_163_wb_clk_i clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_163_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_105_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15050_ net1491 vssd1 vssd1 vccd1 vccd1 gpio_oeb[2] sky130_fd_sc_hd__buf_2
X_12262_ net1337 vssd1 vssd1 vccd1 vccd1 _00026_ sky130_fd_sc_hd__inv_2
XFILLER_0_32_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14001_ clknet_leaf_140_wb_clk_i _01765_ _00366_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[355\]
+ sky130_fd_sc_hd__dfrtp_1
X_11213_ _06456_ _06478_ vssd1 vssd1 vccd1 vccd1 _06681_ sky130_fd_sc_hd__nor2_1
XANTENNA__08568__B1 net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12193_ net1494 vssd1 vssd1 vccd1 vccd1 _02360_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_102_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07240__B1 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11144_ net628 _06648_ vssd1 vssd1 vccd1 vccd1 _06649_ sky130_fd_sc_hd__nor2_1
XFILLER_0_101_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11075_ _06615_ net2584 net417 vssd1 vssd1 vccd1 vccd1 _02268_ sky130_fd_sc_hd__mux2_1
X_14903_ clknet_leaf_86_wb_clk_i _02666_ _01268_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.pc.current_pc\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_10026_ net101 net99 net102 _05902_ vssd1 vssd1 vccd1 vccd1 _05903_ sky130_fd_sc_hd__and4_1
XANTENNA__09532__A2 _04354_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input28_X net28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10888__X _06483_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07543__A1 net1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08740__B1 net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11924__S net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14834_ clknet_leaf_90_wb_clk_i _02598_ _01199_ vssd1 vssd1 vccd1 vccd1 net155 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11890__A3 net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08718__S1 net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11627__B1 net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15053__1439 vssd1 vssd1 vccd1 vccd1 _15053__1439/HI net1439 sky130_fd_sc_hd__conb_1
X_14765_ clknet_leaf_48_wb_clk_i _02529_ _01130_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_11977_ _06413_ net2502 net443 vssd1 vssd1 vccd1 vccd1 _01567_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_336 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13716_ clknet_leaf_132_wb_clk_i _01480_ _00081_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[70\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10928_ net312 net310 net318 _02781_ vssd1 vssd1 vccd1 vccd1 _06515_ sky130_fd_sc_hd__a31o_1
X_14696_ clknet_leaf_63_wb_clk_i _02460_ _01061_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.ADR_I\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_156_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_758 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13647_ clknet_leaf_134_wb_clk_i _01411_ _00012_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09048__A1 net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10859_ team_03_WB.instance_to_wrap.core.decoder.inst\[10\] _06389_ _06390_ vssd1
+ vssd1 vccd1 vccd1 _06458_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_116_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12052__A0 _06454_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08256__C1 net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13578_ net1424 vssd1 vssd1 vccd1 vccd1 _01342_ sky130_fd_sc_hd__inv_2
XANTENNA__08534__A net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10275__S net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_964 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12529_ net1271 vssd1 vssd1 vccd1 vccd1 _00293_ sky130_fd_sc_hd__inv_2
XFILLER_0_169_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09917__X _05859_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_140_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11158__A2 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09220__A1 _03280_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08023__A2 net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10905__A2 _05697_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout308 _06396_ vssd1 vssd1 vccd1 vccd1 net308 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__07782__A1 team_03_WB.instance_to_wrap.core.decoder.inst\[12\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09740_ net537 _05679_ _05681_ vssd1 vssd1 vccd1 vccd1 _05682_ sky130_fd_sc_hd__o21ai_1
X_06952_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[165\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[133\]
+ net787 vssd1 vssd1 vccd1 vccd1 _02894_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
.ends

